module fake_aes_7106_n_780 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_780);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_780;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_227;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_76), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_99), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_78), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_138), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_1), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_153), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_48), .Y(n_199) );
NOR2xp67_ASAP7_75t_L g200 ( .A(n_65), .B(n_186), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_115), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_124), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_49), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_90), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_37), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_179), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_116), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_23), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_175), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_41), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_120), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_128), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_185), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_64), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_101), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_1), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_172), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_98), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_109), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_114), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_111), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_11), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_11), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_121), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_123), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_164), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_80), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_135), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_94), .Y(n_232) );
INVxp33_ASAP7_75t_L g233 ( .A(n_25), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_22), .Y(n_234) );
BUFx10_ASAP7_75t_L g235 ( .A(n_106), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_136), .Y(n_236) );
BUFx10_ASAP7_75t_L g237 ( .A(n_68), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_89), .Y(n_238) );
CKINVDCx14_ASAP7_75t_R g239 ( .A(n_156), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_53), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_102), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_31), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_139), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_118), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_66), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_77), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_61), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_60), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_70), .Y(n_249) );
BUFx2_ASAP7_75t_SL g250 ( .A(n_147), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_7), .Y(n_251) );
NOR2xp67_ASAP7_75t_L g252 ( .A(n_0), .B(n_180), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_84), .Y(n_253) );
BUFx5_ASAP7_75t_L g254 ( .A(n_20), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_9), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_19), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_103), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_96), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_162), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_131), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_129), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_170), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_148), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_169), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_57), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_178), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_165), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_108), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_61), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_161), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_146), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_183), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_184), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_157), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_144), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_35), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_158), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_143), .Y(n_278) );
CKINVDCx16_ASAP7_75t_R g279 ( .A(n_119), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_81), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_58), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_95), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_51), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_62), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_163), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_88), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_181), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_19), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_130), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_93), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_122), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_132), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_55), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_52), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_149), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_45), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_24), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_100), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_97), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_87), .B(n_110), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_238), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_235), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
BUFx8_ASAP7_75t_SL g304 ( .A(n_248), .Y(n_304) );
AOI22xp5_ASAP7_75t_SL g305 ( .A1(n_248), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_225), .B(n_3), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_254), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_238), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_235), .Y(n_310) );
BUFx12f_ASAP7_75t_L g311 ( .A(n_235), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_274), .B(n_4), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_238), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_243), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_233), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_225), .B(n_5), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_254), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_271), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_233), .B(n_8), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_271), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_269), .B(n_8), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_234), .B(n_9), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_272), .B(n_10), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_199), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_269), .B(n_10), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_273), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_199), .Y(n_329) );
INVx4_ASAP7_75t_L g330 ( .A(n_202), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_192), .Y(n_331) );
INVx5_ASAP7_75t_L g332 ( .A(n_202), .Y(n_332) );
OAI22x1_ASAP7_75t_SL g333 ( .A1(n_249), .A2(n_14), .B1(n_12), .B2(n_13), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_192), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_241), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_189), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_191), .Y(n_337) );
NAND2xp33_ASAP7_75t_SL g338 ( .A(n_324), .B(n_198), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_321), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_321), .Y(n_340) );
INVx8_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_306), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_336), .B(n_241), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_306), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_313), .Y(n_345) );
AND2x6_ASAP7_75t_L g346 ( .A(n_306), .B(n_219), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_332), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_304), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_302), .B(n_239), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_313), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_307), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_323), .A2(n_210), .B1(n_218), .B2(n_205), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_311), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_307), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
AO21x2_ASAP7_75t_L g358 ( .A1(n_325), .A2(n_300), .B(n_193), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_302), .B(n_224), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_336), .B(n_244), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_311), .B(n_250), .Y(n_362) );
NAND2xp33_ASAP7_75t_L g363 ( .A(n_310), .B(n_299), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_310), .B(n_279), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_198), .B1(n_230), .B2(n_201), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_310), .B(n_237), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_332), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_360), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_346), .A2(n_327), .B1(n_323), .B2(n_337), .Y(n_370) );
INVx5_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_366), .B(n_314), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_346), .A2(n_327), .B1(n_337), .B2(n_318), .Y(n_374) );
BUFx8_ASAP7_75t_L g375 ( .A(n_366), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_360), .Y(n_376) );
NAND2xp33_ASAP7_75t_L g377 ( .A(n_346), .B(n_314), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_360), .B(n_364), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_346), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_360), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
AND2x6_ASAP7_75t_SL g382 ( .A(n_348), .B(n_320), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_342), .B(n_328), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_355), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_201), .B1(n_232), .B2(n_230), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_363), .B(n_320), .C(n_312), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_344), .B(n_330), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_344), .B(n_330), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_341), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_354), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_346), .B(n_330), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_341), .B(n_237), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_354), .B(n_194), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_343), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_359), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_359), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g400 ( .A(n_338), .B(n_315), .C(n_265), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_361), .B(n_317), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_340), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_358), .A2(n_334), .B1(n_335), .B2(n_331), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_358), .B(n_326), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_349), .A2(n_329), .B1(n_242), .B2(n_245), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_340), .B(n_329), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_365), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_365), .A2(n_259), .B1(n_260), .B2(n_232), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_352), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_356), .A2(n_247), .B1(n_276), .B2(n_240), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_347), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_357), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_368), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_347), .B(n_204), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_347), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g418 ( .A1(n_367), .A2(n_283), .B(n_284), .C(n_281), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_396), .A2(n_295), .B1(n_292), .B2(n_209), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_396), .B(n_195), .Y(n_420) );
INVx5_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_411), .A2(n_197), .B(n_196), .Y(n_422) );
CKINVDCx8_ASAP7_75t_R g423 ( .A(n_382), .Y(n_423) );
O2A1O1Ixp33_ASAP7_75t_L g424 ( .A1(n_409), .A2(n_293), .B(n_294), .C(n_288), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_402), .B(n_203), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_414), .A2(n_211), .B(n_207), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_397), .B(n_305), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_375), .B(n_333), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_369), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_370), .A2(n_212), .B1(n_222), .B2(n_190), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_385), .A2(n_297), .B(n_252), .C(n_200), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_400), .A2(n_290), .B1(n_333), .B2(n_208), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_415), .A2(n_214), .B(n_213), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_381), .B(n_220), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_376), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_374), .A2(n_217), .B1(n_223), .B2(n_215), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_SL g438 ( .A1(n_406), .A2(n_226), .B(n_229), .C(n_228), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_388), .A2(n_253), .B(n_246), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_390), .A2(n_261), .B(n_257), .Y(n_440) );
BUFx12f_ASAP7_75t_L g441 ( .A(n_384), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_390), .A2(n_266), .B(n_262), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_380), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_374), .A2(n_268), .B1(n_270), .B2(n_267), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_391), .B(n_221), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_389), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_394), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_392), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_398), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_372), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_383), .A2(n_278), .B(n_275), .Y(n_451) );
BUFx4f_ASAP7_75t_L g452 ( .A(n_379), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_408), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_397), .B(n_216), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_378), .A2(n_287), .B(n_289), .C(n_286), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_400), .A2(n_418), .B(n_401), .C(n_377), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_371), .Y(n_457) );
OAI22x1_ASAP7_75t_L g458 ( .A1(n_410), .A2(n_255), .B1(n_256), .B2(n_251), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_405), .A2(n_263), .B(n_298), .C(n_227), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_371), .B(n_219), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_403), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_379), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_404), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_405), .A2(n_285), .B(n_264), .C(n_301), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_412), .B(n_407), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_407), .B(n_296), .Y(n_466) );
BUFx2_ASAP7_75t_SL g467 ( .A(n_417), .Y(n_467) );
NOR2xp33_ASAP7_75t_SL g468 ( .A(n_387), .B(n_236), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
NOR2xp33_ASAP7_75t_SL g470 ( .A(n_413), .B(n_258), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_416), .A2(n_206), .B1(n_231), .B2(n_277), .C(n_280), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_413), .B(n_282), .Y(n_472) );
BUFx12f_ASAP7_75t_L g473 ( .A(n_382), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_396), .B(n_291), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_396), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_411), .A2(n_309), .B(n_301), .Y(n_476) );
INVx2_ASAP7_75t_SL g477 ( .A(n_375), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_396), .Y(n_478) );
INVx4_ASAP7_75t_L g479 ( .A(n_381), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_396), .A2(n_316), .B1(n_322), .B2(n_319), .Y(n_480) );
AND2x4_ASAP7_75t_SL g481 ( .A(n_397), .B(n_316), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_396), .A2(n_316), .B1(n_322), .B2(n_319), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_399), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_373), .A2(n_351), .B(n_345), .C(n_17), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_409), .A2(n_17), .B(n_15), .C(n_16), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_411), .A2(n_351), .B(n_345), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_411), .A2(n_351), .B(n_345), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_375), .B(n_18), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_411), .A2(n_351), .B(n_345), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_373), .A2(n_351), .B(n_24), .C(n_21), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_379), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_411), .A2(n_82), .B(n_83), .C(n_79), .Y(n_492) );
AOI21x1_ASAP7_75t_L g493 ( .A1(n_393), .A2(n_86), .B(n_85), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_375), .B(n_26), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_396), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_456), .A2(n_29), .B(n_27), .C(n_28), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_475), .B(n_27), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_478), .B(n_28), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_453), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_495), .B(n_29), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_465), .B(n_30), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_486), .A2(n_489), .B(n_487), .Y(n_502) );
AOI221x1_ASAP7_75t_L g503 ( .A1(n_431), .A2(n_32), .B1(n_33), .B2(n_34), .C(n_35), .Y(n_503) );
AO32x2_ASAP7_75t_L g504 ( .A1(n_437), .A2(n_36), .A3(n_38), .B1(n_39), .B2(n_40), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_436), .B(n_38), .Y(n_505) );
BUFx10_ASAP7_75t_L g506 ( .A(n_477), .Y(n_506) );
BUFx10_ASAP7_75t_L g507 ( .A(n_488), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_420), .B(n_39), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_424), .A2(n_42), .B(n_43), .C(n_44), .Y(n_509) );
AOI21x1_ASAP7_75t_L g510 ( .A1(n_493), .A2(n_92), .B(n_91), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_422), .A2(n_46), .B(n_47), .C(n_48), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_461), .Y(n_512) );
NOR2xp67_ASAP7_75t_L g513 ( .A(n_473), .B(n_47), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_463), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_427), .B(n_49), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_429), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_427), .B(n_50), .Y(n_517) );
NOR2x1_ASAP7_75t_SL g518 ( .A(n_467), .B(n_54), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_447), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_479), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_435), .Y(n_521) );
NAND3x1_ASAP7_75t_L g522 ( .A(n_432), .B(n_56), .C(n_58), .Y(n_522) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_491), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_425), .B(n_59), .Y(n_524) );
NOR2xp67_ASAP7_75t_L g525 ( .A(n_428), .B(n_59), .Y(n_525) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_439), .A2(n_442), .B(n_440), .Y(n_527) );
AO31x2_ASAP7_75t_L g528 ( .A1(n_455), .A2(n_63), .A3(n_64), .B(n_65), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_443), .B(n_67), .Y(n_529) );
NOR2xp67_ASAP7_75t_L g530 ( .A(n_458), .B(n_69), .Y(n_530) );
CKINVDCx8_ASAP7_75t_R g531 ( .A(n_494), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_423), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g533 ( .A1(n_454), .A2(n_71), .B(n_72), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_460), .Y(n_534) );
BUFx4f_ASAP7_75t_L g535 ( .A(n_469), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_474), .B(n_72), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_444), .B(n_73), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_446), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_448), .Y(n_539) );
INVx4_ASAP7_75t_L g540 ( .A(n_421), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_449), .Y(n_541) );
INVx3_ASAP7_75t_L g542 ( .A(n_457), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_460), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_466), .B(n_74), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_421), .B(n_75), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_485), .Y(n_546) );
BUFx3_ASAP7_75t_L g547 ( .A(n_481), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_491), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_459), .A2(n_104), .B(n_105), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_470), .B(n_107), .Y(n_550) );
AO31x2_ASAP7_75t_L g551 ( .A1(n_480), .A2(n_482), .A3(n_476), .B(n_426), .Y(n_551) );
AND2x6_ASAP7_75t_L g552 ( .A(n_462), .B(n_112), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_433), .B(n_113), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_434), .B(n_187), .Y(n_554) );
HAxp5_ASAP7_75t_L g555 ( .A(n_471), .B(n_117), .CON(n_555), .SN(n_555) );
OAI22x1_ASAP7_75t_L g556 ( .A1(n_438), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_556) );
AOI21xp5_ASAP7_75t_SL g557 ( .A1(n_480), .A2(n_133), .B(n_134), .Y(n_557) );
OR2x6_ASAP7_75t_L g558 ( .A(n_445), .B(n_140), .Y(n_558) );
NAND2xp33_ASAP7_75t_L g559 ( .A(n_483), .B(n_141), .Y(n_559) );
BUFx2_ASAP7_75t_L g560 ( .A(n_452), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_492), .Y(n_561) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_451), .A2(n_150), .B(n_151), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_468), .B(n_152), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_472), .Y(n_564) );
OAI21xp5_ASAP7_75t_SL g565 ( .A1(n_452), .A2(n_154), .B(n_155), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_464), .A2(n_159), .B(n_160), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_450), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_419), .Y(n_568) );
INVx4_ASAP7_75t_L g569 ( .A(n_479), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_475), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_464), .A2(n_166), .B(n_168), .Y(n_571) );
NAND2xp33_ASAP7_75t_R g572 ( .A(n_427), .B(n_171), .Y(n_572) );
BUFx2_ASAP7_75t_SL g573 ( .A(n_477), .Y(n_573) );
AOI21x1_ASAP7_75t_L g574 ( .A1(n_493), .A2(n_173), .B(n_174), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_475), .B(n_177), .Y(n_575) );
AO31x2_ASAP7_75t_L g576 ( .A1(n_464), .A2(n_484), .A3(n_490), .B(n_431), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_568), .B(n_499), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_499), .B(n_516), .Y(n_578) );
OAI21x1_ASAP7_75t_SL g579 ( .A1(n_518), .A2(n_565), .B(n_549), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_569), .B(n_512), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_516), .B(n_514), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_538), .Y(n_582) );
NOR2x1_ASAP7_75t_SL g583 ( .A(n_558), .B(n_540), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_539), .Y(n_584) );
AO31x2_ASAP7_75t_L g585 ( .A1(n_556), .A2(n_503), .A3(n_546), .B(n_496), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_541), .B(n_521), .Y(n_586) );
BUFx2_ASAP7_75t_R g587 ( .A(n_531), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_497), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_532), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_498), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g591 ( .A(n_540), .B(n_560), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_500), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_529), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_519), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_537), .A2(n_544), .B(n_505), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_523), .Y(n_596) );
BUFx12f_ASAP7_75t_L g597 ( .A(n_506), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_528), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_547), .B(n_520), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_515), .B(n_517), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_528), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_528), .Y(n_602) );
INVx4_ASAP7_75t_L g603 ( .A(n_506), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_564), .B(n_524), .Y(n_604) );
OA21x2_ASAP7_75t_L g605 ( .A1(n_536), .A2(n_553), .B(n_575), .Y(n_605) );
AO31x2_ASAP7_75t_L g606 ( .A1(n_509), .A2(n_511), .A3(n_508), .B(n_563), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_542), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_572), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_504), .Y(n_609) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_550), .A2(n_557), .B(n_567), .Y(n_610) );
OA21x2_ASAP7_75t_L g611 ( .A1(n_554), .A2(n_545), .B(n_530), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_504), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_535), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_559), .A2(n_562), .B(n_548), .Y(n_614) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_523), .A2(n_526), .B(n_522), .Y(n_615) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_534), .B(n_543), .Y(n_616) );
OA21x2_ASAP7_75t_L g617 ( .A1(n_576), .A2(n_525), .B(n_555), .Y(n_617) );
OA21x2_ASAP7_75t_L g618 ( .A1(n_551), .A2(n_552), .B(n_513), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_507), .B(n_549), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_533), .A2(n_456), .B(n_527), .C(n_496), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_499), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_527), .A2(n_456), .B(n_501), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_527), .A2(n_456), .B(n_501), .Y(n_623) );
AO21x2_ASAP7_75t_L g624 ( .A1(n_561), .A2(n_571), .B(n_566), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_499), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_502), .A2(n_561), .B(n_464), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_499), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_527), .A2(n_456), .B(n_501), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_527), .A2(n_456), .B(n_501), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_533), .A2(n_456), .B(n_527), .C(n_496), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_499), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_568), .B(n_409), .Y(n_632) );
OR2x6_ASAP7_75t_L g633 ( .A(n_573), .B(n_430), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_570), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_502), .A2(n_561), .B(n_464), .Y(n_635) );
INVx4_ASAP7_75t_L g636 ( .A(n_569), .Y(n_636) );
NOR2xp67_ASAP7_75t_L g637 ( .A(n_569), .B(n_441), .Y(n_637) );
AOI21x1_ASAP7_75t_L g638 ( .A1(n_561), .A2(n_574), .B(n_510), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_502), .A2(n_561), .B(n_464), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_499), .Y(n_640) );
INVx6_ASAP7_75t_L g641 ( .A(n_506), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_519), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_586), .B(n_625), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_634), .Y(n_644) );
AO21x2_ASAP7_75t_L g645 ( .A1(n_626), .A2(n_639), .B(n_635), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_586), .B(n_631), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_621), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_627), .B(n_640), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_627), .B(n_640), .Y(n_649) );
BUFx2_ASAP7_75t_SL g650 ( .A(n_637), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_578), .B(n_581), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_582), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_636), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_598), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_584), .Y(n_655) );
BUFx3_ASAP7_75t_L g656 ( .A(n_597), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_632), .B(n_577), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_583), .B(n_580), .Y(n_658) );
INVx2_ASAP7_75t_SL g659 ( .A(n_641), .Y(n_659) );
OR2x6_ASAP7_75t_L g660 ( .A(n_633), .B(n_615), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_604), .B(n_600), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_594), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_601), .Y(n_663) );
AO21x2_ASAP7_75t_L g664 ( .A1(n_638), .A2(n_622), .B(n_629), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_641), .Y(n_665) );
NOR2xp67_ASAP7_75t_SL g666 ( .A(n_608), .B(n_611), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_642), .B(n_602), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_591), .Y(n_668) );
INVx6_ASAP7_75t_L g669 ( .A(n_603), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_591), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_607), .B(n_596), .Y(n_671) );
AO21x2_ASAP7_75t_L g672 ( .A1(n_622), .A2(n_629), .B(n_623), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_603), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_593), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_588), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_633), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_590), .Y(n_677) );
AO21x2_ASAP7_75t_L g678 ( .A1(n_623), .A2(n_628), .B(n_614), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_592), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_620), .B(n_630), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_609), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_612), .Y(n_682) );
BUFx2_ASAP7_75t_L g683 ( .A(n_618), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_628), .B(n_595), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_617), .Y(n_685) );
OR2x6_ASAP7_75t_L g686 ( .A(n_660), .B(n_579), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_661), .B(n_616), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_662), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_654), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_684), .B(n_617), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_680), .B(n_606), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_663), .Y(n_692) );
INVx5_ASAP7_75t_L g693 ( .A(n_653), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_672), .B(n_606), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_651), .B(n_585), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_667), .B(n_619), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_650), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_653), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_643), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_658), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_648), .B(n_605), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_648), .B(n_624), .Y(n_702) );
INVx4_ASAP7_75t_L g703 ( .A(n_658), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_681), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_682), .Y(n_705) );
INVx3_ASAP7_75t_L g706 ( .A(n_660), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_649), .B(n_646), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_674), .B(n_599), .Y(n_708) );
AND2x4_ASAP7_75t_L g709 ( .A(n_660), .B(n_610), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_675), .B(n_599), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_647), .Y(n_711) );
NAND2x1_ASAP7_75t_L g712 ( .A(n_703), .B(n_666), .Y(n_712) );
INVxp67_ASAP7_75t_L g713 ( .A(n_688), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_693), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_707), .B(n_677), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_699), .B(n_679), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_695), .B(n_678), .Y(n_717) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_703), .B(n_653), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_686), .B(n_685), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_711), .B(n_657), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_700), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_690), .B(n_664), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_691), .B(n_644), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_686), .B(n_683), .Y(n_724) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_698), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_686), .B(n_683), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_704), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_705), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_705), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_702), .B(n_645), .Y(n_730) );
INVxp67_ASAP7_75t_L g731 ( .A(n_708), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_697), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_727), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_728), .Y(n_734) );
AND2x4_ASAP7_75t_L g735 ( .A(n_724), .B(n_706), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_729), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_720), .B(n_701), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_715), .B(n_689), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_723), .B(n_689), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_730), .B(n_696), .Y(n_740) );
INVx2_ASAP7_75t_SL g741 ( .A(n_718), .Y(n_741) );
NOR2xp33_ASAP7_75t_SL g742 ( .A(n_732), .B(n_587), .Y(n_742) );
BUFx3_ASAP7_75t_L g743 ( .A(n_714), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_713), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_716), .B(n_692), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_717), .B(n_696), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_724), .B(n_726), .Y(n_747) );
OR2x6_ASAP7_75t_L g748 ( .A(n_741), .B(n_712), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_747), .B(n_719), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_742), .A2(n_731), .B1(n_676), .B2(n_732), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_733), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_734), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_736), .Y(n_753) );
INVxp67_ASAP7_75t_L g754 ( .A(n_744), .Y(n_754) );
OAI21xp33_ASAP7_75t_SL g755 ( .A1(n_741), .A2(n_725), .B(n_721), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_743), .Y(n_756) );
O2A1O1Ixp33_ASAP7_75t_L g757 ( .A1(n_755), .A2(n_710), .B(n_673), .C(n_687), .Y(n_757) );
AOI211xp5_ASAP7_75t_L g758 ( .A1(n_755), .A2(n_747), .B(n_743), .C(n_735), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_756), .Y(n_759) );
OAI322xp33_ASAP7_75t_L g760 ( .A1(n_754), .A2(n_740), .A3(n_746), .B1(n_738), .B2(n_745), .C1(n_737), .C2(n_739), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_751), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_752), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_753), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_758), .A2(n_750), .B1(n_748), .B2(n_749), .Y(n_764) );
NOR2xp67_ASAP7_75t_SL g765 ( .A(n_759), .B(n_656), .Y(n_765) );
AOI21xp33_ASAP7_75t_L g766 ( .A1(n_757), .A2(n_665), .B(n_659), .Y(n_766) );
NOR3xp33_ASAP7_75t_SL g767 ( .A(n_760), .B(n_589), .C(n_613), .Y(n_767) );
AOI211xp5_ASAP7_75t_SL g768 ( .A1(n_764), .A2(n_706), .B(n_670), .C(n_668), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_767), .A2(n_763), .B1(n_762), .B2(n_761), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_768), .B(n_765), .C(n_766), .Y(n_770) );
XNOR2xp5_ASAP7_75t_L g771 ( .A(n_770), .B(n_769), .Y(n_771) );
NOR2xp33_ASAP7_75t_R g772 ( .A(n_771), .B(n_669), .Y(n_772) );
BUFx2_ASAP7_75t_L g773 ( .A(n_772), .Y(n_773) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_773), .Y(n_774) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_774), .A2(n_655), .B(n_652), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_775), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_776), .Y(n_777) );
OR2x6_ASAP7_75t_L g778 ( .A(n_777), .B(n_671), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_778), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_779), .A2(n_694), .B1(n_722), .B2(n_709), .Y(n_780) );
endmodule