module fake_jpeg_652_n_688 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_688);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_688;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_514;
wire n_242;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_63),
.Y(n_219)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_64),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_65),
.B(n_116),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_9),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_66),
.B(n_75),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_70),
.Y(n_198)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_73),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_9),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_76),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_18),
.B(n_8),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_80),
.B(n_82),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_84),
.B(n_98),
.Y(n_169)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_89),
.Y(n_191)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_91),
.Y(n_222)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_95),
.Y(n_226)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_8),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_20),
.B(n_21),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_99),
.B(n_112),
.Y(n_174)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_10),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_124),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_20),
.B(n_10),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_47),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_117),
.B(n_118),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_31),
.B(n_7),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_22),
.Y(n_119)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_120),
.B(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_21),
.B(n_7),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_23),
.B(n_11),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_33),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_39),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_60),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_31),
.Y(n_129)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_129),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_41),
.Y(n_132)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_78),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_134),
.B(n_161),
.Y(n_255)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_80),
.B(n_53),
.CON(n_139),
.SN(n_139)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_139),
.B(n_170),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_75),
.A2(n_28),
.B(n_55),
.C(n_50),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_144),
.B(n_225),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_60),
.B1(n_59),
.B2(n_48),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_158),
.A2(n_215),
.B1(n_33),
.B2(n_44),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_61),
.B(n_28),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_77),
.B(n_23),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_166),
.B(n_178),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_85),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_95),
.B(n_55),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_179),
.B(n_192),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_62),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_190),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_125),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_209),
.Y(n_228)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_67),
.Y(n_197)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_69),
.Y(n_199)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_129),
.A2(n_43),
.B1(n_31),
.B2(n_40),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g299 ( 
.A1(n_200),
.A2(n_1),
.B1(n_18),
.B2(n_160),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_74),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_204),
.Y(n_306)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_72),
.Y(n_205)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_79),
.Y(n_207)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_74),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_111),
.B(n_132),
.C(n_91),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_59),
.C(n_42),
.Y(n_238)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_106),
.A2(n_60),
.B1(n_59),
.B2(n_42),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_216),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_113),
.Y(n_217)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_115),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_142),
.Y(n_233)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_92),
.Y(n_223)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_63),
.Y(n_224)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_86),
.B(n_50),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_154),
.A2(n_96),
.B1(n_32),
.B2(n_44),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_227),
.A2(n_253),
.B1(n_269),
.B2(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_32),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_229),
.B(n_234),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_230),
.A2(n_245),
.B1(n_248),
.B2(n_303),
.Y(n_357)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_233),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_104),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_169),
.B(n_103),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_236),
.B(n_240),
.Y(n_324)
);

CKINVDCx12_ASAP7_75t_R g237 ( 
.A(n_221),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_237),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_238),
.B(n_281),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_239),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_174),
.B(n_102),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_174),
.B(n_110),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_241),
.B(n_244),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_181),
.B(n_110),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_203),
.A2(n_48),
.B1(n_42),
.B2(n_31),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_154),
.A2(n_48),
.B1(n_93),
.B2(n_86),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_247),
.A2(n_299),
.B1(n_137),
.B2(n_138),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_209),
.A2(n_40),
.B1(n_101),
.B2(n_93),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_101),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_249),
.B(n_250),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_40),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_40),
.B1(n_52),
.B2(n_2),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_254),
.Y(n_323)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_257),
.Y(n_346)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_150),
.Y(n_258)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_261),
.Y(n_353)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_165),
.Y(n_265)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_148),
.A2(n_52),
.B(n_13),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_267),
.B(n_159),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_173),
.B(n_146),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_268),
.B(n_270),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_184),
.A2(n_6),
.B1(n_17),
.B2(n_2),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_141),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_148),
.B(n_0),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_271),
.B(n_276),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_162),
.A2(n_6),
.B1(n_17),
.B2(n_2),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_273),
.A2(n_289),
.B1(n_295),
.B2(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_151),
.Y(n_274)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_156),
.B(n_13),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_142),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_279),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_152),
.B(n_18),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_245),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_141),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_280),
.A2(n_176),
.B(n_189),
.C(n_172),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_222),
.B(n_0),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_206),
.A2(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_136),
.B(n_14),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_287),
.Y(n_319)
);

CKINVDCx12_ASAP7_75t_R g284 ( 
.A(n_221),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_284),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_163),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_165),
.Y(n_288)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_191),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_202),
.Y(n_291)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_15),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_300),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_164),
.A2(n_4),
.B1(n_5),
.B2(n_13),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_140),
.Y(n_296)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_208),
.A2(n_5),
.B1(n_16),
.B2(n_17),
.Y(n_297)
);

INVx5_ASAP7_75t_SL g298 ( 
.A(n_168),
.Y(n_298)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_171),
.Y(n_301)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_175),
.B(n_18),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_140),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_200),
.A2(n_133),
.B1(n_135),
.B2(n_199),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_133),
.Y(n_304)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g305 ( 
.A(n_172),
.Y(n_305)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

OA22x2_ASAP7_75t_L g307 ( 
.A1(n_186),
.A2(n_185),
.B1(n_167),
.B2(n_217),
.Y(n_307)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_307),
.A2(n_196),
.B1(n_140),
.B2(n_157),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_313),
.B(n_326),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_275),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_328),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_300),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_255),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_285),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_262),
.A2(n_186),
.B1(n_190),
.B2(n_145),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_332),
.A2(n_369),
.B1(n_348),
.B2(n_350),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_262),
.A2(n_135),
.B1(n_183),
.B2(n_145),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_333),
.A2(n_348),
.B1(n_352),
.B2(n_298),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_296),
.Y(n_394)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_235),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_336),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_278),
.B(n_155),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_337),
.B(n_338),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_254),
.B(n_155),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_235),
.Y(n_339)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_341),
.A2(n_246),
.B(n_306),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_256),
.B(n_183),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_358),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_290),
.A2(n_147),
.B1(n_149),
.B2(n_153),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_157),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_271),
.A2(n_147),
.B1(n_149),
.B2(n_153),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_243),
.Y(n_354)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_354),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_292),
.C(n_259),
.Y(n_387)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_243),
.Y(n_356)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_280),
.B(n_281),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_228),
.B(n_196),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_270),
.C(n_279),
.Y(n_374)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_252),
.Y(n_361)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_252),
.Y(n_362)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_362),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_SL g363 ( 
.A(n_248),
.B(n_267),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_363),
.A2(n_306),
.B(n_301),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_281),
.B(n_238),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_364),
.Y(n_376)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_259),
.Y(n_366)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_229),
.A2(n_167),
.B1(n_177),
.B2(n_180),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

AO22x1_ASAP7_75t_SL g371 ( 
.A1(n_344),
.A2(n_303),
.B1(n_230),
.B2(n_307),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_371),
.A2(n_397),
.B(n_345),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_341),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_374),
.B(n_361),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_274),
.C(n_258),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_416),
.C(n_368),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_357),
.A2(n_273),
.B1(n_299),
.B2(n_307),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_377),
.B(n_381),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_316),
.A2(n_264),
.B1(n_307),
.B2(n_299),
.Y(n_378)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_378),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_379),
.A2(n_388),
.B1(n_334),
.B2(n_331),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_357),
.A2(n_299),
.B1(n_177),
.B2(n_180),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_382),
.B(n_394),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_287),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_383),
.B(n_398),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_385),
.A2(n_400),
.B(n_315),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_176),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_393),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_387),
.B(n_366),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g393 ( 
.A(n_324),
.B(n_189),
.Y(n_393)
);

INVx8_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_323),
.B(n_272),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_294),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_399),
.B(n_362),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_327),
.B(n_272),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_403),
.B(n_411),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_337),
.B(n_266),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_406),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_344),
.B(n_266),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_292),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_410),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_327),
.B(n_231),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_319),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_317),
.B(n_291),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_412),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_294),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_417),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_342),
.B(n_231),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_414),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_308),
.Y(n_415)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_415),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_355),
.B(n_257),
.C(n_232),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_304),
.Y(n_417)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_359),
.Y(n_418)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_418),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_392),
.A2(n_313),
.B1(n_358),
.B2(n_363),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_419),
.B(n_451),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_400),
.A2(n_312),
.B(n_350),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_424),
.A2(n_426),
.B(n_397),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g475 ( 
.A(n_425),
.B(n_443),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_385),
.A2(n_246),
.B(n_347),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_392),
.A2(n_325),
.B(n_340),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_427),
.A2(n_440),
.B(n_452),
.Y(n_476)
);

OA22x2_ASAP7_75t_L g429 ( 
.A1(n_379),
.A2(n_351),
.B1(n_349),
.B2(n_353),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_429),
.A2(n_371),
.B(n_381),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_433),
.A2(n_370),
.B1(n_374),
.B2(n_399),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_376),
.B(n_318),
.C(n_367),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_439),
.B(n_446),
.C(n_450),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_392),
.A2(n_365),
.B(n_346),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_441),
.B(n_397),
.Y(n_464)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_384),
.Y(n_444)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_445),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_311),
.C(n_343),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_447),
.B(n_456),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_375),
.B(n_322),
.C(n_309),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_388),
.A2(n_263),
.B1(n_260),
.B2(n_286),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_322),
.C(n_309),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_453),
.B(n_415),
.C(n_401),
.Y(n_491)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_396),
.B(n_391),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_458),
.B(n_387),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_411),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_460),
.B(n_461),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_449),
.B(n_373),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_462),
.A2(n_480),
.B(n_493),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_464),
.A2(n_419),
.B(n_429),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_420),
.A2(n_396),
.B1(n_395),
.B2(n_371),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_466),
.A2(n_478),
.B1(n_482),
.B2(n_441),
.Y(n_504)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_435),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_468),
.B(n_439),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_469),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_454),
.Y(n_470)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_405),
.Y(n_471)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_472),
.B(n_436),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_459),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_473),
.B(n_484),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_449),
.B(n_422),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_474),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_420),
.A2(n_395),
.B1(n_371),
.B2(n_386),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_422),
.B(n_391),
.Y(n_479)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_479),
.Y(n_511)
);

A2O1A1O1Ixp25_ASAP7_75t_L g480 ( 
.A1(n_427),
.A2(n_413),
.B(n_406),
.C(n_409),
.D(n_399),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_441),
.A2(n_417),
.B1(n_377),
.B2(n_393),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_448),
.B(n_457),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_483),
.B(n_486),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_430),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_432),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_448),
.Y(n_488)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_428),
.A2(n_394),
.B1(n_387),
.B2(n_410),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_489),
.A2(n_445),
.B1(n_437),
.B2(n_431),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_491),
.B(n_490),
.C(n_496),
.Y(n_530)
);

NOR2x1_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_408),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_492),
.B(n_496),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_452),
.A2(n_407),
.B(n_345),
.Y(n_493)
);

INVx13_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_494),
.Y(n_501)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_442),
.Y(n_495)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_495),
.Y(n_521)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_446),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_444),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_497),
.A2(n_434),
.B1(n_335),
.B2(n_455),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_425),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_498),
.B(n_520),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_423),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_499),
.B(n_506),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_462),
.A2(n_424),
.B(n_426),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_503),
.A2(n_532),
.B(n_480),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_504),
.A2(n_522),
.B1(n_533),
.B2(n_469),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_505),
.B(n_510),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_432),
.Y(n_506)
);

INVxp33_ASAP7_75t_SL g507 ( 
.A(n_486),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_507),
.B(n_509),
.Y(n_539)
);

OAI32xp33_ASAP7_75t_L g509 ( 
.A1(n_479),
.A2(n_429),
.A3(n_447),
.B1(n_440),
.B2(n_443),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_488),
.B(n_453),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_514),
.B(n_517),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_464),
.A2(n_434),
.B1(n_438),
.B2(n_429),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_515),
.A2(n_469),
.B1(n_493),
.B2(n_464),
.Y(n_535)
);

OAI21xp33_ASAP7_75t_L g516 ( 
.A1(n_476),
.A2(n_450),
.B(n_438),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_516),
.B(n_528),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_474),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_475),
.B(n_456),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_466),
.A2(n_482),
.B1(n_469),
.B2(n_478),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_487),
.B(n_436),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_523),
.B(n_404),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_483),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_524),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_527),
.B(n_408),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_484),
.B(n_421),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_487),
.C(n_491),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_460),
.B(n_437),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_431),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_535),
.A2(n_543),
.B1(n_547),
.B2(n_553),
.Y(n_587)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_536),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_537),
.B(n_559),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_503),
.A2(n_476),
.B(n_492),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_538),
.A2(n_548),
.B(n_549),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_540),
.A2(n_545),
.B1(n_551),
.B2(n_557),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_518),
.A2(n_463),
.B1(n_481),
.B2(n_471),
.Y(n_542)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_542),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_500),
.A2(n_489),
.B1(n_463),
.B2(n_470),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_521),
.Y(n_544)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_544),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_522),
.A2(n_492),
.B1(n_480),
.B2(n_467),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_500),
.A2(n_490),
.B1(n_495),
.B2(n_497),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_513),
.A2(n_526),
.B(n_512),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_523),
.B(n_472),
.C(n_485),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_550),
.B(n_554),
.C(n_556),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_504),
.A2(n_465),
.B1(n_485),
.B2(n_477),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_513),
.A2(n_418),
.B(n_477),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_552),
.B(n_505),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_529),
.A2(n_467),
.B1(n_465),
.B2(n_494),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_308),
.C(n_320),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_498),
.B(n_520),
.C(n_514),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_517),
.A2(n_524),
.B1(n_511),
.B2(n_508),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_SL g571 ( 
.A(n_558),
.B(n_509),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_527),
.B(n_320),
.C(n_404),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_560),
.B(n_501),
.C(n_533),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_515),
.A2(n_494),
.B1(n_380),
.B2(n_402),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_561),
.A2(n_567),
.B1(n_501),
.B2(n_335),
.Y(n_589)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_562),
.Y(n_588)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_519),
.Y(n_564)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_564),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_505),
.A2(n_380),
.B1(n_390),
.B2(n_401),
.Y(n_567)
);

AOI21xp33_ASAP7_75t_L g568 ( 
.A1(n_541),
.A2(n_526),
.B(n_525),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_568),
.B(n_572),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_571),
.B(n_573),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_546),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_519),
.C(n_502),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_575),
.B(n_584),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_SL g576 ( 
.A(n_558),
.B(n_518),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_576),
.B(n_578),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_577),
.A2(n_549),
.B(n_539),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_SL g578 ( 
.A(n_563),
.B(n_502),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_534),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_582),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_534),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_546),
.B(n_525),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_556),
.B(n_511),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_585),
.B(n_586),
.C(n_593),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_508),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_589),
.A2(n_561),
.B1(n_551),
.B2(n_545),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_390),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_591),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_554),
.B(n_321),
.C(n_261),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_555),
.B(n_380),
.Y(n_594)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_594),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_580),
.B(n_560),
.C(n_547),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_596),
.B(n_597),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_580),
.B(n_570),
.C(n_575),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_570),
.B(n_585),
.C(n_582),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_600),
.B(n_613),
.C(n_616),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_601),
.A2(n_329),
.B(n_242),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_594),
.B(n_555),
.Y(n_605)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_605),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_607),
.A2(n_609),
.B1(n_592),
.B2(n_576),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_574),
.A2(n_566),
.B1(n_535),
.B2(n_543),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_608),
.A2(n_607),
.B1(n_604),
.B2(n_609),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_579),
.A2(n_539),
.B1(n_557),
.B2(n_566),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_589),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_610),
.B(n_615),
.Y(n_635)
);

AOI322xp5_ASAP7_75t_L g612 ( 
.A1(n_569),
.A2(n_548),
.A3(n_552),
.B1(n_564),
.B2(n_538),
.C1(n_544),
.C2(n_562),
.Y(n_612)
);

OAI321xp33_ASAP7_75t_L g633 ( 
.A1(n_612),
.A2(n_571),
.A3(n_359),
.B1(n_305),
.B2(n_242),
.C(n_239),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_573),
.B(n_553),
.C(n_567),
.Y(n_613)
);

BUFx12_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_614),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_583),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_581),
.B(n_565),
.C(n_321),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_590),
.Y(n_617)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_617),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_587),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_618),
.B(n_626),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_613),
.B(n_578),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_619),
.B(n_631),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_601),
.A2(n_592),
.B(n_574),
.Y(n_621)
);

AO21x1_ASAP7_75t_L g640 ( 
.A1(n_621),
.A2(n_634),
.B(n_625),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_588),
.Y(n_625)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_625),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_598),
.B(n_587),
.Y(n_626)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_616),
.Y(n_627)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_627),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_628),
.A2(n_637),
.B1(n_608),
.B2(n_602),
.Y(n_645)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_617),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_630),
.B(n_632),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_603),
.B(n_593),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_604),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_633),
.A2(n_636),
.B(n_634),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_606),
.B(n_329),
.Y(n_636)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_640),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_622),
.B(n_597),
.C(n_620),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_641),
.B(n_642),
.Y(n_663)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_622),
.B(n_611),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_635),
.A2(n_623),
.B1(n_637),
.B2(n_621),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_643),
.B(n_646),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_SL g655 ( 
.A1(n_644),
.A2(n_647),
.B1(n_624),
.B2(n_629),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_645),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_618),
.B(n_600),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_628),
.A2(n_599),
.B1(n_602),
.B2(n_596),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_627),
.A2(n_599),
.B1(n_614),
.B2(n_595),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_649),
.B(n_650),
.Y(n_658)
);

BUFx24_ASAP7_75t_SL g650 ( 
.A(n_619),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_631),
.B(n_595),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_653),
.A2(n_636),
.B(n_614),
.Y(n_656)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_655),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_656),
.B(n_659),
.Y(n_666)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_642),
.B(n_286),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_641),
.B(n_260),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_660),
.B(n_661),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_652),
.B(n_263),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_651),
.B(n_356),
.C(n_354),
.Y(n_664)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_664),
.Y(n_669)
);

AOI31xp67_ASAP7_75t_L g665 ( 
.A1(n_648),
.A2(n_640),
.A3(n_638),
.B(n_645),
.Y(n_665)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_665),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_657),
.B(n_639),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_667),
.B(n_336),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_654),
.A2(n_647),
.B(n_651),
.Y(n_670)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_670),
.A2(n_657),
.B(n_658),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_663),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_672),
.A2(n_674),
.B(n_305),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_662),
.A2(n_251),
.B(n_305),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_675),
.B(n_676),
.Y(n_681)
);

BUFx24_ASAP7_75t_SL g676 ( 
.A(n_671),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_670),
.A2(n_664),
.B(n_659),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_677),
.B(n_669),
.C(n_668),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_SL g682 ( 
.A1(n_678),
.A2(n_679),
.B(n_673),
.C(n_674),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_680),
.B(n_682),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_681),
.A2(n_666),
.B(n_339),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_684),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_685),
.A2(n_683),
.B(n_265),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_686),
.B(n_288),
.C(n_157),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_687),
.A2(n_188),
.B(n_311),
.C(n_284),
.Y(n_688)
);


endmodule