module fake_jpeg_3529_n_179 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_0),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_51),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_67),
.B1(n_52),
.B2(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_66),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_44),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_67),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_54),
.B1(n_47),
.B2(n_46),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_68),
.B1(n_51),
.B2(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_53),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_86),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_57),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_64),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_33),
.C(n_29),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_71),
.B1(n_74),
.B2(n_53),
.Y(n_99)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_62),
.B(n_56),
.C(n_45),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_85),
.B(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_68),
.B1(n_60),
.B2(n_52),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_108),
.B1(n_95),
.B2(n_4),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_106),
.B1(n_95),
.B2(n_4),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_91),
.B1(n_97),
.B2(n_85),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_1),
.B(n_6),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_8),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_59),
.B1(n_58),
.B2(n_3),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_59),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_7),
.Y(n_128)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_6),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_123),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_89),
.B(n_93),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_124),
.B(n_127),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_1),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_28),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_128),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_7),
.B(n_8),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_105),
.B(n_10),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_131),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_25),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.C(n_104),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_24),
.C(n_23),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_141),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_125),
.B(n_13),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_104),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_9),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_149),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_156),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_137),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_136),
.B(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_161),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_12),
.B(n_14),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_135),
.C(n_144),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_163),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_157),
.B1(n_154),
.B2(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_149),
.C(n_150),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_160),
.B(n_154),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_171),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_167),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_165),
.B(n_158),
.C(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_170),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_168),
.B1(n_17),
.B2(n_18),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_19),
.B1(n_15),
.B2(n_16),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_15),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_16),
.Y(n_179)
);


endmodule