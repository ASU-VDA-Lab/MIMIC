module real_aes_536_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g186 ( .A(n_0), .B(n_133), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_1), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_2), .B(n_117), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_3), .B(n_135), .Y(n_535) );
INVx1_ASAP7_75t_L g124 ( .A(n_4), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_5), .B(n_117), .Y(n_116) );
NAND2xp33_ASAP7_75t_SL g230 ( .A(n_6), .B(n_123), .Y(n_230) );
INVx1_ASAP7_75t_L g222 ( .A(n_7), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_8), .Y(n_443) );
AND2x2_ASAP7_75t_L g111 ( .A(n_9), .B(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g473 ( .A(n_10), .B(n_228), .Y(n_473) );
AND2x2_ASAP7_75t_L g537 ( .A(n_11), .B(n_162), .Y(n_537) );
INVx2_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_13), .B(n_135), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_14), .Y(n_428) );
AOI221x1_ASAP7_75t_L g225 ( .A1(n_15), .A2(n_126), .B1(n_226), .B2(n_228), .C(n_229), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_16), .B(n_117), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_17), .B(n_117), .Y(n_492) );
INVx1_ASAP7_75t_L g432 ( .A(n_18), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_19), .A2(n_65), .B1(n_422), .B2(n_423), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_19), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_20), .A2(n_89), .B1(n_117), .B2(n_166), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_21), .A2(n_126), .B(n_131), .Y(n_125) );
AOI221xp5_ASAP7_75t_SL g196 ( .A1(n_22), .A2(n_36), .B1(n_117), .B2(n_126), .C(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_23), .B(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g114 ( .A(n_24), .B(n_88), .Y(n_114) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_24), .A2(n_88), .B(n_113), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_25), .B(n_135), .Y(n_213) );
INVxp67_ASAP7_75t_L g224 ( .A(n_26), .Y(n_224) );
AND2x2_ASAP7_75t_L g157 ( .A(n_27), .B(n_147), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_28), .A2(n_126), .B(n_185), .Y(n_184) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_29), .A2(n_228), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_30), .B(n_135), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_31), .A2(n_126), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_32), .B(n_135), .Y(n_508) );
AND2x2_ASAP7_75t_L g123 ( .A(n_33), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g127 ( .A(n_33), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g174 ( .A(n_33), .Y(n_174) );
OR2x6_ASAP7_75t_L g430 ( .A(n_34), .B(n_431), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_35), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_37), .B(n_117), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_38), .A2(n_81), .B1(n_126), .B2(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_39), .B(n_135), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_40), .B(n_117), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_41), .B(n_133), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_42), .A2(n_126), .B(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_43), .A2(n_50), .B1(n_759), .B2(n_760), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_43), .Y(n_760) );
AND2x2_ASAP7_75t_L g189 ( .A(n_44), .B(n_147), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_45), .B(n_133), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_46), .B(n_147), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_47), .B(n_117), .Y(n_516) );
INVx1_ASAP7_75t_L g120 ( .A(n_48), .Y(n_120) );
INVx1_ASAP7_75t_L g130 ( .A(n_48), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_49), .B(n_135), .Y(n_471) );
INVx1_ASAP7_75t_L g759 ( .A(n_50), .Y(n_759) );
AND2x2_ASAP7_75t_L g483 ( .A(n_51), .B(n_147), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_52), .B(n_117), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_53), .B(n_133), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_54), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_55), .B(n_133), .Y(n_507) );
AND2x2_ASAP7_75t_L g148 ( .A(n_56), .B(n_147), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_57), .B(n_117), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_58), .B(n_135), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_59), .B(n_117), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_60), .A2(n_126), .B(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_61), .B(n_133), .Y(n_144) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_62), .B(n_112), .Y(n_214) );
AND2x2_ASAP7_75t_L g498 ( .A(n_63), .B(n_112), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_64), .A2(n_126), .B(n_153), .Y(n_152) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_65), .A2(n_101), .B1(n_438), .B2(n_445), .C1(n_772), .C2(n_778), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_65), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_66), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_67), .B(n_162), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_68), .B(n_133), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_69), .B(n_133), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_70), .A2(n_91), .B1(n_126), .B2(n_172), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_71), .B(n_135), .Y(n_495) );
INVx1_ASAP7_75t_L g122 ( .A(n_72), .Y(n_122) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_73), .B(n_133), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_74), .A2(n_126), .B(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_75), .A2(n_126), .B(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_76), .A2(n_126), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g510 ( .A(n_77), .B(n_112), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_78), .B(n_147), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_79), .B(n_117), .Y(n_145) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_80), .A2(n_83), .B1(n_117), .B2(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g433 ( .A(n_82), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_84), .B(n_133), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_85), .B(n_133), .Y(n_199) );
AND2x2_ASAP7_75t_L g464 ( .A(n_86), .B(n_162), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_87), .A2(n_126), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_90), .B(n_135), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_92), .A2(n_126), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_93), .B(n_135), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_94), .B(n_117), .Y(n_188) );
INVxp67_ASAP7_75t_L g227 ( .A(n_95), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_96), .B(n_135), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_97), .A2(n_126), .B(n_211), .Y(n_210) );
BUFx2_ASAP7_75t_L g497 ( .A(n_98), .Y(n_497) );
BUFx2_ASAP7_75t_L g444 ( .A(n_99), .Y(n_444) );
BUFx2_ASAP7_75t_SL g782 ( .A(n_99), .Y(n_782) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_424), .B(n_434), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
XNOR2x1_ASAP7_75t_L g104 ( .A(n_105), .B(n_421), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_105), .A2(n_448), .B1(n_450), .B2(n_755), .Y(n_447) );
INVx3_ASAP7_75t_SL g762 ( .A(n_105), .Y(n_762) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_351), .Y(n_105) );
NOR4xp25_ASAP7_75t_SL g106 ( .A(n_107), .B(n_244), .C(n_288), .D(n_315), .Y(n_106) );
OAI221xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_205), .B1(n_215), .B2(n_232), .C(n_234), .Y(n_107) );
AOI32xp33_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_158), .A3(n_178), .B1(n_190), .B2(n_201), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_109), .B(n_387), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_109), .A2(n_357), .B1(n_415), .B2(n_418), .Y(n_414) );
AND2x4_ASAP7_75t_SL g109 ( .A(n_110), .B(n_138), .Y(n_109) );
INVx5_ASAP7_75t_L g204 ( .A(n_110), .Y(n_204) );
OR2x2_ASAP7_75t_L g233 ( .A(n_110), .B(n_203), .Y(n_233) );
AND2x4_ASAP7_75t_L g235 ( .A(n_110), .B(n_150), .Y(n_235) );
INVx2_ASAP7_75t_L g250 ( .A(n_110), .Y(n_250) );
OR2x2_ASAP7_75t_L g262 ( .A(n_110), .B(n_159), .Y(n_262) );
AND2x2_ASAP7_75t_L g269 ( .A(n_110), .B(n_149), .Y(n_269) );
AND2x2_ASAP7_75t_SL g311 ( .A(n_110), .B(n_192), .Y(n_311) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_110), .Y(n_368) );
OR2x6_ASAP7_75t_L g110 ( .A(n_111), .B(n_115), .Y(n_110) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_112), .Y(n_147) );
AND2x2_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x4_ASAP7_75t_L g137 ( .A(n_113), .B(n_114), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_125), .B(n_137), .Y(n_115) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_123), .Y(n_117) );
INVx1_ASAP7_75t_L g231 ( .A(n_118), .Y(n_231) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
AND2x6_ASAP7_75t_L g133 ( .A(n_119), .B(n_128), .Y(n_133) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g135 ( .A(n_121), .B(n_130), .Y(n_135) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx5_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
AND2x2_ASAP7_75t_L g129 ( .A(n_124), .B(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
AND2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
BUFx3_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
INVx2_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
AND2x4_ASAP7_75t_L g172 ( .A(n_129), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g168 ( .A(n_130), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_134), .B(n_136), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_133), .B(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_136), .A2(n_143), .B(n_144), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_136), .A2(n_154), .B(n_155), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_136), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_136), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_136), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_136), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_136), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_136), .A2(n_488), .B(n_489), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_136), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_136), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_136), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_136), .A2(n_534), .B(n_535), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_137), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_137), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_137), .B(n_227), .Y(n_226) );
NOR3xp33_ASAP7_75t_L g229 ( .A(n_137), .B(n_230), .C(n_231), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_137), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_137), .A2(n_516), .B(n_517), .Y(n_515) );
INVx3_ASAP7_75t_SL g263 ( .A(n_138), .Y(n_263) );
AND2x2_ASAP7_75t_L g282 ( .A(n_138), .B(n_204), .Y(n_282) );
AOI32xp33_ASAP7_75t_L g397 ( .A1(n_138), .A2(n_268), .A3(n_298), .B1(n_328), .B2(n_363), .Y(n_397) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_149), .Y(n_138) );
AND2x2_ASAP7_75t_L g237 ( .A(n_139), .B(n_159), .Y(n_237) );
OR2x2_ASAP7_75t_L g253 ( .A(n_139), .B(n_150), .Y(n_253) );
INVx1_ASAP7_75t_L g276 ( .A(n_139), .Y(n_276) );
INVx2_ASAP7_75t_L g292 ( .A(n_139), .Y(n_292) );
AND2x2_ASAP7_75t_L g329 ( .A(n_139), .B(n_192), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_139), .B(n_150), .Y(n_348) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_139), .Y(n_417) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_146), .B(n_148), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
AO21x2_ASAP7_75t_L g150 ( .A1(n_146), .A2(n_151), .B(n_157), .Y(n_150) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_146), .A2(n_151), .B(n_157), .Y(n_203) );
AOI21x1_ASAP7_75t_L g530 ( .A1(n_146), .A2(n_531), .B(n_537), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_147), .Y(n_146) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_147), .A2(n_196), .B(n_200), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_147), .A2(n_459), .B(n_460), .Y(n_458) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_147), .A2(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g384 ( .A(n_150), .B(n_159), .Y(n_384) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_150), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_156), .Y(n_151) );
OR2x2_ASAP7_75t_L g232 ( .A(n_158), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g238 ( .A(n_158), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g251 ( .A(n_158), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g413 ( .A(n_158), .B(n_282), .Y(n_413) );
BUFx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g342 ( .A(n_159), .B(n_292), .Y(n_342) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_160), .Y(n_192) );
AOI21x1_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_164), .B(n_177), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_162), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_162), .A2(n_492), .B(n_493), .Y(n_491) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g182 ( .A(n_163), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_165), .B(n_171), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_166), .A2(n_172), .B1(n_221), .B2(n_223), .Y(n_220) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_170), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2x1p5_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_178), .B(n_309), .Y(n_411) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_179), .B(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g194 ( .A(n_180), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g216 ( .A(n_180), .Y(n_216) );
AND2x2_ASAP7_75t_L g242 ( .A(n_180), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_180), .B(n_218), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_180), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g300 ( .A(n_180), .Y(n_300) );
OR2x2_ASAP7_75t_L g319 ( .A(n_180), .B(n_246), .Y(n_319) );
INVx1_ASAP7_75t_L g326 ( .A(n_180), .Y(n_326) );
NOR2xp33_ASAP7_75t_R g378 ( .A(n_180), .B(n_207), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_180), .B(n_219), .Y(n_382) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI21x1_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_181) );
INVx4_ASAP7_75t_L g228 ( .A(n_182), .Y(n_228) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_182), .A2(n_467), .B(n_473), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
AOI32xp33_ASAP7_75t_L g405 ( .A1(n_190), .A2(n_241), .A3(n_406), .B1(n_407), .B2(n_408), .Y(n_405) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx2_ASAP7_75t_L g272 ( .A(n_192), .Y(n_272) );
AND2x4_ASAP7_75t_L g291 ( .A(n_192), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_192), .B(n_263), .Y(n_320) );
OR2x2_ASAP7_75t_L g374 ( .A(n_192), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g332 ( .A(n_193), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g390 ( .A(n_193), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_194), .B(n_207), .Y(n_356) );
AND2x2_ASAP7_75t_L g393 ( .A(n_194), .B(n_359), .Y(n_393) );
INVx2_ASAP7_75t_L g243 ( .A(n_195), .Y(n_243) );
INVx2_ASAP7_75t_L g246 ( .A(n_195), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_195), .B(n_207), .Y(n_266) );
INVx1_ASAP7_75t_L g297 ( .A(n_195), .Y(n_297) );
OR2x2_ASAP7_75t_L g323 ( .A(n_195), .B(n_207), .Y(n_323) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_195), .Y(n_375) );
BUFx3_ASAP7_75t_L g404 ( .A(n_195), .Y(n_404) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g273 ( .A(n_202), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_202), .B(n_291), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_202), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_203), .B(n_276), .Y(n_275) );
OAI21xp33_ASAP7_75t_L g305 ( .A1(n_203), .A2(n_272), .B(n_290), .Y(n_305) );
OAI32xp33_ASAP7_75t_L g327 ( .A1(n_204), .A2(n_328), .A3(n_330), .B1(n_332), .B2(n_334), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_204), .B(n_291), .Y(n_400) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g333 ( .A(n_206), .Y(n_333) );
NOR2x1p5_ASAP7_75t_L g403 ( .A(n_206), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x4_ASAP7_75t_L g217 ( .A(n_207), .B(n_218), .Y(n_217) );
AND2x4_ASAP7_75t_SL g241 ( .A(n_207), .B(n_219), .Y(n_241) );
OR2x2_ASAP7_75t_L g245 ( .A(n_207), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g280 ( .A(n_207), .Y(n_280) );
AND2x2_ASAP7_75t_L g298 ( .A(n_207), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g309 ( .A(n_207), .B(n_219), .Y(n_309) );
OR2x2_ASAP7_75t_L g371 ( .A(n_207), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g388 ( .A(n_207), .B(n_319), .Y(n_388) );
INVx1_ASAP7_75t_L g420 ( .A(n_207), .Y(n_420) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_214), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_216), .B(n_297), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_217), .B(n_331), .Y(n_330) );
AOI222xp33_ASAP7_75t_L g335 ( .A1(n_217), .A2(n_336), .B1(n_341), .B2(n_343), .C1(n_346), .C2(n_349), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_217), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g363 ( .A(n_217), .B(n_242), .Y(n_363) );
AND2x2_ASAP7_75t_L g325 ( .A(n_218), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g340 ( .A(n_218), .B(n_245), .Y(n_340) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_219), .B(n_246), .Y(n_278) );
AND2x4_ASAP7_75t_L g299 ( .A(n_219), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g359 ( .A(n_219), .B(n_280), .Y(n_359) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_225), .Y(n_219) );
INVx3_ASAP7_75t_L g503 ( .A(n_228), .Y(n_503) );
INVx1_ASAP7_75t_SL g239 ( .A(n_233), .Y(n_239) );
NAND2xp33_ASAP7_75t_SL g408 ( .A(n_233), .B(n_263), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_238), .C(n_240), .Y(n_234) );
INVx2_ASAP7_75t_SL g285 ( .A(n_235), .Y(n_285) );
AND2x2_ASAP7_75t_L g289 ( .A(n_236), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_237), .B(n_285), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_237), .A2(n_275), .B(n_311), .C(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g387 ( .A(n_237), .B(n_368), .Y(n_387) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
AND2x4_ASAP7_75t_L g286 ( .A(n_241), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_SL g391 ( .A(n_241), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .B(n_254), .C(n_281), .Y(n_244) );
INVx2_ASAP7_75t_L g256 ( .A(n_245), .Y(n_256) );
OR2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_246), .Y(n_287) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_249), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g341 ( .A(n_249), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_249), .B(n_329), .Y(n_395) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_251), .A2(n_354), .B1(n_355), .B2(n_357), .C1(n_360), .C2(n_363), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_252), .A2(n_317), .B1(n_320), .B2(n_321), .C(n_327), .Y(n_316) );
AND2x2_ASAP7_75t_L g354 ( .A(n_252), .B(n_311), .Y(n_354) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp33_ASAP7_75t_SL g267 ( .A(n_253), .B(n_268), .Y(n_267) );
AOI221x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_259), .B1(n_264), .B2(n_267), .C(n_270), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g407 ( .A(n_257), .B(n_345), .Y(n_407) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g265 ( .A(n_258), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
OAI32xp33_ASAP7_75t_L g373 ( .A1(n_263), .A2(n_304), .A3(n_374), .B1(n_376), .B2(n_380), .Y(n_373) );
OAI21xp33_ASAP7_75t_SL g392 ( .A1(n_264), .A2(n_393), .B(n_394), .Y(n_392) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI21xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .B(n_277), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OR2x2_ASAP7_75t_L g274 ( .A(n_272), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g347 ( .A(n_272), .B(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_276), .A2(n_302), .B1(n_305), .B2(n_306), .C(n_310), .Y(n_301) );
INVx1_ASAP7_75t_L g377 ( .A(n_276), .Y(n_377) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_276), .Y(n_383) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OAI21xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_286), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_285), .B(n_350), .Y(n_349) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_293), .B(n_301), .Y(n_288) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_292), .Y(n_362) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_295), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g314 ( .A(n_297), .Y(n_314) );
INVx1_ASAP7_75t_L g304 ( .A(n_299), .Y(n_304) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_299), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_299), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_299), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g318 ( .A(n_309), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_314), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_335), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g331 ( .A(n_319), .Y(n_331) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_SL g345 ( .A(n_323), .Y(n_345) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_325), .B(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_326), .Y(n_339) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_337), .B(n_340), .Y(n_336) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g350 ( .A(n_342), .Y(n_350) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g369 ( .A(n_348), .Y(n_369) );
NOR4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_385), .C(n_396), .D(n_409), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_364), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_354), .A2(n_365), .B(n_370), .C(n_373), .Y(n_364) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_369), .Y(n_366) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_367), .A2(n_377), .B(n_378), .C(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OAI21xp33_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_383), .B(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_384), .B(n_416), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_388), .B1(n_389), .B2(n_390), .C(n_392), .Y(n_385) );
INVx1_ASAP7_75t_SL g389 ( .A(n_387), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND3xp33_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .C(n_405), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp33_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
CKINVDCx11_ASAP7_75t_R g424 ( .A(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g777 ( .A(n_427), .Y(n_777) );
BUFx2_ASAP7_75t_L g784 ( .A(n_427), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AND2x6_ASAP7_75t_SL g449 ( .A(n_428), .B(n_430), .Y(n_449) );
OR2x6_ASAP7_75t_SL g757 ( .A(n_428), .B(n_429), .Y(n_757) );
OR2x2_ASAP7_75t_L g771 ( .A(n_428), .B(n_430), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_SL g441 ( .A(n_442), .B(n_444), .Y(n_441) );
INVx2_ASAP7_75t_L g776 ( .A(n_442), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_442), .A2(n_780), .B(n_783), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_444), .B(n_776), .Y(n_775) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_758), .B1(n_761), .B2(n_766), .C(n_767), .Y(n_446) );
CKINVDCx11_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_449), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_450), .Y(n_764) );
AND2x4_ASAP7_75t_L g450 ( .A(n_451), .B(n_680), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_452), .B(n_599), .Y(n_451) );
NAND5xp2_ASAP7_75t_L g452 ( .A(n_453), .B(n_543), .C(n_553), .D(n_570), .E(n_586), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_479), .B1(n_521), .B2(n_525), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g527 ( .A(n_457), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g545 ( .A(n_457), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g566 ( .A(n_457), .B(n_567), .Y(n_566) );
INVx4_ASAP7_75t_L g580 ( .A(n_457), .Y(n_580) );
AND2x2_ASAP7_75t_L g589 ( .A(n_457), .B(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_SL g611 ( .A(n_457), .B(n_529), .Y(n_611) );
BUFx2_ASAP7_75t_L g654 ( .A(n_457), .Y(n_654) );
AND2x2_ASAP7_75t_L g669 ( .A(n_457), .B(n_466), .Y(n_669) );
OR2x2_ASAP7_75t_L g701 ( .A(n_457), .B(n_702), .Y(n_701) );
NOR4xp25_ASAP7_75t_L g750 ( .A(n_457), .B(n_751), .C(n_752), .D(n_753), .Y(n_750) );
OR2x6_ASAP7_75t_L g457 ( .A(n_458), .B(n_464), .Y(n_457) );
AOI31xp33_ASAP7_75t_L g618 ( .A1(n_465), .A2(n_619), .A3(n_621), .B(n_623), .Y(n_618) );
INVx2_ASAP7_75t_SL g735 ( .A(n_465), .Y(n_735) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_474), .Y(n_465) );
INVx2_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
AND2x2_ASAP7_75t_L g546 ( .A(n_466), .B(n_530), .Y(n_546) );
INVx2_ASAP7_75t_L g569 ( .A(n_466), .Y(n_569) );
AND2x2_ASAP7_75t_L g588 ( .A(n_466), .B(n_529), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .Y(n_467) );
AND2x2_ASAP7_75t_L g540 ( .A(n_474), .B(n_541), .Y(n_540) );
BUFx3_ASAP7_75t_L g547 ( .A(n_474), .Y(n_547) );
INVx2_ASAP7_75t_L g565 ( .A(n_474), .Y(n_565) );
AND2x2_ASAP7_75t_L g620 ( .A(n_474), .B(n_580), .Y(n_620) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AND2x4_ASAP7_75t_L g591 ( .A(n_475), .B(n_476), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_511), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_499), .Y(n_480) );
OR2x2_ASAP7_75t_L g521 ( .A(n_481), .B(n_522), .Y(n_521) );
INVx3_ASAP7_75t_L g672 ( .A(n_481), .Y(n_672) );
OR2x2_ASAP7_75t_L g720 ( .A(n_481), .B(n_721), .Y(n_720) );
NAND2x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
OR2x2_ASAP7_75t_SL g512 ( .A(n_482), .B(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g550 ( .A(n_482), .Y(n_550) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_482), .Y(n_594) );
INVx2_ASAP7_75t_L g602 ( .A(n_482), .Y(n_602) );
OR2x2_ASAP7_75t_L g637 ( .A(n_482), .B(n_501), .Y(n_637) );
AND2x2_ASAP7_75t_L g749 ( .A(n_482), .B(n_604), .Y(n_749) );
AND2x2_ASAP7_75t_L g754 ( .A(n_482), .B(n_514), .Y(n_754) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
OR2x2_ASAP7_75t_L g513 ( .A(n_490), .B(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g578 ( .A(n_490), .B(n_500), .Y(n_578) );
OR2x2_ASAP7_75t_L g585 ( .A(n_490), .B(n_550), .Y(n_585) );
NOR2x1_ASAP7_75t_SL g604 ( .A(n_490), .B(n_524), .Y(n_604) );
BUFx2_ASAP7_75t_L g636 ( .A(n_490), .Y(n_636) );
AND2x2_ASAP7_75t_L g645 ( .A(n_490), .B(n_550), .Y(n_645) );
AND2x2_ASAP7_75t_L g678 ( .A(n_490), .B(n_598), .Y(n_678) );
INVx2_ASAP7_75t_SL g687 ( .A(n_490), .Y(n_687) );
AND2x2_ASAP7_75t_L g690 ( .A(n_490), .B(n_501), .Y(n_690) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_498), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_499), .B(n_555), .C(n_640), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_499), .B(n_602), .Y(n_705) );
INVxp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_500), .B(n_687), .Y(n_708) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_501), .Y(n_552) );
AND2x2_ASAP7_75t_L g596 ( .A(n_501), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g661 ( .A(n_501), .B(n_662), .Y(n_661) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_510), .Y(n_502) );
AO21x1_ASAP7_75t_SL g524 ( .A1(n_503), .A2(n_504), .B(n_510), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
AND2x4_ASAP7_75t_L g556 ( .A(n_511), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g692 ( .A(n_513), .B(n_637), .Y(n_692) );
AND2x2_ASAP7_75t_L g523 ( .A(n_514), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
INVx2_ASAP7_75t_L g598 ( .A(n_514), .Y(n_598) );
INVx1_ASAP7_75t_L g662 ( .A(n_514), .Y(n_662) );
INVx2_ASAP7_75t_L g744 ( .A(n_521), .Y(n_744) );
OR2x2_ASAP7_75t_L g608 ( .A(n_522), .B(n_585), .Y(n_608) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g748 ( .A(n_523), .B(n_645), .Y(n_748) );
AND2x2_ASAP7_75t_L g641 ( .A(n_524), .B(n_598), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_538), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_527), .A2(n_655), .B1(n_672), .B2(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g568 ( .A(n_529), .Y(n_568) );
AND2x2_ASAP7_75t_L g622 ( .A(n_529), .B(n_542), .Y(n_622) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_529), .Y(n_649) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_530), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
INVxp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_540), .B(n_654), .Y(n_653) );
OAI32xp33_ASAP7_75t_L g670 ( .A1(n_540), .A2(n_671), .A3(n_673), .B1(n_674), .B2(n_676), .Y(n_670) );
BUFx2_ASAP7_75t_L g555 ( .A(n_541), .Y(n_555) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g697 ( .A(n_542), .B(n_591), .Y(n_697) );
OR4x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_547), .C(n_548), .D(n_551), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_544), .A2(n_635), .B1(n_729), .B2(n_730), .Y(n_728) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_545), .Y(n_737) );
AND2x2_ASAP7_75t_L g579 ( .A(n_546), .B(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g659 ( .A(n_546), .Y(n_659) );
INVx1_ASAP7_75t_L g675 ( .A(n_546), .Y(n_675) );
INVx1_ASAP7_75t_L g710 ( .A(n_546), .Y(n_710) );
OR2x2_ASAP7_75t_L g667 ( .A(n_547), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g711 ( .A(n_547), .B(n_712), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_548), .A2(n_585), .B1(n_629), .B2(n_648), .Y(n_650) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g694 ( .A(n_549), .B(n_603), .Y(n_694) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g561 ( .A(n_550), .Y(n_561) );
NOR2xp67_ASAP7_75t_L g576 ( .A(n_550), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g557 ( .A(n_551), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_551), .B(n_555), .C(n_636), .D(n_648), .Y(n_684) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g721 ( .A(n_552), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_556), .B1(n_558), .B2(n_562), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_554), .A2(n_555), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx3_ASAP7_75t_L g583 ( .A(n_560), .Y(n_583) );
AOI32xp33_ASAP7_75t_L g699 ( .A1(n_560), .A2(n_700), .A3(n_704), .B1(n_709), .B2(n_713), .Y(n_699) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g605 ( .A(n_563), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g658 ( .A(n_563), .B(n_659), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_563), .A2(n_571), .B1(n_683), .B2(n_688), .C(n_691), .Y(n_682) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g615 ( .A(n_564), .B(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g730 ( .A(n_564), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_565), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g572 ( .A(n_567), .Y(n_572) );
AND2x2_ASAP7_75t_L g590 ( .A(n_567), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_SL g630 ( .A(n_568), .Y(n_630) );
INVx1_ASAP7_75t_L g614 ( .A(n_569), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B1(n_579), .B2(n_581), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g716 ( .A(n_572), .B(n_646), .Y(n_716) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g656 ( .A(n_575), .Y(n_656) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
AND2x2_ASAP7_75t_L g587 ( .A(n_580), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_580), .B(n_617), .Y(n_616) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_580), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_580), .B(n_622), .Y(n_743) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_581), .A2(n_741), .B1(n_742), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
OR2x2_ASAP7_75t_L g623 ( .A(n_583), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g633 ( .A(n_583), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_583), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_583), .B(n_687), .Y(n_686) );
AND2x4_ASAP7_75t_SL g688 ( .A(n_583), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g664 ( .A(n_585), .B(n_665), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_589), .B(n_592), .Y(n_586) );
INVx1_ASAP7_75t_L g606 ( .A(n_588), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_589), .A2(n_626), .B1(n_633), .B2(n_638), .Y(n_625) );
INVx3_ASAP7_75t_L g628 ( .A(n_591), .Y(n_628) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
OAI32xp33_ASAP7_75t_SL g683 ( .A1(n_594), .A2(n_654), .A3(n_684), .B1(n_685), .B2(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g603 ( .A(n_597), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND4xp25_ASAP7_75t_SL g599 ( .A(n_600), .B(n_625), .C(n_642), .D(n_657), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_605), .B1(n_607), .B2(n_609), .C(n_618), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx2_ASAP7_75t_L g640 ( .A(n_602), .Y(n_640) );
AND2x2_ASAP7_75t_L g689 ( .A(n_602), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_602), .B(n_641), .Y(n_727) );
AND2x2_ASAP7_75t_L g738 ( .A(n_602), .B(n_661), .Y(n_738) );
INVx2_ASAP7_75t_L g624 ( .A(n_604), .Y(n_624) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B(n_615), .Y(n_609) );
AND2x2_ASAP7_75t_L g741 ( .A(n_610), .B(n_612), .Y(n_741) );
INVx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_611), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g718 ( .A(n_616), .Y(n_718) );
INVx1_ASAP7_75t_L g703 ( .A(n_617), .Y(n_703) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_620), .B(n_675), .Y(n_674) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_621), .B(n_628), .Y(n_632) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g731 ( .A(n_622), .Y(n_731) );
INVx1_ASAP7_75t_L g713 ( .A(n_624), .Y(n_713) );
OR2x2_ASAP7_75t_L g729 ( .A(n_624), .B(n_640), .Y(n_729) );
NAND2xp33_ASAP7_75t_SL g626 ( .A(n_627), .B(n_631), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx2_ASAP7_75t_L g646 ( .A(n_628), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_628), .B(n_641), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_628), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g725 ( .A(n_629), .Y(n_725) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_634), .A2(n_715), .B1(n_717), .B2(n_719), .Y(n_714) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g679 ( .A(n_637), .Y(n_679) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g665 ( .A(n_641), .Y(n_665) );
AOI322xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .A3(n_647), .B1(n_650), .B2(n_651), .C1(n_652), .C2(n_655), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_643), .A2(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g660 ( .A(n_645), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g717 ( .A(n_646), .B(n_718), .Y(n_717) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_653), .B(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g673 ( .A(n_654), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_654), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_663), .B2(n_666), .C(n_670), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_659), .A2(n_746), .B1(n_748), .B2(n_749), .C(n_750), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_661), .B(n_672), .Y(n_671) );
BUFx2_ASAP7_75t_L g712 ( .A(n_662), .Y(n_712) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_666), .A2(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp33_ASAP7_75t_SL g746 ( .A(n_675), .B(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NOR4xp75_ASAP7_75t_L g680 ( .A(n_681), .B(n_698), .C(n_722), .D(n_739), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_693), .Y(n_681) );
INVx1_ASAP7_75t_L g752 ( .A(n_690), .Y(n_752) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g724 ( .A(n_697), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g751 ( .A(n_697), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_699), .B(n_714), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g747 ( .A(n_718), .Y(n_747) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND3x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_732), .C(n_736), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_726), .B(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_745), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_756), .Y(n_765) );
CKINVDCx11_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g766 ( .A(n_758), .Y(n_766) );
OAI22x1_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx2_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx4f_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_777), .Y(n_773) );
INVxp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
CKINVDCx11_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
CKINVDCx8_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
endmodule