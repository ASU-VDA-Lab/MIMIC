module fake_jpeg_26342_n_246 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_40),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_16),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_23),
.Y(n_71)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_36),
.B1(n_27),
.B2(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_63),
.B1(n_66),
.B2(n_18),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_27),
.B1(n_20),
.B2(n_36),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_74),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_33),
.Y(n_102)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_29),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_76),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_39),
.A2(n_0),
.B(n_1),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_78),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_91),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_103),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_53),
.A2(n_31),
.B1(n_21),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_96),
.B1(n_64),
.B2(n_73),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_42),
.C(n_19),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_100),
.C(n_108),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_31),
.B1(n_22),
.B2(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_26),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_35),
.C(n_26),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_107),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_33),
.B1(n_29),
.B2(n_34),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_106),
.B1(n_62),
.B2(n_76),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_0),
.B(n_1),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_0),
.Y(n_108)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_13),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_2),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_108),
.C(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_118),
.B1(n_104),
.B2(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_117),
.B(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_73),
.B1(n_67),
.B2(n_60),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_127),
.B1(n_126),
.B2(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_3),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_13),
.A3(n_12),
.B1(n_11),
.B2(n_8),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_10),
.C(n_88),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_132),
.A2(n_100),
.B1(n_102),
.B2(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_5),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_10),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_139),
.B(n_149),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_161),
.B1(n_123),
.B2(n_125),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_83),
.B(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_143),
.B1(n_158),
.B2(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_147),
.Y(n_163)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_83),
.B(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_91),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_156),
.Y(n_168)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_101),
.Y(n_156)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_95),
.B1(n_89),
.B2(n_94),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_89),
.B1(n_94),
.B2(n_88),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_159),
.A2(n_131),
.B1(n_116),
.B2(n_117),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_177),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_173),
.B1(n_157),
.B2(n_160),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_170),
.B1(n_180),
.B2(n_155),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_116),
.C(n_135),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_181),
.C(n_144),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_125),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_118),
.B1(n_112),
.B2(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_10),
.B(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_159),
.B1(n_146),
.B2(n_149),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_141),
.C(n_152),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_185),
.B(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_151),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_188),
.B(n_192),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_194),
.C(n_197),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_181),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_198),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_147),
.C(n_153),
.Y(n_194)
);

OA21x2_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_148),
.B(n_145),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_SL g200 ( 
.A(n_195),
.B(n_172),
.C(n_178),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_154),
.C(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_202),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_209),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_178),
.B(n_180),
.Y(n_207)
);

HAxp5_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_191),
.CON(n_219),
.SN(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_196),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_190),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_218),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_189),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_187),
.C(n_198),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_219),
.A2(n_220),
.B1(n_209),
.B2(n_177),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_197),
.B1(n_173),
.B2(n_196),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_167),
.C(n_168),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_211),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_210),
.B(n_205),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_227),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_210),
.B(n_201),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_226),
.B(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_201),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_230),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_226),
.A2(n_162),
.B1(n_179),
.B2(n_219),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_166),
.B1(n_218),
.B2(n_225),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_162),
.B1(n_164),
.B2(n_166),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_214),
.B1(n_203),
.B2(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_232),
.B(n_231),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_217),
.Y(n_243)
);

XNOR2x2_ASAP7_75t_SL g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_208),
.Y(n_246)
);


endmodule