module real_jpeg_22219_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_0),
.A2(n_42),
.B1(n_49),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_1),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_48),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_82)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_6),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_6),
.A2(n_42),
.B1(n_49),
.B2(n_117),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_117),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_117),
.Y(n_206)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_8),
.A2(n_68),
.B1(n_69),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_8),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_42),
.B1(n_49),
.B2(n_77),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_77),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_10),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_10),
.B(n_74),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_31),
.B(n_34),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_135),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_56),
.B1(n_108),
.B2(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_10),
.B(n_89),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_10),
.A2(n_49),
.B(n_221),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_11),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_42),
.B1(n_49),
.B2(n_137),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_137),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_137),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_68),
.B1(n_69),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_13),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_42),
.B1(n_49),
.B2(n_94),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_94),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_94),
.Y(n_224)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_14),
.A2(n_30),
.A3(n_49),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_15),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_15),
.A2(n_42),
.B1(n_49),
.B2(n_70),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_208)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_97),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_22),
.B(n_97),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_79),
.B2(n_96),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_53),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_40),
.B(n_52),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_27),
.A2(n_33),
.B1(n_36),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_27),
.A2(n_33),
.B1(n_62),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_27),
.A2(n_33),
.B1(n_84),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_27),
.A2(n_33),
.B1(n_110),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_27),
.A2(n_33),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_27),
.A2(n_33),
.B1(n_186),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_27),
.A2(n_33),
.B1(n_206),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_27),
.A2(n_33),
.B1(n_128),
.B2(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_29),
.B(n_43),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_30),
.A2(n_32),
.B(n_135),
.C(n_182),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx9p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_33),
.B(n_135),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_35),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_40)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_41),
.A2(n_45),
.B1(n_87),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_41),
.A2(n_45),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_41),
.A2(n_45),
.B1(n_113),
.B2(n_132),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_41),
.A2(n_45),
.B1(n_159),
.B2(n_220),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_49),
.B1(n_72),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_42),
.A2(n_73),
.B1(n_134),
.B2(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_42),
.B(n_135),
.Y(n_217)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_49),
.B(n_72),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_61),
.B1(n_78),
.B2(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B(n_60),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_82),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_56),
.A2(n_58),
.B1(n_107),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_56),
.A2(n_57),
.B1(n_149),
.B2(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_56),
.A2(n_58),
.B1(n_175),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_56),
.A2(n_108),
.B1(n_178),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_56),
.A2(n_58),
.B1(n_164),
.B2(n_208),
.Y(n_214)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_61),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_72),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g134 ( 
.A(n_69),
.B(n_135),
.CON(n_134),
.SN(n_134)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_71),
.A2(n_74),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.C(n_90),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_81),
.B(n_83),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_88),
.A2(n_89),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_92),
.A2(n_95),
.B1(n_116),
.B2(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_104),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_102),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_104),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_111),
.C(n_114),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_105),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_109),
.Y(n_124)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_135),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_262),
.B(n_267),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_165),
.B(n_249),
.C(n_261),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_150),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_122),
.B(n_150),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_138),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_124),
.B(n_125),
.C(n_138),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_133),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_136),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_140),
.B(n_144),
.C(n_145),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_143),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_151),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.C(n_162),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_161),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_248),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_243),
.B(n_247),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_229),
.B(n_242),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_210),
.B(n_228),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_198),
.B(n_209),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_187),
.B(n_197),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_179),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_183),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_192),
.B(n_196),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_191),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_200),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_218),
.B1(n_226),
.B2(n_227),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_213),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_215),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_231),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_239),
.C(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_238),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_251),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_260),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_252),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_258),
.C(n_260),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);


endmodule