module real_jpeg_16479_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AO22x1_ASAP7_75t_SL g9 ( 
.A1(n_0),
.A2(n_1),
.B1(n_10),
.B2(n_11),
.Y(n_9)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

OA22x2_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_4),
.B1(n_11),
.B2(n_15),
.Y(n_14)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

OR2x4_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_16),
.B1(n_19),
.B2(n_25),
.C(n_30),
.Y(n_6)
);

CKINVDCx16_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

AOI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_12),
.B(n_13),
.Y(n_8)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_17),
.B(n_21),
.Y(n_20)
);

OR2x4_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_18),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_26),
.B(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);


endmodule