module fake_jpeg_2052_n_225 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_225);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_13),
.B(n_32),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_12),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_33),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_1),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_36),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_71),
.B1(n_81),
.B2(n_64),
.Y(n_95)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_72),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_99),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_104),
.B1(n_82),
.B2(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_56),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_63),
.B1(n_64),
.B2(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_80),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_119),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_88),
.B1(n_85),
.B2(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_124),
.Y(n_147)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_82),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_75),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_70),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_83),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_57),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_77),
.B1(n_85),
.B2(n_55),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_27),
.B1(n_50),
.B2(n_47),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_89),
.B1(n_68),
.B2(n_65),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_138),
.Y(n_152)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_88),
.B1(n_83),
.B2(n_97),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_137),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_58),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_62),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_61),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_110),
.B1(n_77),
.B2(n_76),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_161),
.B1(n_53),
.B2(n_23),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_155),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_151),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_68),
.B1(n_59),
.B2(n_65),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_154),
.A2(n_158),
.B1(n_171),
.B2(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_68),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_0),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_164),
.Y(n_184)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_132),
.B(n_4),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_4),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_172),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_126),
.A2(n_26),
.B1(n_46),
.B2(n_45),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_136),
.C(n_25),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_5),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_143),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_176),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_148),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_189),
.B1(n_162),
.B2(n_10),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_192),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_24),
.B(n_43),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_187),
.B1(n_18),
.B2(n_37),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_171),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_165),
.C(n_153),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_199),
.B1(n_39),
.B2(n_34),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_165),
.C(n_151),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.C(n_197),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_29),
.C(n_42),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_28),
.C(n_40),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_187),
.B1(n_181),
.B2(n_182),
.Y(n_205)
);

OAI322xp33_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_188),
.A3(n_184),
.B1(n_186),
.B2(n_176),
.C1(n_179),
.C2(n_181),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_209),
.C(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_202),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_182),
.B1(n_10),
.B2(n_11),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_30),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_209),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_35),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_31),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_213),
.B(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_7),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g218 ( 
.A1(n_215),
.A2(n_204),
.B(n_206),
.C(n_15),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_217),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_211),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_218),
.B(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_221),
.B(n_212),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_222),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_16),
.Y(n_225)
);


endmodule