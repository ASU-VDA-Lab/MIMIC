module fake_netlist_1_5876_n_455 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_455);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_455;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_123;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g69 ( .A(n_13), .Y(n_69) );
INVxp67_ASAP7_75t_SL g70 ( .A(n_53), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_35), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_64), .Y(n_72) );
CKINVDCx16_ASAP7_75t_R g73 ( .A(n_10), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_24), .Y(n_74) );
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_61), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_8), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_18), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_16), .Y(n_78) );
BUFx2_ASAP7_75t_L g79 ( .A(n_26), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_39), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
INVxp67_ASAP7_75t_L g82 ( .A(n_54), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_31), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_25), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_66), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_1), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_41), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_33), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_48), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_60), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_36), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_17), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_12), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_45), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_50), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_58), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_3), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_44), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_29), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_11), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_14), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_52), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_79), .B(n_0), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_79), .B(n_0), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_75), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_89), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_71), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_91), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_87), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_81), .B(n_1), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_93), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_91), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_90), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_99), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_71), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_90), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_72), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_72), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_98), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_86), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_73), .B(n_2), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_96), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_107), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_110), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_108), .B(n_78), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_108), .A2(n_102), .B1(n_99), .B2(n_103), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_110), .Y(n_131) );
BUFx8_ASAP7_75t_SL g132 ( .A(n_111), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_115), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_123), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_114), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_123), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_116), .B(n_96), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_114), .Y(n_139) );
INVx8_ASAP7_75t_L g140 ( .A(n_118), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_116), .B(n_101), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_109), .B(n_103), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_109), .B(n_101), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_125), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_117), .B(n_69), .Y(n_146) );
OR2x2_ASAP7_75t_L g147 ( .A(n_106), .B(n_85), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_117), .B(n_119), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_122), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_128), .Y(n_151) );
BUFx4f_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_138), .B(n_106), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_141), .B(n_119), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_131), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_144), .B(n_120), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
OAI221xp5_ASAP7_75t_L g160 ( .A1(n_147), .A2(n_124), .B1(n_121), .B2(n_120), .C(n_105), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_144), .B(n_121), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_142), .B(n_124), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_133), .B(n_113), .Y(n_163) );
NAND2xp33_ASAP7_75t_SL g164 ( .A(n_147), .B(n_145), .Y(n_164) );
NOR2xp33_ASAP7_75t_R g165 ( .A(n_127), .B(n_76), .Y(n_165) );
NOR3xp33_ASAP7_75t_SL g166 ( .A(n_130), .B(n_112), .C(n_95), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_142), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_135), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
NOR2xp33_ASAP7_75t_SL g175 ( .A(n_140), .B(n_102), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_146), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_146), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
AOI222xp33_ASAP7_75t_L g182 ( .A1(n_164), .A2(n_129), .B1(n_88), .B2(n_148), .C1(n_140), .C2(n_139), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_169), .Y(n_183) );
BUFx12f_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_153), .B(n_140), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_169), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_162), .B(n_139), .Y(n_187) );
BUFx2_ASAP7_75t_SL g188 ( .A(n_162), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_169), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_171), .B(n_149), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_152), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_172), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_152), .B(n_149), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_152), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_154), .A2(n_150), .B(n_134), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_180), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_158), .B(n_122), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_155), .B(n_126), .Y(n_201) );
BUFx2_ASAP7_75t_L g202 ( .A(n_162), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_162), .A2(n_86), .B1(n_126), .B2(n_77), .Y(n_204) );
INVx5_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_162), .B(n_126), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_161), .B(n_82), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_179), .B(n_70), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_155), .B(n_74), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_173), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_179), .B(n_100), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_172), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_190), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_205), .B(n_171), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_182), .B(n_166), .C(n_175), .Y(n_215) );
OAI21x1_ASAP7_75t_L g216 ( .A1(n_183), .A2(n_181), .B(n_178), .Y(n_216) );
OAI221xp5_ASAP7_75t_L g217 ( .A1(n_182), .A2(n_163), .B1(n_160), .B2(n_174), .C(n_170), .Y(n_217) );
NAND2xp33_ASAP7_75t_R g218 ( .A(n_190), .B(n_165), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_184), .A2(n_173), .B1(n_176), .B2(n_170), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_183), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_184), .A2(n_173), .B1(n_176), .B2(n_174), .Y(n_221) );
OR2x6_ASAP7_75t_L g222 ( .A(n_188), .B(n_184), .Y(n_222) );
NOR2x1_ASAP7_75t_SL g223 ( .A(n_188), .B(n_176), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_205), .Y(n_224) );
INVx5_ASAP7_75t_L g225 ( .A(n_190), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_205), .B(n_157), .Y(n_226) );
AOI21xp33_ASAP7_75t_L g227 ( .A1(n_206), .A2(n_177), .B(n_157), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_186), .B(n_167), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_210), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_186), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_205), .B(n_181), .Y(n_232) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_190), .A2(n_178), .B1(n_167), .B2(n_180), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_190), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_189), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_185), .B(n_177), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_189), .B(n_180), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_231), .B(n_192), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_215), .A2(n_202), .B1(n_209), .B2(n_132), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_225), .A2(n_205), .B1(n_192), .B2(n_212), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_225), .B(n_205), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_218), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_215), .A2(n_202), .B1(n_209), .B2(n_210), .Y(n_244) );
OAI211xp5_ASAP7_75t_L g245 ( .A1(n_217), .A2(n_204), .B(n_201), .C(n_207), .Y(n_245) );
AOI21xp33_ASAP7_75t_L g246 ( .A1(n_233), .A2(n_199), .B(n_201), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_212), .B1(n_197), .B2(n_187), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_235), .A2(n_210), .B1(n_203), .B2(n_200), .Y(n_248) );
OAI211xp5_ASAP7_75t_L g249 ( .A1(n_219), .A2(n_211), .B(n_208), .C(n_193), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_225), .A2(n_197), .B1(n_187), .B2(n_200), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_231), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_235), .A2(n_210), .B1(n_203), .B2(n_200), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_231), .B(n_180), .Y(n_253) );
NOR2xp67_ASAP7_75t_L g254 ( .A(n_225), .B(n_191), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_225), .B(n_198), .Y(n_255) );
AOI22xp33_ASAP7_75t_SL g256 ( .A1(n_213), .A2(n_194), .B1(n_191), .B2(n_203), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_216), .A2(n_196), .B(n_151), .Y(n_257) );
AOI33xp33_ASAP7_75t_L g258 ( .A1(n_221), .A2(n_77), .A3(n_80), .B1(n_84), .B2(n_92), .B3(n_94), .Y(n_258) );
OR2x2_ASAP7_75t_SL g259 ( .A(n_236), .B(n_86), .Y(n_259) );
NOR2xp33_ASAP7_75t_R g260 ( .A(n_251), .B(n_213), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_251), .Y(n_261) );
AND2x6_ASAP7_75t_SL g262 ( .A(n_242), .B(n_222), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_259), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_239), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_239), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_259), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_253), .B(n_236), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_253), .B(n_236), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_240), .B(n_228), .C(n_229), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_257), .A2(n_216), .B(n_220), .Y(n_270) );
OAI211xp5_ASAP7_75t_L g271 ( .A1(n_243), .A2(n_229), .B(n_237), .C(n_97), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_244), .B(n_228), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_242), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_247), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_247), .Y(n_275) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_257), .A2(n_227), .B(n_228), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g277 ( .A1(n_250), .A2(n_223), .B1(n_220), .B2(n_222), .Y(n_277) );
OAI22xp33_ASAP7_75t_L g278 ( .A1(n_250), .A2(n_222), .B1(n_237), .B2(n_230), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_242), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
INVx4_ASAP7_75t_L g281 ( .A(n_262), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_261), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_278), .A2(n_241), .B(n_246), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_266), .Y(n_285) );
OAI21xp5_ASAP7_75t_SL g286 ( .A1(n_263), .A2(n_242), .B(n_256), .Y(n_286) );
NAND5xp2_ASAP7_75t_SL g287 ( .A(n_271), .B(n_245), .C(n_249), .D(n_248), .E(n_252), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_264), .B(n_220), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
OAI22xp5_ASAP7_75t_SL g291 ( .A1(n_263), .A2(n_222), .B1(n_214), .B2(n_224), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_260), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_270), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_262), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_264), .B(n_220), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_279), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_271), .A2(n_86), .B1(n_227), .B2(n_80), .C(n_104), .Y(n_297) );
OAI211xp5_ASAP7_75t_L g298 ( .A1(n_277), .A2(n_86), .B(n_254), .C(n_83), .Y(n_298) );
OAI21xp5_ASAP7_75t_SL g299 ( .A1(n_277), .A2(n_214), .B(n_226), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_265), .B(n_267), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_275), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_267), .B(n_238), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_279), .B(n_254), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_265), .B(n_238), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_270), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_268), .B(n_230), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_270), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_276), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_285), .B(n_274), .Y(n_309) );
NAND2xp33_ASAP7_75t_SL g310 ( .A(n_281), .B(n_274), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_300), .B(n_268), .Y(n_311) );
XNOR2xp5_ASAP7_75t_L g312 ( .A(n_292), .B(n_269), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_302), .B(n_275), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_287), .A2(n_269), .B1(n_273), .B2(n_279), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_285), .B(n_279), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_283), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_288), .B(n_290), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_302), .B(n_304), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_281), .B(n_3), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_281), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_294), .A2(n_273), .B1(n_279), .B2(n_272), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_304), .Y(n_323) );
NAND2xp33_ASAP7_75t_SL g324 ( .A(n_294), .B(n_279), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_301), .B(n_276), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_291), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_306), .B(n_273), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_306), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_289), .Y(n_329) );
INVx3_ASAP7_75t_SL g330 ( .A(n_294), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_296), .B(n_276), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_296), .B(n_276), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_289), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_295), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_308), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_293), .B(n_273), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_286), .B(n_258), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_291), .B(n_280), .Y(n_339) );
OA21x2_ASAP7_75t_L g340 ( .A1(n_284), .A2(n_280), .B(n_226), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_303), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_299), .B(n_280), .Y(n_342) );
NOR2xp33_ASAP7_75t_R g343 ( .A(n_287), .B(n_4), .Y(n_343) );
NAND2x1_ASAP7_75t_SL g344 ( .A(n_330), .B(n_303), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_338), .A2(n_326), .B1(n_320), .B2(n_312), .Y(n_345) );
OAI21xp33_ASAP7_75t_SL g346 ( .A1(n_339), .A2(n_297), .B(n_305), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g347 ( .A(n_339), .B(n_298), .C(n_123), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_343), .A2(n_83), .B1(n_299), .B2(n_307), .C(n_305), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_328), .B(n_303), .Y(n_349) );
NAND4xp25_ASAP7_75t_SL g350 ( .A(n_330), .B(n_293), .C(n_5), .D(n_6), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_321), .A2(n_222), .B1(n_230), .B2(n_224), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_323), .B(n_4), .Y(n_352) );
OAI31xp33_ASAP7_75t_L g353 ( .A1(n_310), .A2(n_214), .A3(n_230), .B(n_226), .Y(n_353) );
AOI21xp33_ASAP7_75t_SL g354 ( .A1(n_322), .A2(n_5), .B(n_6), .Y(n_354) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_314), .A2(n_226), .B(n_232), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_319), .A2(n_232), .B1(n_214), .B2(n_224), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_329), .B(n_7), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_316), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_313), .B(n_7), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_324), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_311), .B(n_333), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_310), .A2(n_232), .B(n_194), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_317), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_334), .B(n_8), .Y(n_364) );
OAI321xp33_ASAP7_75t_L g365 ( .A1(n_342), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_12), .C(n_13), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_335), .B(n_9), .Y(n_366) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_318), .B(n_234), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_324), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_309), .B(n_14), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_327), .B(n_15), .Y(n_371) );
AOI32xp33_ASAP7_75t_L g372 ( .A1(n_309), .A2(n_232), .A3(n_195), .B1(n_223), .B2(n_159), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_195), .B(n_234), .C(n_198), .Y(n_373) );
OAI21xp5_ASAP7_75t_SL g374 ( .A1(n_315), .A2(n_234), .B(n_198), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_340), .A2(n_195), .B(n_198), .C(n_234), .Y(n_375) );
OAI32xp33_ASAP7_75t_L g376 ( .A1(n_325), .A2(n_159), .A3(n_151), .B1(n_20), .B2(n_21), .Y(n_376) );
NOR2xp33_ASAP7_75t_SL g377 ( .A(n_315), .B(n_234), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_315), .B(n_19), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_337), .A2(n_198), .B1(n_156), .B2(n_159), .Y(n_379) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_325), .B(n_332), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_368), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_344), .Y(n_382) );
NOR2xp67_ASAP7_75t_SL g383 ( .A(n_365), .B(n_340), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_349), .B(n_337), .Y(n_384) );
OR3x1_ASAP7_75t_L g385 ( .A(n_350), .B(n_340), .C(n_331), .Y(n_385) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_362), .B(n_336), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_361), .B(n_331), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
NOR3xp33_ASAP7_75t_SL g389 ( .A(n_346), .B(n_22), .C(n_23), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_363), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_353), .A2(n_27), .B(n_28), .C(n_32), .Y(n_391) );
NOR2xp33_ASAP7_75t_R g392 ( .A(n_367), .B(n_34), .Y(n_392) );
NOR3xp33_ASAP7_75t_SL g393 ( .A(n_365), .B(n_37), .C(n_38), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_370), .B(n_40), .Y(n_394) );
AOI21xp5_ASAP7_75t_SL g395 ( .A1(n_362), .A2(n_42), .B(n_43), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_360), .B(n_156), .Y(n_396) );
AND2x4_ASAP7_75t_SL g397 ( .A(n_357), .B(n_156), .Y(n_397) );
NAND2xp33_ASAP7_75t_SL g398 ( .A(n_378), .B(n_156), .Y(n_398) );
NOR3xp33_ASAP7_75t_SL g399 ( .A(n_348), .B(n_46), .C(n_47), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_371), .B(n_49), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_359), .B(n_51), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_352), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_360), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_369), .B(n_55), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_366), .Y(n_406) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_377), .B(n_156), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_369), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_388), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_385), .A2(n_347), .B1(n_356), .B2(n_351), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_390), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_385), .A2(n_372), .B1(n_354), .B2(n_374), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_382), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_389), .A2(n_355), .B(n_375), .C(n_373), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_393), .A2(n_376), .B(n_377), .Y(n_415) );
XNOR2xp5_ASAP7_75t_L g416 ( .A(n_401), .B(n_379), .Y(n_416) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_395), .B(n_56), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_402), .A2(n_134), .B1(n_143), .B2(n_137), .C(n_63), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_404), .A2(n_143), .B1(n_137), .B2(n_62), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_387), .B(n_57), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_381), .B(n_59), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_65), .B(n_67), .C(n_68), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_406), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_403), .Y(n_425) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_395), .B(n_396), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
AOI211xp5_ASAP7_75t_SL g428 ( .A1(n_424), .A2(n_391), .B(n_405), .C(n_400), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_426), .A2(n_391), .B(n_396), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_412), .A2(n_386), .B1(n_397), .B2(n_394), .Y(n_430) );
XNOR2xp5_ASAP7_75t_L g431 ( .A(n_416), .B(n_397), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_413), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_424), .A2(n_393), .B(n_399), .C(n_408), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_410), .A2(n_398), .B1(n_399), .B2(n_407), .Y(n_434) );
NOR2x1_ASAP7_75t_SL g435 ( .A(n_425), .B(n_392), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_425), .A2(n_427), .B1(n_409), .B2(n_411), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_415), .A2(n_414), .B1(n_417), .B2(n_422), .C(n_419), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g438 ( .A1(n_414), .A2(n_421), .B(n_419), .C(n_420), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_418), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_424), .A2(n_380), .B1(n_423), .B2(n_412), .C(n_402), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g441 ( .A1(n_424), .A2(n_345), .B1(n_380), .B2(n_410), .C(n_413), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_440), .A2(n_430), .B1(n_432), .B2(n_437), .Y(n_442) );
CKINVDCx12_ASAP7_75t_R g443 ( .A(n_431), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_439), .B(n_430), .Y(n_444) );
OR3x2_ASAP7_75t_L g445 ( .A(n_441), .B(n_435), .C(n_428), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_436), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_445), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_442), .A2(n_433), .B1(n_434), .B2(n_429), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_444), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_447), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_449), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_450), .A2(n_448), .B1(n_443), .B2(n_446), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_450), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_453), .A2(n_451), .B1(n_433), .B2(n_429), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_454), .A2(n_452), .B(n_438), .Y(n_455) );
endmodule