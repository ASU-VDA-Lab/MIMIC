module fake_jpeg_29221_n_552 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_552);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_88),
.Y(n_114)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g156 ( 
.A(n_60),
.Y(n_156)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_9),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_79),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_20),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_80),
.Y(n_122)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_9),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_29),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_105),
.Y(n_133)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_107),
.Y(n_131)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_43),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_48),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_31),
.C(n_43),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_126),
.B(n_142),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_61),
.A2(n_39),
.B1(n_34),
.B2(n_50),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_139),
.B1(n_140),
.B2(n_144),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_80),
.B(n_46),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_130),
.B(n_162),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_70),
.A2(n_39),
.B1(n_34),
.B2(n_50),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_39),
.B1(n_93),
.B2(n_83),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_57),
.A2(n_39),
.B1(n_50),
.B2(n_27),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_141),
.A2(n_28),
.B1(n_67),
.B2(n_78),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_39),
.B1(n_34),
.B2(n_27),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_53),
.A2(n_33),
.B1(n_46),
.B2(n_30),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_149),
.A2(n_170),
.B1(n_44),
.B2(n_28),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_79),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_33),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_60),
.B(n_30),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_166),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_38),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_58),
.A2(n_42),
.B1(n_36),
.B2(n_26),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_109),
.A2(n_48),
.B(n_23),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_174),
.A2(n_0),
.B(n_1),
.Y(n_237)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_176),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_102),
.B1(n_99),
.B2(n_91),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_177),
.A2(n_220),
.B1(n_230),
.B2(n_160),
.Y(n_284)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_114),
.B(n_42),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_179),
.B(n_199),
.Y(n_278)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_182),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_36),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_204),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_65),
.B1(n_64),
.B2(n_81),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_184),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_243)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_185),
.Y(n_268)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_189),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVx6_ASAP7_75t_SL g251 ( 
.A(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_196),
.Y(n_271)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_124),
.B(n_26),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_200),
.Y(n_280)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_136),
.Y(n_202)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_124),
.A2(n_27),
.A3(n_44),
.B1(n_24),
.B2(n_26),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_23),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_205),
.B(n_206),
.Y(n_260)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_224),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_210),
.Y(n_262)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_215),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_141),
.A2(n_77),
.B1(n_73),
.B2(n_90),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_128),
.A2(n_87),
.B1(n_44),
.B2(n_28),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_23),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_146),
.B(n_23),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_217),
.Y(n_282)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_139),
.A2(n_48),
.B1(n_23),
.B2(n_3),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_218),
.A2(n_221),
.B1(n_0),
.B2(n_1),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_111),
.A2(n_48),
.B1(n_10),
.B2(n_3),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_144),
.A2(n_48),
.B1(n_10),
.B2(n_4),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_123),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_222),
.Y(n_275)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_223),
.Y(n_281)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_156),
.B(n_8),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_8),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_227),
.A2(n_228),
.B1(n_231),
.B2(n_232),
.Y(n_267)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_148),
.A2(n_8),
.B1(n_16),
.B2(n_4),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_140),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_115),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

OR2x2_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_151),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_186),
.A2(n_158),
.B1(n_164),
.B2(n_167),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_245),
.A2(n_250),
.B1(n_243),
.B2(n_267),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_171),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_247),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_191),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_184),
.A2(n_173),
.B1(n_169),
.B2(n_151),
.Y(n_250)
);

MAJx3_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_283),
.C(n_208),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_171),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_257),
.B(n_259),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g258 ( 
.A(n_237),
.B(n_152),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_258),
.B(n_7),
.CI(n_12),
.CON(n_325),
.SN(n_325)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_192),
.B(n_168),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_177),
.A2(n_118),
.B1(n_168),
.B2(n_172),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_209),
.B1(n_203),
.B2(n_217),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_219),
.B(n_118),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_274),
.B(n_285),
.Y(n_302)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_230),
.B1(n_201),
.B2(n_200),
.Y(n_295)
);

OR2x4_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_116),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_284),
.A2(n_7),
.B(n_11),
.C(n_12),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_155),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_182),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_286),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_298),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_288),
.A2(n_297),
.B1(n_305),
.B2(n_313),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_251),
.A2(n_224),
.B1(n_210),
.B2(n_231),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_289),
.A2(n_317),
.B1(n_266),
.B2(n_239),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_290),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_312),
.Y(n_331)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_296),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_240),
.A2(n_228),
.B1(n_196),
.B2(n_112),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_263),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_220),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_303),
.C(n_315),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_242),
.A2(n_185),
.B(n_187),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_300),
.A2(n_304),
.B(n_264),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_208),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_301),
.B(n_314),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_190),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_240),
.A2(n_258),
.B1(n_243),
.B2(n_270),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_260),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_309),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_307),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_319),
.B1(n_323),
.B2(n_251),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_240),
.B(n_235),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_258),
.A2(n_195),
.B1(n_194),
.B2(n_202),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_275),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_113),
.C(n_0),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_325),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_276),
.A2(n_113),
.B1(n_5),
.B2(n_6),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_249),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_241),
.B(n_4),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_324),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_259),
.B(n_5),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_264),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_322),
.A2(n_238),
.B1(n_268),
.B2(n_269),
.Y(n_340)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_249),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_241),
.B(n_7),
.C(n_11),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_312),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_328),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_278),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_335),
.Y(n_367)
);

AO21x1_ASAP7_75t_L g386 ( 
.A1(n_334),
.A2(n_280),
.B(n_271),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_281),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_283),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_315),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_244),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_344),
.C(n_354),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_304),
.A2(n_264),
.B(n_277),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_339),
.A2(n_347),
.B(n_307),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_340),
.A2(n_311),
.B1(n_310),
.B2(n_312),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_304),
.A2(n_239),
.B(n_252),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_342),
.A2(n_355),
.B(n_14),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_343),
.A2(n_297),
.B1(n_288),
.B2(n_313),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_244),
.C(n_252),
.Y(n_344)
);

AOI32xp33_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_268),
.A3(n_272),
.B1(n_253),
.B2(n_261),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_272),
.C(n_261),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_300),
.A2(n_273),
.B(n_253),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_273),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_301),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_362),
.A2(n_374),
.B1(n_375),
.B2(n_346),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_363),
.A2(n_377),
.B(n_383),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_287),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_364),
.B(n_380),
.Y(n_405)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_366),
.A2(n_371),
.B1(n_373),
.B2(n_389),
.Y(n_410)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_384),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_376),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_331),
.A2(n_295),
.B1(n_305),
.B2(n_317),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_324),
.C(n_325),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_385),
.C(n_387),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_331),
.A2(n_295),
.B1(n_293),
.B2(n_322),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_330),
.A2(n_295),
.B1(n_322),
.B2(n_325),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_343),
.A2(n_322),
.B1(n_266),
.B2(n_316),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_331),
.A2(n_255),
.B(n_254),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_351),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_378),
.Y(n_400)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

NAND3xp33_ASAP7_75t_SL g380 ( 
.A(n_334),
.B(n_255),
.C(n_254),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_359),
.Y(n_381)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_381),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_351),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_382),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_290),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_338),
.B(n_280),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_388),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_271),
.C(n_308),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_328),
.B(n_12),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_392),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_350),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_391),
.A2(n_327),
.B1(n_345),
.B2(n_352),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_16),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_335),
.Y(n_395)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_419),
.Y(n_438)
);

XNOR2x1_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_339),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_397),
.B(n_423),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_336),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_399),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_401),
.A2(n_403),
.B1(n_413),
.B2(n_414),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_337),
.B1(n_333),
.B2(n_346),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_349),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_406),
.B(n_407),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_360),
.B(n_354),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_333),
.B1(n_346),
.B2(n_347),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_376),
.A2(n_341),
.B1(n_329),
.B2(n_348),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_358),
.C(n_357),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_369),
.C(n_385),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_383),
.A2(n_341),
.B1(n_329),
.B2(n_348),
.Y(n_418)
);

INVx13_ASAP7_75t_L g426 ( 
.A(n_418),
.Y(n_426)
);

NAND3xp33_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_352),
.C(n_358),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_420),
.B(n_422),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_345),
.Y(n_421)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_421),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_367),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_361),
.B(n_17),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_402),
.Y(n_457)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_427),
.Y(n_455)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_421),
.Y(n_431)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_373),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_432),
.Y(n_452)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_434),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_395),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_400),
.B(n_388),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_442),
.Y(n_465)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_393),
.B(n_390),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_440),
.B(n_411),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_387),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_409),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_445),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_408),
.B(n_363),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_393),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_447),
.Y(n_463)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_448),
.B(n_449),
.Y(n_459)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_412),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_450),
.A2(n_451),
.B1(n_416),
.B2(n_365),
.Y(n_454)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_402),
.C(n_404),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_460),
.C(n_461),
.Y(n_482)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_462),
.Y(n_475)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_458),
.B(n_466),
.CI(n_411),
.CON(n_481),
.SN(n_481)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_404),
.C(n_415),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_397),
.C(n_423),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_417),
.Y(n_462)
);

XNOR2x2_ASAP7_75t_SL g466 ( 
.A(n_440),
.B(n_394),
.Y(n_466)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_428),
.B(n_403),
.CI(n_413),
.CON(n_470),
.SN(n_470)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_470),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_417),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_472),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_401),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_410),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_371),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_410),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_438),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_468),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_487),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_484),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_492),
.Y(n_500)
);

BUFx5_ASAP7_75t_L g483 ( 
.A(n_455),
.Y(n_483)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_483),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g485 ( 
.A1(n_455),
.A2(n_427),
.B1(n_449),
.B2(n_452),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_431),
.C(n_430),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_490),
.C(n_479),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_473),
.A2(n_425),
.B1(n_436),
.B2(n_429),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_474),
.A2(n_446),
.B1(n_434),
.B2(n_429),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_488),
.A2(n_464),
.B1(n_463),
.B2(n_459),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_466),
.A2(n_430),
.B(n_396),
.C(n_433),
.Y(n_489)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_489),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_426),
.C(n_451),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_419),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_491),
.B(n_471),
.Y(n_494)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_499),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_496),
.B(n_488),
.Y(n_511)
);

OAI21xp33_ASAP7_75t_L g497 ( 
.A1(n_477),
.A2(n_458),
.B(n_467),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_497),
.A2(n_484),
.B(n_481),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_480),
.A2(n_472),
.B1(n_462),
.B2(n_470),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_505),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_460),
.C(n_470),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_507),
.C(n_482),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_483),
.B(n_469),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_508),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_476),
.A2(n_426),
.B1(n_411),
.B2(n_392),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_475),
.B(n_461),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_479),
.B(n_475),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_490),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_518),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_512),
.Y(n_528)
);

XOR2x1_ASAP7_75t_SL g513 ( 
.A(n_495),
.B(n_489),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_513),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_514),
.A2(n_496),
.B(n_502),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_482),
.C(n_481),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_515),
.B(n_516),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_504),
.A2(n_450),
.B(n_439),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_448),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_520),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_372),
.C(n_447),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_500),
.A2(n_443),
.B1(n_444),
.B2(n_379),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_522),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_386),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_513),
.A2(n_498),
.B1(n_505),
.B2(n_493),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_523),
.B(n_528),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_527),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_502),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_511),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_444),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_389),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_529),
.B(n_516),
.Y(n_534)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_534),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_530),
.B(n_368),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_536),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_524),
.A2(n_514),
.B(n_512),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_539),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_528),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_540),
.B(n_533),
.C(n_525),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_541),
.B(n_537),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_544),
.A2(n_545),
.B(n_543),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_546),
.A2(n_547),
.B(n_527),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_531),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_540),
.B(n_542),
.Y(n_549)
);

MAJx2_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_526),
.C(n_381),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_392),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_391),
.Y(n_552)
);


endmodule