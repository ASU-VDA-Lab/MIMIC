module fake_netlist_6_2369_n_1985 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1985);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1985;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_48),
.Y(n_193)
);

INVx4_ASAP7_75t_R g194 ( 
.A(n_34),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_44),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_35),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_49),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_43),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_61),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_13),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_134),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_86),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_26),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_24),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_173),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_132),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_22),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_5),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_37),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_139),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_95),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_14),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_75),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_63),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_48),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_146),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_74),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_123),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_30),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_107),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_88),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_114),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_142),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_20),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_144),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_89),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_110),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_97),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_151),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_12),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_45),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_155),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_147),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_116),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_32),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_133),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_28),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_56),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_186),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_115),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_96),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_58),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_94),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_106),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_5),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_56),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_69),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_113),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_41),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_67),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_71),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_125),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_34),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_190),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_87),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_7),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_162),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_69),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_172),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_76),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_183),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_73),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_18),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_154),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_128),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_145),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_7),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_120),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_82),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_62),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_189),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_41),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_38),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_148),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_168),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_156),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_20),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_14),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_92),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_51),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_30),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_188),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_105),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_90),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_141),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_99),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_138),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_80),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_61),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_117),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_63),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_129),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_191),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_16),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_50),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_79),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_149),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_85),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_70),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_25),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_18),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_121),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_35),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_26),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_10),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_10),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_135),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_157),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_55),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_21),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_136),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_182),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_27),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_37),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_15),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_179),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_49),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_2),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_46),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_150),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_185),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_50),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_6),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_124),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_164),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_51),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_140),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_15),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_111),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_171),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_27),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_24),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_36),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_31),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_38),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_161),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_169),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_143),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_137),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_78),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_130),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_174),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_19),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_8),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_187),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_33),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_12),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_29),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_81),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_52),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_21),
.Y(n_373)
);

BUFx8_ASAP7_75t_SL g374 ( 
.A(n_52),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_23),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_16),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_104),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_25),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_68),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_131),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_102),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_108),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_31),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_160),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_240),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_374),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_281),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_217),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_352),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_199),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_288),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_318),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_245),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_275),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_193),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_234),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_236),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_238),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_289),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_197),
.B(n_308),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_289),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_289),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_199),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_289),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_239),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_241),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_242),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_200),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_200),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_197),
.B(n_0),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_359),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_289),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_308),
.B(n_0),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_251),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_360),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_254),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_382),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_311),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_311),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_311),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_332),
.B(n_1),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_311),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_215),
.B(n_2),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_272),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_311),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_192),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_367),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_256),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_215),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_266),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_231),
.Y(n_440)
);

BUFx6f_ASAP7_75t_SL g441 ( 
.A(n_268),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_266),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_345),
.B(n_3),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_332),
.B(n_3),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_258),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_207),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_198),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_265),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_269),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_206),
.B(n_4),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_221),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_224),
.B(n_4),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_237),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_252),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_271),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_263),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_264),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_270),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_274),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_278),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_276),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_283),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_282),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_230),
.B(n_6),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_292),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_284),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_212),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_287),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_295),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_302),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_303),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_212),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_231),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_297),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_305),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_306),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_300),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_307),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_207),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_321),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_322),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_280),
.B(n_371),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_196),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_440),
.B(n_474),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_408),
.B(n_196),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_421),
.B(n_255),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_421),
.B(n_255),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_408),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_401),
.A2(n_201),
.B(n_195),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_385),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_431),
.B(n_294),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_431),
.B(n_294),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_436),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_385),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_390),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_402),
.A2(n_232),
.B1(n_356),
.B2(n_339),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_390),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_396),
.B(n_203),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_411),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_417),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_397),
.B(n_205),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_435),
.B(n_192),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_428),
.B(n_429),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_428),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_429),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_399),
.B(n_210),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_418),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_400),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_434),
.B(n_202),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_447),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_400),
.B(n_220),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_407),
.B(n_222),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_457),
.B(n_235),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_457),
.B(n_243),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_435),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_422),
.B(n_202),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_444),
.B(n_209),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_480),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_439),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_430),
.B(n_192),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_442),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g543 ( 
.A(n_387),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_473),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_432),
.B(n_192),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_412),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_446),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_446),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_448),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_448),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_483),
.B(n_209),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_452),
.B(n_246),
.Y(n_553)
);

OR2x2_ASAP7_75t_SL g554 ( 
.A(n_395),
.B(n_419),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_482),
.B(n_481),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_452),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_454),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_454),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_455),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_455),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_458),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_458),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_459),
.A2(n_248),
.B(n_247),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_530),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_485),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_500),
.A2(n_468),
.B1(n_441),
.B2(n_395),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_531),
.B(n_532),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_488),
.Y(n_568)
);

NOR2x1p5_ASAP7_75t_L g569 ( 
.A(n_552),
.B(n_391),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_552),
.B(n_433),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_503),
.B(n_465),
.C(n_453),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_530),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_486),
.Y(n_574)
);

AND2x2_ASAP7_75t_SL g575 ( 
.A(n_541),
.B(n_192),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_522),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_500),
.A2(n_441),
.B1(n_211),
.B2(n_334),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_486),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_514),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_514),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_485),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_514),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_534),
.B(n_404),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_514),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_543),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_503),
.B(n_204),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_514),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_534),
.B(n_433),
.Y(n_592)
);

NOR2x1p5_ASAP7_75t_L g593 ( 
.A(n_535),
.B(n_344),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_496),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_493),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_522),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_493),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_488),
.B(n_249),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_503),
.B(n_519),
.C(n_512),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_488),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_493),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_493),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_498),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_535),
.B(n_405),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_496),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_498),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_498),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_498),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_484),
.B(n_406),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_484),
.B(n_414),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_499),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_499),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_499),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_488),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_499),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_501),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_547),
.Y(n_618)
);

AND3x2_ASAP7_75t_L g619 ( 
.A(n_544),
.B(n_412),
.C(n_547),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_501),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_501),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_506),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_522),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_501),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_505),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_522),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_489),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_543),
.B(n_451),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_541),
.B(n_415),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_416),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_505),
.Y(n_631)
);

INVx4_ASAP7_75t_SL g632 ( 
.A(n_541),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_522),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_522),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_522),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_554),
.A2(n_479),
.B1(n_477),
.B2(n_437),
.Y(n_636)
);

INVx6_ASAP7_75t_L g637 ( 
.A(n_495),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_505),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_545),
.Y(n_640)
);

AND2x6_ASAP7_75t_L g641 ( 
.A(n_503),
.B(n_204),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_521),
.B(n_423),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_489),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_522),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_512),
.B(n_527),
.C(n_519),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_541),
.B(n_489),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_489),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_516),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_544),
.B(n_425),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_544),
.B(n_445),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_522),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_533),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_543),
.B(n_259),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_543),
.B(n_260),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_531),
.B(n_482),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_494),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_547),
.B(n_449),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_516),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g659 ( 
.A(n_506),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_487),
.B(n_450),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_502),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_533),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_SL g663 ( 
.A1(n_500),
.A2(n_441),
.B1(n_394),
.B2(n_386),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_516),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_496),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_520),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_520),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_541),
.A2(n_443),
.B1(n_432),
.B2(n_392),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_487),
.B(n_456),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_533),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_512),
.A2(n_443),
.B1(n_325),
.B2(n_326),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_524),
.B(n_460),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_502),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_524),
.B(n_461),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_509),
.B(n_463),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_520),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_509),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_545),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_525),
.B(n_467),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_494),
.B(n_469),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_520),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_494),
.B(n_471),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_494),
.B(n_476),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_512),
.B(n_312),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_495),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_525),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_523),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_495),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_531),
.B(n_532),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_SL g692 ( 
.A(n_538),
.B(n_470),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_523),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_523),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_538),
.B(n_472),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_490),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_506),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_554),
.B(n_403),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_545),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_533),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_560),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_495),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_533),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_554),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_519),
.B(n_268),
.Y(n_706)
);

AO22x2_ASAP7_75t_L g707 ( 
.A1(n_545),
.A2(n_378),
.B1(n_335),
.B2(n_353),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_490),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_490),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_519),
.B(n_462),
.C(n_459),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_560),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_495),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_553),
.A2(n_227),
.B1(n_226),
.B2(n_216),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_527),
.B(n_464),
.C(n_462),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_565),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_568),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_618),
.B(n_560),
.Y(n_717)
);

NOR2x1p5_ASAP7_75t_L g718 ( 
.A(n_682),
.B(n_208),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_599),
.B(n_527),
.Y(n_719)
);

BUFx8_ASAP7_75t_L g720 ( 
.A(n_675),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_599),
.B(n_645),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_572),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_568),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_615),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_571),
.B(n_560),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_574),
.B(n_527),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_615),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_575),
.A2(n_528),
.B1(n_563),
.B2(n_553),
.Y(n_728)
);

INVx8_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_579),
.B(n_528),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_572),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_574),
.B(n_528),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_586),
.B(n_528),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_600),
.B(n_561),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_575),
.A2(n_563),
.B1(n_553),
.B2(n_375),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_600),
.B(n_627),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_627),
.B(n_561),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_571),
.B(n_561),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_588),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_605),
.A2(n_563),
.B(n_491),
.C(n_553),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_628),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_647),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_645),
.B(n_204),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_575),
.A2(n_563),
.B1(n_366),
.B2(n_491),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_618),
.Y(n_745)
);

BUFx6f_ASAP7_75t_SL g746 ( 
.A(n_688),
.Y(n_746)
);

AND2x4_ASAP7_75t_SL g747 ( 
.A(n_688),
.B(n_388),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_584),
.Y(n_748)
);

BUFx5_ASAP7_75t_L g749 ( 
.A(n_595),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_647),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_687),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_643),
.B(n_561),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_699),
.B(n_532),
.C(n_531),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_643),
.B(n_545),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_656),
.B(n_555),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_688),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_687),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_640),
.B(n_204),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_584),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_656),
.B(n_610),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_590),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_690),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_611),
.B(n_545),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_690),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_590),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_660),
.B(n_545),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_671),
.B(n_532),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_630),
.B(n_250),
.C(n_244),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_602),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_688),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_676),
.B(n_495),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_653),
.B(n_555),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_629),
.A2(n_420),
.B1(n_424),
.B2(n_426),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_567),
.B(n_495),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_567),
.B(n_492),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_691),
.B(n_492),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_691),
.B(n_492),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_702),
.B(n_497),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_702),
.B(n_497),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_711),
.B(n_497),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_711),
.B(n_504),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_679),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_679),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_684),
.B(n_213),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_675),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_686),
.B(n_504),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_707),
.A2(n_491),
.B1(n_559),
.B2(n_558),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_703),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_602),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_685),
.B(n_213),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_640),
.B(n_204),
.Y(n_791)
);

CKINVDCx11_ASAP7_75t_R g792 ( 
.A(n_594),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_640),
.B(n_290),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_703),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_649),
.B(n_393),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_593),
.B(n_507),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_655),
.B(n_555),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_580),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_570),
.B(n_214),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_603),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_666),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_650),
.B(n_214),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_680),
.B(n_290),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_655),
.B(n_555),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_569),
.B(n_313),
.Y(n_805)
);

BUFx5_ASAP7_75t_L g806 ( 
.A(n_595),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_603),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_653),
.B(n_464),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_661),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_581),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_607),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_607),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_592),
.B(n_218),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_593),
.B(n_507),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_582),
.B(n_508),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_582),
.B(n_508),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_585),
.B(n_508),
.Y(n_817)
);

BUFx5_ASAP7_75t_L g818 ( 
.A(n_597),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_608),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_674),
.B(n_218),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_637),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_587),
.B(n_510),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_608),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_569),
.A2(n_398),
.B1(n_298),
.B2(n_293),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_637),
.Y(n_825)
);

BUFx10_ASAP7_75t_L g826 ( 
.A(n_619),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_707),
.A2(n_491),
.B1(n_559),
.B2(n_558),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_587),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_713),
.B(n_550),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_680),
.B(n_290),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_653),
.B(n_466),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_591),
.B(n_510),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_609),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_710),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_646),
.A2(n_515),
.B(n_511),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_564),
.B(n_573),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_700),
.B(n_290),
.Y(n_837)
);

NAND2x1p5_ASAP7_75t_L g838 ( 
.A(n_700),
.B(n_261),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_606),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_L g840 ( 
.A(n_670),
.B(n_257),
.C(n_253),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_583),
.B(n_290),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_653),
.B(n_466),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_564),
.B(n_510),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_573),
.B(n_511),
.Y(n_844)
);

INVx8_ASAP7_75t_L g845 ( 
.A(n_628),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_583),
.B(n_279),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_609),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_583),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_577),
.B(n_511),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_712),
.A2(n_285),
.B1(n_304),
.B2(n_323),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_577),
.B(n_513),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_707),
.A2(n_562),
.B1(n_559),
.B2(n_558),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_632),
.B(n_328),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_642),
.B(n_219),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_705),
.B(n_219),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_705),
.B(n_223),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_637),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_632),
.B(n_363),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_606),
.B(n_550),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_598),
.B(n_513),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_612),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_636),
.B(n_556),
.Y(n_862)
);

INVx8_ASAP7_75t_L g863 ( 
.A(n_628),
.Y(n_863)
);

INVx8_ASAP7_75t_L g864 ( 
.A(n_628),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_712),
.A2(n_515),
.B(n_533),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_637),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_598),
.B(n_513),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_598),
.B(n_622),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_612),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_710),
.A2(n_562),
.B(n_556),
.C(n_557),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_614),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_598),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_657),
.B(n_223),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_697),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_659),
.B(n_517),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_677),
.B(n_225),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_698),
.B(n_517),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_760),
.B(n_566),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_745),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_733),
.B(n_706),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_798),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_766),
.A2(n_623),
.B(n_576),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_724),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_733),
.B(n_673),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_763),
.A2(n_623),
.B(n_576),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_730),
.A2(n_623),
.B(n_576),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_771),
.A2(n_623),
.B(n_576),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_724),
.B(n_653),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_742),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_742),
.B(n_654),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_726),
.B(n_732),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_782),
.B(n_663),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_726),
.B(n_708),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_782),
.B(n_692),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_732),
.B(n_708),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_810),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_729),
.B(n_654),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_767),
.B(n_709),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_821),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_802),
.A2(n_681),
.B1(n_696),
.B2(n_654),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_736),
.B(n_709),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_802),
.A2(n_714),
.B(n_377),
.C(n_380),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_755),
.B(n_597),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_755),
.B(n_604),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_721),
.A2(n_714),
.B(n_616),
.C(n_613),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_721),
.A2(n_707),
.B1(n_589),
.B2(n_641),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_783),
.B(n_578),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_821),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_740),
.A2(n_613),
.B(n_604),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_745),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_754),
.A2(n_634),
.B(n_633),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_735),
.A2(n_654),
.B1(n_365),
.B2(n_357),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_784),
.B(n_616),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_784),
.B(n_625),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_790),
.B(n_625),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_719),
.A2(n_634),
.B(n_633),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_790),
.B(n_638),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_834),
.B(n_638),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_735),
.A2(n_834),
.B1(n_728),
.B2(n_744),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_719),
.A2(n_634),
.B(n_633),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_774),
.A2(n_669),
.B(n_634),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_797),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_725),
.B(n_648),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_743),
.A2(n_668),
.B(n_658),
.C(n_648),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_797),
.B(n_658),
.Y(n_925)
);

NAND2x1_ASAP7_75t_L g926 ( 
.A(n_848),
.B(n_669),
.Y(n_926)
);

INVx1_ASAP7_75t_SL g927 ( 
.A(n_785),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_804),
.B(n_668),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_859),
.B(n_654),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_828),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_839),
.B(n_225),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_804),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_717),
.B(n_212),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_801),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_716),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_740),
.A2(n_694),
.B(n_689),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_762),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_723),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_738),
.B(n_689),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_809),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_868),
.A2(n_669),
.B(n_596),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_728),
.A2(n_368),
.B1(n_341),
.B2(n_348),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_727),
.B(n_632),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_872),
.A2(n_632),
.B1(n_589),
.B2(n_641),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_773),
.B(n_556),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_786),
.B(n_694),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_743),
.A2(n_669),
.B(n_596),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_753),
.A2(n_757),
.B1(n_764),
.B2(n_751),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_750),
.B(n_734),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_737),
.B(n_614),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_752),
.A2(n_596),
.B(n_704),
.Y(n_951)
);

OAI321xp33_ASAP7_75t_L g952 ( 
.A1(n_799),
.A2(n_478),
.A3(n_475),
.B1(n_481),
.B2(n_562),
.C(n_194),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_775),
.B(n_617),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_776),
.B(n_617),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_718),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_744),
.A2(n_621),
.B(n_620),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_777),
.B(n_620),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_862),
.B(n_228),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_795),
.B(n_475),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_855),
.B(n_228),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_792),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_729),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_855),
.B(n_229),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_L g964 ( 
.A(n_876),
.B(n_233),
.C(n_229),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_796),
.B(n_621),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_814),
.B(n_624),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_SL g967 ( 
.A1(n_758),
.A2(n_639),
.B(n_624),
.C(n_695),
.Y(n_967)
);

AOI21xp33_ASAP7_75t_L g968 ( 
.A1(n_820),
.A2(n_639),
.B(n_631),
.Y(n_968)
);

AOI21xp33_ASAP7_75t_L g969 ( 
.A1(n_820),
.A2(n_664),
.B(n_631),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_758),
.A2(n_665),
.B(n_664),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_720),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_829),
.B(n_601),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_835),
.A2(n_667),
.B(n_665),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_860),
.A2(n_596),
.B(n_704),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_788),
.A2(n_794),
.B1(n_805),
.B2(n_762),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_867),
.A2(n_626),
.B(n_601),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_856),
.B(n_478),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_865),
.A2(n_704),
.B(n_635),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_854),
.B(n_233),
.Y(n_979)
);

AOI21xp33_ASAP7_75t_L g980 ( 
.A1(n_799),
.A2(n_813),
.B(n_854),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_848),
.A2(n_701),
.B(n_635),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_836),
.A2(n_683),
.B(n_678),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_874),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_825),
.B(n_626),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_825),
.A2(n_701),
.B(n_635),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_852),
.B(n_678),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_815),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_720),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_857),
.A2(n_701),
.B(n_644),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_852),
.B(n_683),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_756),
.B(n_342),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_813),
.B(n_693),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_787),
.A2(n_827),
.B1(n_840),
.B2(n_873),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_856),
.B(n_342),
.Y(n_994)
);

INVx11_ASAP7_75t_L g995 ( 
.A(n_746),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_770),
.B(n_343),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_715),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_873),
.B(n_343),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_876),
.A2(n_693),
.B(n_695),
.C(n_672),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_857),
.A2(n_672),
.B(n_644),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_816),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_875),
.B(n_626),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_729),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_768),
.B(n_346),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_866),
.A2(n_651),
.B(n_644),
.Y(n_1005)
);

AO21x1_ASAP7_75t_L g1006 ( 
.A1(n_838),
.A2(n_518),
.B(n_517),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_L g1007 ( 
.A(n_808),
.B(n_651),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_741),
.B(n_551),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_877),
.B(n_651),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_L g1010 ( 
.A(n_741),
.B(n_589),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_870),
.A2(n_518),
.B(n_529),
.C(n_551),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_787),
.A2(n_662),
.B(n_652),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_866),
.A2(n_672),
.B(n_662),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_747),
.B(n_824),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_850),
.A2(n_518),
.B(n_529),
.C(n_551),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_791),
.A2(n_662),
.B(n_652),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_747),
.B(n_551),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_808),
.B(n_548),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_791),
.A2(n_652),
.B(n_533),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_808),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_846),
.A2(n_641),
.B1(n_589),
.B2(n_557),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_749),
.B(n_589),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_749),
.B(n_589),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_817),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_769),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_793),
.A2(n_533),
.B(n_526),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_822),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_793),
.A2(n_533),
.B(n_526),
.Y(n_1028)
);

NOR2xp67_ASAP7_75t_L g1029 ( 
.A(n_739),
.B(n_789),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_SL g1030 ( 
.A1(n_803),
.A2(n_529),
.B(n_548),
.C(n_557),
.Y(n_1030)
);

AOI33xp33_ASAP7_75t_L g1031 ( 
.A1(n_827),
.A2(n_548),
.A3(n_557),
.B1(n_208),
.B2(n_369),
.B3(n_348),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_845),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_722),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_838),
.B(n_346),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_832),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_803),
.A2(n_539),
.B(n_542),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_843),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_831),
.B(n_347),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_749),
.B(n_347),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_846),
.A2(n_364),
.B(n_362),
.C(n_361),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_831),
.B(n_349),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_806),
.B(n_818),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_830),
.A2(n_837),
.B(n_841),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_806),
.B(n_349),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_844),
.A2(n_364),
.B(n_362),
.C(n_361),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_778),
.A2(n_641),
.B(n_539),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_831),
.A2(n_365),
.B1(n_357),
.B2(n_355),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_826),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_806),
.B(n_818),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_806),
.B(n_641),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_842),
.B(n_216),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_842),
.B(n_358),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_842),
.A2(n_226),
.B1(n_227),
.B2(n_340),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_806),
.B(n_358),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_772),
.A2(n_316),
.B1(n_317),
.B2(n_320),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1042),
.A2(n_837),
.B(n_830),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_980),
.A2(n_963),
.B(n_994),
.C(n_960),
.Y(n_1057)
);

OAI22x1_ASAP7_75t_L g1058 ( 
.A1(n_900),
.A2(n_907),
.B1(n_892),
.B2(n_878),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1042),
.A2(n_841),
.B(n_853),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_882),
.A2(n_858),
.B(n_853),
.Y(n_1060)
);

AND2x4_ASAP7_75t_SL g1061 ( 
.A(n_1003),
.B(n_826),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_910),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_980),
.A2(n_845),
.B(n_864),
.C(n_863),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_879),
.B(n_934),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_962),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_922),
.B(n_863),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_922),
.B(n_863),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_962),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_922),
.B(n_864),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_885),
.A2(n_858),
.B(n_780),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_902),
.A2(n_781),
.B(n_779),
.C(n_849),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_887),
.A2(n_1049),
.B(n_898),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_880),
.A2(n_851),
.B(n_772),
.C(n_800),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_927),
.B(n_746),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_932),
.B(n_864),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_993),
.A2(n_772),
.B1(n_806),
.B2(n_818),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_891),
.B(n_818),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_886),
.A2(n_871),
.B(n_869),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_930),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_940),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_L g1081 ( 
.A1(n_894),
.A2(n_340),
.B1(n_341),
.B2(n_383),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_943),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_987),
.B(n_818),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_SL g1084 ( 
.A1(n_1004),
.A2(n_861),
.B(n_847),
.C(n_833),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_983),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_881),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_1003),
.B(n_962),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1001),
.B(n_818),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_932),
.B(n_807),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1024),
.B(n_1027),
.Y(n_1090)
);

AOI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_884),
.A2(n_823),
.B(n_819),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_964),
.A2(n_350),
.B1(n_354),
.B2(n_383),
.C(n_355),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1043),
.A2(n_919),
.B(n_921),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1035),
.B(n_811),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_959),
.B(n_262),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_919),
.A2(n_946),
.B(n_895),
.Y(n_1096)
);

BUFx8_ASAP7_75t_SL g1097 ( 
.A(n_961),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_932),
.B(n_812),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_977),
.B(n_731),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_929),
.B(n_889),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_993),
.A2(n_765),
.B(n_761),
.C(n_759),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1037),
.A2(n_748),
.B(n_384),
.C(n_381),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_1048),
.B(n_329),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_972),
.A2(n_333),
.B1(n_338),
.B2(n_337),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_SL g1105 ( 
.A1(n_955),
.A2(n_1020),
.B1(n_971),
.B2(n_988),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_893),
.A2(n_895),
.B(n_913),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_889),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_893),
.A2(n_506),
.B(n_526),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_889),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_896),
.B(n_384),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1017),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_998),
.A2(n_542),
.B(n_539),
.C(n_506),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_933),
.B(n_267),
.Y(n_1113)
);

AOI33xp33_ASAP7_75t_L g1114 ( 
.A1(n_1014),
.A2(n_379),
.A3(n_369),
.B1(n_368),
.B2(n_354),
.B3(n_350),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_914),
.A2(n_330),
.B1(n_296),
.B2(n_299),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_979),
.A2(n_542),
.B(n_539),
.C(n_526),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_931),
.B(n_273),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_915),
.A2(n_506),
.B(n_526),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1032),
.B(n_542),
.Y(n_1119)
);

OAI21xp33_ASAP7_75t_SL g1120 ( 
.A1(n_1012),
.A2(n_268),
.B(n_310),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_925),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_1032),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_949),
.B(n_277),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_918),
.B(n_286),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1031),
.A2(n_336),
.B(n_301),
.C(n_309),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_1038),
.B(n_373),
.C(n_314),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_917),
.A2(n_526),
.B(n_546),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_992),
.A2(n_954),
.B(n_953),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_SL g1129 ( 
.A(n_1032),
.B(n_379),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_945),
.B(n_291),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_901),
.B(n_372),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_888),
.B(n_91),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_957),
.A2(n_549),
.B(n_546),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_911),
.A2(n_549),
.B(n_546),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_888),
.B(n_310),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1025),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_928),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_972),
.A2(n_310),
.B1(n_331),
.B2(n_327),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_956),
.A2(n_549),
.B(n_546),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_956),
.A2(n_549),
.B(n_546),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_972),
.A2(n_912),
.B1(n_938),
.B2(n_1018),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1051),
.B(n_315),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_L g1143 ( 
.A(n_1041),
.B(n_376),
.C(n_324),
.Y(n_1143)
);

NOR3xp33_ASAP7_75t_L g1144 ( 
.A(n_1052),
.B(n_319),
.C(n_9),
.Y(n_1144)
);

CKINVDCx6p67_ASAP7_75t_R g1145 ( 
.A(n_897),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_883),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_916),
.A2(n_549),
.B(n_546),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1025),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_890),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_912),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1045),
.A2(n_11),
.B(n_13),
.C(n_17),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_920),
.A2(n_549),
.B(n_546),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_890),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1018),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_972),
.A2(n_546),
.B1(n_540),
.B2(n_537),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_935),
.B(n_549),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_883),
.Y(n_1157)
);

NAND2xp33_ASAP7_75t_L g1158 ( 
.A(n_1007),
.B(n_549),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_905),
.A2(n_549),
.B(n_546),
.C(n_540),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_958),
.B(n_23),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_SL g1161 ( 
.A(n_1055),
.B(n_32),
.C(n_33),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1047),
.B(n_36),
.C(n_39),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_903),
.B(n_549),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_997),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_942),
.B(n_546),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_986),
.A2(n_540),
.B1(n_537),
.B2(n_536),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_937),
.B(n_540),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_904),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_937),
.B(n_540),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1002),
.A2(n_540),
.B(n_537),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_943),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1033),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_948),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_899),
.B(n_540),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1029),
.Y(n_1175)
);

OR2x6_ASAP7_75t_SL g1176 ( 
.A(n_942),
.B(n_1047),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1008),
.Y(n_1177)
);

AO22x1_ASAP7_75t_L g1178 ( 
.A1(n_1053),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_995),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_899),
.B(n_540),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_908),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_908),
.B(n_540),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_965),
.B(n_540),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_984),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1009),
.A2(n_537),
.B(n_536),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1034),
.A2(n_1054),
.B1(n_1039),
.B2(n_1044),
.Y(n_1186)
);

INVx8_ASAP7_75t_L g1187 ( 
.A(n_1008),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_991),
.A2(n_536),
.B1(n_537),
.B2(n_184),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_926),
.B(n_537),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_966),
.B(n_537),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_990),
.B(n_537),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_SL g1192 ( 
.A(n_996),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_950),
.B(n_537),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_923),
.B(n_975),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_952),
.A2(n_119),
.B(n_100),
.C(n_167),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1053),
.B(n_537),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_984),
.Y(n_1197)
);

OAI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1040),
.A2(n_536),
.B(n_43),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_978),
.A2(n_536),
.B(n_166),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1011),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_906),
.A2(n_536),
.B1(n_159),
.B2(n_158),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_939),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_909),
.B(n_40),
.C(n_44),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1022),
.B(n_536),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1050),
.B(n_536),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1108),
.A2(n_970),
.B(n_1036),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1108),
.A2(n_909),
.B(n_936),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1122),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1134),
.A2(n_936),
.B(n_976),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1095),
.B(n_1130),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1093),
.A2(n_999),
.B(n_973),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1057),
.A2(n_973),
.B(n_969),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1139),
.A2(n_1140),
.B(n_1170),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1072),
.A2(n_1010),
.B(n_1023),
.Y(n_1214)
);

AOI221xp5_ASAP7_75t_L g1215 ( 
.A1(n_1058),
.A2(n_969),
.B1(n_968),
.B2(n_1015),
.C(n_1030),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1139),
.A2(n_1016),
.B(n_982),
.Y(n_1216)
);

BUFx4f_ASAP7_75t_SL g1217 ( 
.A(n_1107),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1090),
.B(n_982),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1117),
.A2(n_968),
.B(n_967),
.C(n_924),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1079),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1085),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1140),
.A2(n_941),
.B(n_951),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1170),
.A2(n_974),
.B(n_1019),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_1125),
.A2(n_1063),
.B(n_1102),
.C(n_1083),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1176),
.A2(n_944),
.B1(n_1046),
.B2(n_1012),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1072),
.A2(n_1046),
.B(n_947),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1080),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1128),
.A2(n_981),
.B(n_1000),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1143),
.A2(n_984),
.B1(n_1021),
.B2(n_1005),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1185),
.A2(n_1013),
.B(n_989),
.Y(n_1230)
);

BUFx8_ASAP7_75t_L g1231 ( 
.A(n_1154),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1128),
.A2(n_985),
.B(n_1026),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1185),
.A2(n_1028),
.B(n_984),
.Y(n_1233)
);

CKINVDCx8_ASAP7_75t_R g1234 ( 
.A(n_1179),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1160),
.A2(n_984),
.B(n_536),
.C(n_53),
.Y(n_1235)
);

NAND3x1_ASAP7_75t_L g1236 ( 
.A(n_1144),
.B(n_46),
.C(n_47),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1164),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1078),
.A2(n_122),
.B(n_118),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1106),
.A2(n_536),
.B(n_112),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1096),
.A2(n_103),
.B(n_101),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1120),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1106),
.A2(n_98),
.B(n_57),
.Y(n_1242)
);

NOR2x1_ASAP7_75t_R g1243 ( 
.A(n_1065),
.B(n_54),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1172),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1147),
.A2(n_57),
.B(n_58),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1184),
.B(n_59),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1062),
.B(n_59),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1093),
.A2(n_60),
.B(n_62),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1064),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1070),
.A2(n_60),
.B(n_64),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1147),
.A2(n_64),
.B(n_65),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1184),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1152),
.A2(n_1070),
.B(n_1060),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1109),
.Y(n_1254)
);

AND2x6_ASAP7_75t_L g1255 ( 
.A(n_1132),
.B(n_65),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1168),
.B(n_68),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1065),
.Y(n_1257)
);

AO32x2_ASAP7_75t_L g1258 ( 
.A1(n_1201),
.A2(n_66),
.A3(n_67),
.B1(n_1166),
.B2(n_1115),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1161),
.A2(n_66),
.B1(n_1173),
.B2(n_1203),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1152),
.A2(n_1060),
.B(n_1133),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1094),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1097),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1192),
.A2(n_1092),
.B1(n_1142),
.B2(n_1111),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1136),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1157),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1077),
.A2(n_1056),
.B(n_1059),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1148),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1175),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1056),
.A2(n_1059),
.B(n_1194),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1159),
.A2(n_1199),
.A3(n_1101),
.B(n_1200),
.Y(n_1270)
);

AOI211x1_ASAP7_75t_L g1271 ( 
.A1(n_1178),
.A2(n_1198),
.B(n_1137),
.C(n_1121),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1133),
.A2(n_1118),
.B(n_1127),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1073),
.A2(n_1071),
.B(n_1088),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1124),
.B(n_1123),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1150),
.A2(n_1151),
.B(n_1135),
.C(n_1162),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1118),
.A2(n_1127),
.B(n_1199),
.Y(n_1276)
);

AOI221x1_ASAP7_75t_L g1277 ( 
.A1(n_1081),
.A2(n_1153),
.B1(n_1091),
.B2(n_1126),
.C(n_1196),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1131),
.A2(n_1113),
.B(n_1100),
.C(n_1110),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1149),
.B(n_1132),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1186),
.A2(n_1202),
.B(n_1138),
.C(n_1188),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1099),
.A2(n_1076),
.B(n_1190),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1184),
.A2(n_1183),
.B(n_1193),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1068),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1114),
.B(n_1149),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1184),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1156),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1141),
.B(n_1181),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1191),
.A2(n_1163),
.B(n_1189),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1181),
.B(n_1171),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1158),
.A2(n_1084),
.B(n_1204),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1068),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1165),
.A2(n_1145),
.B1(n_1177),
.B2(n_1187),
.Y(n_1292)
);

INVxp67_ASAP7_75t_SL g1293 ( 
.A(n_1082),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1068),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1082),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1187),
.A2(n_1177),
.B1(n_1066),
.B2(n_1067),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1171),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1205),
.A2(n_1174),
.B(n_1180),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1155),
.A2(n_1169),
.B(n_1167),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1177),
.Y(n_1300)
);

AO31x2_ASAP7_75t_L g1301 ( 
.A1(n_1146),
.A2(n_1116),
.A3(n_1112),
.B(n_1074),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1119),
.B(n_1087),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1182),
.A2(n_1098),
.B(n_1089),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1119),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1069),
.A2(n_1075),
.B(n_1187),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1189),
.A2(n_1104),
.B(n_1103),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1146),
.A2(n_1105),
.B1(n_1061),
.B2(n_1129),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1065),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1108),
.A2(n_1134),
.B(n_1139),
.Y(n_1309)
);

AOI31xp67_ASAP7_75t_L g1310 ( 
.A1(n_1194),
.A2(n_913),
.A3(n_915),
.B(n_914),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1057),
.A2(n_919),
.B1(n_1176),
.B2(n_1090),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1086),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1159),
.A2(n_1057),
.A3(n_1006),
.B(n_1093),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1090),
.B(n_891),
.Y(n_1314)
);

BUFx4_ASAP7_75t_SL g1315 ( 
.A(n_1122),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1057),
.B(n_386),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1090),
.B(n_891),
.Y(n_1317)
);

AO22x2_ASAP7_75t_L g1318 ( 
.A1(n_1161),
.A2(n_919),
.B1(n_993),
.B2(n_912),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1090),
.B(n_891),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1072),
.A2(n_1042),
.B(n_1057),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1072),
.A2(n_1042),
.B(n_1057),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1108),
.A2(n_1134),
.B(n_1139),
.Y(n_1322)
);

OAI22x1_ASAP7_75t_L g1323 ( 
.A1(n_1117),
.A2(n_900),
.B1(n_1130),
.B2(n_878),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1090),
.B(n_891),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_SL g1325 ( 
.A1(n_1057),
.A2(n_980),
.B(n_919),
.C(n_1195),
.Y(n_1325)
);

INVx5_ASAP7_75t_L g1326 ( 
.A(n_1184),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1087),
.B(n_1149),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_SL g1328 ( 
.A(n_1184),
.B(n_745),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1108),
.A2(n_1134),
.B(n_1139),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1072),
.A2(n_1042),
.B(n_1057),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1117),
.A2(n_795),
.B1(n_963),
.B2(n_960),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1108),
.A2(n_1134),
.B(n_1139),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1090),
.B(n_891),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1072),
.A2(n_1042),
.B(n_1128),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1086),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1057),
.B(n_386),
.Y(n_1336)
);

OAI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1176),
.A2(n_900),
.B1(n_606),
.B2(n_980),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1086),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1159),
.A2(n_1057),
.A3(n_1006),
.B(n_1093),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1095),
.B(n_959),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1062),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1197),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_SL g1343 ( 
.A1(n_1150),
.A2(n_1151),
.B(n_1006),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1057),
.A2(n_980),
.B(n_733),
.C(n_963),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1057),
.B(n_839),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1072),
.A2(n_1042),
.B(n_1057),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1072),
.A2(n_1042),
.B(n_1057),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_1074),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1057),
.A2(n_980),
.B1(n_1058),
.B2(n_1198),
.C(n_1093),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1117),
.A2(n_980),
.B1(n_960),
.B2(n_963),
.Y(n_1350)
);

BUFx10_ASAP7_75t_L g1351 ( 
.A(n_1074),
.Y(n_1351)
);

NOR2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1179),
.B(n_961),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1086),
.Y(n_1353)
);

INVx3_ASAP7_75t_SL g1354 ( 
.A(n_1179),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1057),
.A2(n_1096),
.B(n_1093),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1057),
.A2(n_980),
.B(n_733),
.C(n_963),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1331),
.A2(n_1350),
.B1(n_1314),
.B2(n_1317),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1318),
.A2(n_1336),
.B1(n_1316),
.B2(n_1323),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1262),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1312),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1327),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1327),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1353),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1257),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1337),
.A2(n_1318),
.B1(n_1311),
.B2(n_1210),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1311),
.A2(n_1259),
.B1(n_1248),
.B2(n_1345),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1231),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1259),
.A2(n_1248),
.B1(n_1340),
.B2(n_1274),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1246),
.A2(n_1314),
.B1(n_1317),
.B2(n_1319),
.Y(n_1369)
);

OAI21xp33_ASAP7_75t_L g1370 ( 
.A1(n_1344),
.A2(n_1356),
.B(n_1324),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1263),
.A2(n_1284),
.B1(n_1255),
.B2(n_1355),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1231),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1255),
.A2(n_1355),
.B1(n_1246),
.B2(n_1324),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1319),
.B(n_1333),
.Y(n_1374)
);

BUFx4f_ASAP7_75t_SL g1375 ( 
.A(n_1354),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1352),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1333),
.A2(n_1256),
.B1(n_1349),
.B2(n_1277),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1315),
.Y(n_1378)
);

BUFx8_ASAP7_75t_SL g1379 ( 
.A(n_1208),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1234),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1237),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1255),
.A2(n_1247),
.B1(n_1212),
.B2(n_1343),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1255),
.A2(n_1212),
.B1(n_1250),
.B2(n_1261),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1250),
.A2(n_1225),
.B1(n_1256),
.B2(n_1242),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1227),
.Y(n_1385)
);

INVx4_ASAP7_75t_SL g1386 ( 
.A(n_1301),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1348),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1236),
.A2(n_1249),
.B1(n_1243),
.B2(n_1258),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1348),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1258),
.A2(n_1292),
.B1(n_1335),
.B2(n_1338),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1268),
.A2(n_1296),
.B1(n_1265),
.B2(n_1279),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1254),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1220),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1257),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1341),
.A2(n_1287),
.B1(n_1304),
.B2(n_1292),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1257),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1258),
.A2(n_1265),
.B1(n_1307),
.B2(n_1351),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1291),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1351),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1326),
.B(n_1328),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1283),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1300),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1221),
.B(n_1302),
.Y(n_1403)
);

BUFx4_ASAP7_75t_R g1404 ( 
.A(n_1295),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1218),
.A2(n_1244),
.B1(n_1302),
.B2(n_1286),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1264),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1278),
.B(n_1271),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1267),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1294),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1275),
.B(n_1280),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1291),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1307),
.A2(n_1326),
.B1(n_1251),
.B2(n_1245),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1291),
.Y(n_1413)
);

INVx8_ASAP7_75t_L g1414 ( 
.A(n_1326),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1297),
.Y(n_1415)
);

INVx8_ASAP7_75t_L g1416 ( 
.A(n_1326),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1289),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1289),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1320),
.A2(n_1347),
.B1(n_1330),
.B2(n_1346),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1308),
.Y(n_1420)
);

BUFx2_ASAP7_75t_R g1421 ( 
.A(n_1252),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1293),
.Y(n_1422)
);

BUFx8_ASAP7_75t_SL g1423 ( 
.A(n_1308),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1215),
.A2(n_1281),
.B1(n_1269),
.B2(n_1347),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1342),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1215),
.A2(n_1281),
.B1(n_1346),
.B2(n_1321),
.Y(n_1426)
);

INVx6_ASAP7_75t_L g1427 ( 
.A(n_1305),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1320),
.A2(n_1321),
.B1(n_1330),
.B2(n_1207),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1229),
.A2(n_1239),
.B1(n_1303),
.B2(n_1299),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1273),
.A2(n_1303),
.B1(n_1298),
.B2(n_1285),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1235),
.A2(n_1241),
.B1(n_1273),
.B2(n_1285),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1299),
.A2(n_1306),
.B1(n_1290),
.B2(n_1211),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1211),
.A2(n_1266),
.B1(n_1226),
.B2(n_1334),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1325),
.B(n_1339),
.Y(n_1434)
);

CKINVDCx8_ASAP7_75t_R g1435 ( 
.A(n_1224),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1226),
.A2(n_1209),
.B1(n_1213),
.B2(n_1290),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1270),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1219),
.A2(n_1282),
.B1(n_1214),
.B2(n_1228),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1309),
.A2(n_1332),
.B1(n_1329),
.B2(n_1322),
.Y(n_1439)
);

INVx6_ASAP7_75t_L g1440 ( 
.A(n_1301),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1313),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1313),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1339),
.B(n_1301),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1339),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1270),
.Y(n_1445)
);

BUFx10_ASAP7_75t_L g1446 ( 
.A(n_1240),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1238),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1253),
.A2(n_1216),
.B1(n_1260),
.B2(n_1276),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1272),
.A2(n_1232),
.B1(n_1288),
.B2(n_1222),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1310),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1230),
.A2(n_1233),
.B1(n_1223),
.B2(n_1206),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1327),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1312),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1314),
.B(n_1317),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1340),
.B(n_1210),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1350),
.A2(n_980),
.B1(n_1318),
.B2(n_1331),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1340),
.B(n_1210),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1350),
.A2(n_980),
.B1(n_1318),
.B2(n_1331),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_1207),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1217),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1217),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1350),
.A2(n_980),
.B1(n_1318),
.B2(n_1331),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1312),
.Y(n_1463)
);

BUFx12f_ASAP7_75t_L g1464 ( 
.A(n_1262),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1331),
.A2(n_1350),
.B1(n_1057),
.B2(n_802),
.Y(n_1465)
);

INVx6_ASAP7_75t_L g1466 ( 
.A(n_1231),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1312),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1246),
.A2(n_1336),
.B1(n_1316),
.B2(n_919),
.Y(n_1468)
);

BUFx4f_ASAP7_75t_SL g1469 ( 
.A(n_1354),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1327),
.B(n_1087),
.Y(n_1470)
);

CKINVDCx6p67_ASAP7_75t_R g1471 ( 
.A(n_1354),
.Y(n_1471)
);

BUFx10_ASAP7_75t_L g1472 ( 
.A(n_1262),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1350),
.A2(n_980),
.B1(n_1318),
.B2(n_1331),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1246),
.A2(n_1336),
.B1(n_1316),
.B2(n_919),
.Y(n_1475)
);

CKINVDCx11_ASAP7_75t_R g1476 ( 
.A(n_1234),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1249),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1246),
.A2(n_1336),
.B1(n_1316),
.B2(n_919),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1312),
.Y(n_1479)
);

INVx4_ASAP7_75t_L g1480 ( 
.A(n_1217),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1327),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1331),
.A2(n_1350),
.B1(n_1316),
.B2(n_1336),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1331),
.A2(n_1246),
.B1(n_1176),
.B2(n_919),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1340),
.B(n_1210),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1312),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1331),
.A2(n_1350),
.B1(n_1057),
.B2(n_802),
.Y(n_1486)
);

INVx3_ASAP7_75t_SL g1487 ( 
.A(n_1354),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1217),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1327),
.Y(n_1489)
);

BUFx10_ASAP7_75t_L g1490 ( 
.A(n_1262),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1312),
.Y(n_1491)
);

CKINVDCx6p67_ASAP7_75t_R g1492 ( 
.A(n_1354),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1350),
.A2(n_980),
.B1(n_1336),
.B2(n_1316),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1314),
.B(n_1317),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1246),
.A2(n_1336),
.B1(n_1316),
.B2(n_919),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1331),
.A2(n_1246),
.B1(n_1176),
.B2(n_919),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1350),
.A2(n_980),
.B1(n_1336),
.B2(n_1316),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1312),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1417),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1418),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1414),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1414),
.B(n_1416),
.Y(n_1502)
);

AO21x1_ASAP7_75t_SL g1503 ( 
.A1(n_1373),
.A2(n_1383),
.B(n_1410),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1477),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1465),
.A2(n_1486),
.B(n_1482),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1414),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1365),
.B(n_1443),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1476),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1455),
.Y(n_1509)
);

OAI21xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1373),
.A2(n_1497),
.B(n_1493),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1441),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1359),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1442),
.B(n_1444),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1451),
.A2(n_1438),
.B(n_1439),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1403),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1437),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1423),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1445),
.B(n_1434),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1374),
.B(n_1454),
.Y(n_1519)
);

BUFx8_ASAP7_75t_L g1520 ( 
.A(n_1464),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1416),
.B(n_1427),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1416),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1363),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1445),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1468),
.A2(n_1475),
.B1(n_1478),
.B2(n_1495),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1451),
.A2(n_1439),
.B(n_1449),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1401),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1459),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1459),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1450),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1393),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1453),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1440),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1463),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1467),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1440),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1427),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1386),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1479),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1435),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1485),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1408),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1411),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1386),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1447),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1390),
.B(n_1358),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1498),
.Y(n_1548)
);

AO31x2_ASAP7_75t_L g1549 ( 
.A1(n_1431),
.A2(n_1407),
.A3(n_1357),
.B(n_1386),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1360),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1468),
.A2(n_1495),
.B(n_1478),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1491),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1422),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1381),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1406),
.Y(n_1555)
);

AO21x2_ASAP7_75t_L g1556 ( 
.A1(n_1430),
.A2(n_1377),
.B(n_1405),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1394),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1457),
.B(n_1484),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1425),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1415),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1394),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1400),
.B(n_1447),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1377),
.A2(n_1405),
.B(n_1496),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1494),
.B(n_1368),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1390),
.B(n_1358),
.Y(n_1565)
);

AND2x4_ASAP7_75t_SL g1566 ( 
.A(n_1471),
.B(n_1492),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1391),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1447),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1428),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1428),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1392),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1419),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1370),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1369),
.A2(n_1475),
.B1(n_1466),
.B2(n_1367),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1397),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1397),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1447),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1446),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1395),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1367),
.A2(n_1466),
.B1(n_1372),
.B2(n_1388),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1400),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1366),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1446),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1364),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1364),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1489),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1483),
.A2(n_1496),
.B1(n_1456),
.B2(n_1458),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1364),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1489),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1483),
.A2(n_1462),
.B1(n_1458),
.B2(n_1473),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1364),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1394),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1456),
.B(n_1462),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1426),
.B(n_1424),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1473),
.B(n_1426),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1383),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1452),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1452),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1449),
.A2(n_1433),
.B(n_1436),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1404),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1371),
.B(n_1382),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1396),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1385),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1402),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1433),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1448),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1448),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1432),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1409),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1396),
.Y(n_1614)
);

OAI222xp33_ASAP7_75t_L g1615 ( 
.A1(n_1412),
.A2(n_1399),
.B1(n_1429),
.B2(n_1375),
.C1(n_1469),
.C2(n_1378),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1412),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1474),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1470),
.A2(n_1481),
.B(n_1420),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1367),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1541),
.B(n_1487),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1515),
.B(n_1487),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1505),
.A2(n_1470),
.B(n_1481),
.C(n_1488),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1553),
.B(n_1481),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1588),
.A2(n_1421),
.B1(n_1466),
.B2(n_1372),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1510),
.A2(n_1461),
.B(n_1380),
.C(n_1387),
.Y(n_1625)
);

AOI221x1_ASAP7_75t_SL g1626 ( 
.A1(n_1576),
.A2(n_1372),
.B1(n_1389),
.B2(n_1379),
.C(n_1376),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1551),
.A2(n_1375),
.B(n_1469),
.C(n_1490),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_SL g1628 ( 
.A1(n_1579),
.A2(n_1396),
.B(n_1398),
.C(n_1413),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1553),
.B(n_1460),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_R g1630 ( 
.A(n_1508),
.B(n_1472),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1570),
.B(n_1480),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1509),
.B(n_1398),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1525),
.A2(n_1472),
.B1(n_1490),
.B2(n_1398),
.Y(n_1633)
);

O2A1O1Ixp33_ASAP7_75t_SL g1634 ( 
.A1(n_1615),
.A2(n_1602),
.B(n_1601),
.C(n_1567),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1558),
.B(n_1507),
.Y(n_1635)
);

AO21x1_ASAP7_75t_L g1636 ( 
.A1(n_1610),
.A2(n_1583),
.B(n_1574),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1591),
.A2(n_1610),
.B1(n_1607),
.B2(n_1594),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1607),
.A2(n_1594),
.B(n_1575),
.C(n_1596),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1547),
.A2(n_1565),
.B1(n_1574),
.B2(n_1577),
.C(n_1616),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1541),
.B(n_1604),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1541),
.B(n_1606),
.Y(n_1641)
);

AOI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1565),
.A2(n_1564),
.B(n_1596),
.C(n_1580),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1582),
.B(n_1534),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1595),
.A2(n_1581),
.B(n_1597),
.C(n_1616),
.Y(n_1644)
);

OA21x2_ASAP7_75t_L g1645 ( 
.A1(n_1600),
.A2(n_1514),
.B(n_1526),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1571),
.B(n_1518),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_SL g1647 ( 
.A(n_1619),
.B(n_1501),
.Y(n_1647)
);

NAND2x1_ASAP7_75t_L g1648 ( 
.A(n_1521),
.B(n_1538),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1617),
.B(n_1599),
.Y(n_1649)
);

AND2x6_ASAP7_75t_L g1650 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1519),
.A2(n_1504),
.B1(n_1605),
.B2(n_1500),
.Y(n_1651)
);

AND2x4_ASAP7_75t_SL g1652 ( 
.A(n_1512),
.B(n_1613),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1563),
.A2(n_1556),
.B1(n_1612),
.B2(n_1608),
.C(n_1573),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1573),
.A2(n_1612),
.B(n_1514),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1500),
.B(n_1499),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_SL g1656 ( 
.A(n_1503),
.B(n_1521),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1600),
.A2(n_1579),
.B(n_1584),
.Y(n_1657)
);

AOI22x1_ASAP7_75t_SL g1658 ( 
.A1(n_1508),
.A2(n_1619),
.B1(n_1512),
.B2(n_1539),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1572),
.A2(n_1619),
.B1(n_1527),
.B2(n_1606),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1499),
.B(n_1533),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1526),
.A2(n_1611),
.B(n_1609),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1513),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1549),
.B(n_1533),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1538),
.A2(n_1611),
.B(n_1609),
.C(n_1503),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1584),
.A2(n_1618),
.B(n_1590),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1537),
.B(n_1545),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1535),
.B(n_1536),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1549),
.B(n_1535),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1572),
.A2(n_1544),
.B(n_1566),
.C(n_1563),
.Y(n_1669)
);

AO32x2_ASAP7_75t_L g1670 ( 
.A1(n_1557),
.A2(n_1593),
.A3(n_1603),
.B1(n_1561),
.B2(n_1522),
.Y(n_1670)
);

AO21x1_ASAP7_75t_L g1671 ( 
.A1(n_1523),
.A2(n_1542),
.B(n_1592),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1527),
.B(n_1566),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1587),
.A2(n_1590),
.B(n_1555),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1531),
.A2(n_1530),
.B(n_1528),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1536),
.B(n_1540),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1531),
.A2(n_1530),
.B(n_1524),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1524),
.A2(n_1511),
.B(n_1516),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1614),
.B(n_1517),
.Y(n_1678)
);

NAND2x1_ASAP7_75t_L g1679 ( 
.A(n_1521),
.B(n_1562),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1563),
.A2(n_1556),
.B1(n_1548),
.B2(n_1552),
.C(n_1560),
.Y(n_1680)
);

INVxp67_ASAP7_75t_L g1681 ( 
.A(n_1614),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1517),
.B(n_1529),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1544),
.Y(n_1683)
);

AO32x2_ASAP7_75t_L g1684 ( 
.A1(n_1557),
.A2(n_1593),
.A3(n_1603),
.B1(n_1561),
.B2(n_1522),
.Y(n_1684)
);

OAI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1532),
.A2(n_1543),
.B(n_1550),
.C(n_1559),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1529),
.A2(n_1568),
.B1(n_1521),
.B2(n_1587),
.Y(n_1686)
);

NAND2x1_ASAP7_75t_L g1687 ( 
.A(n_1562),
.B(n_1502),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1661),
.B(n_1645),
.Y(n_1688)
);

NOR2xp67_ASAP7_75t_L g1689 ( 
.A(n_1685),
.B(n_1546),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.B(n_1646),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1677),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1677),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1654),
.B(n_1549),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1663),
.B(n_1668),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1674),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1676),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1676),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1687),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1653),
.B(n_1549),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1679),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1651),
.B(n_1662),
.Y(n_1701)
);

NOR3xp33_ASAP7_75t_L g1702 ( 
.A(n_1624),
.B(n_1501),
.C(n_1598),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1657),
.B(n_1578),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1621),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1650),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1671),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1631),
.B(n_1586),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1667),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1657),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1675),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1629),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1650),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1670),
.Y(n_1713)
);

NOR2x1_ASAP7_75t_SL g1714 ( 
.A(n_1623),
.B(n_1562),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1670),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1684),
.B(n_1569),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1680),
.B(n_1550),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1546),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1660),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1704),
.B(n_1620),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1720),
.B(n_1636),
.Y(n_1722)
);

OAI31xp33_ASAP7_75t_SL g1723 ( 
.A1(n_1693),
.A2(n_1639),
.A3(n_1659),
.B(n_1642),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1690),
.B(n_1635),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1696),
.Y(n_1725)
);

AO21x2_ASAP7_75t_L g1726 ( 
.A1(n_1706),
.A2(n_1669),
.B(n_1665),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1713),
.B(n_1649),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1691),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1711),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_L g1730 ( 
.A1(n_1699),
.A2(n_1642),
.B(n_1638),
.C(n_1637),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1713),
.B(n_1715),
.Y(n_1731)
);

OAI31xp33_ASAP7_75t_L g1732 ( 
.A1(n_1699),
.A2(n_1634),
.A3(n_1644),
.B(n_1627),
.Y(n_1732)
);

AOI33xp33_ASAP7_75t_L g1733 ( 
.A1(n_1706),
.A2(n_1637),
.A3(n_1633),
.B1(n_1625),
.B2(n_1652),
.B3(n_1632),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1689),
.A2(n_1664),
.B(n_1622),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1696),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1693),
.A2(n_1626),
.B1(n_1641),
.B2(n_1640),
.C(n_1665),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1702),
.A2(n_1626),
.B1(n_1648),
.B2(n_1686),
.C(n_1630),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1691),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1697),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1692),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1705),
.B(n_1712),
.Y(n_1741)
);

OAI33xp33_ASAP7_75t_L g1742 ( 
.A1(n_1718),
.A2(n_1655),
.A3(n_1681),
.B1(n_1589),
.B2(n_1585),
.B3(n_1554),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1702),
.A2(n_1568),
.B1(n_1666),
.B2(n_1643),
.Y(n_1743)
);

INVx4_ASAP7_75t_L g1744 ( 
.A(n_1705),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1717),
.B(n_1656),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1705),
.Y(n_1746)
);

INVx5_ASAP7_75t_SL g1747 ( 
.A(n_1703),
.Y(n_1747)
);

CKINVDCx9p33_ASAP7_75t_R g1748 ( 
.A(n_1707),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1692),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1704),
.B(n_1682),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1720),
.B(n_1673),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1717),
.B(n_1719),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1701),
.B(n_1673),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1700),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1700),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1716),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1700),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1700),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1745),
.B(n_1752),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1725),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1728),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1729),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1725),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1735),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1735),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1724),
.B(n_1690),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1745),
.B(n_1714),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1756),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1722),
.B(n_1701),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1745),
.B(n_1714),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1756),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1739),
.Y(n_1773)
);

NOR2xp67_ASAP7_75t_L g1774 ( 
.A(n_1722),
.B(n_1709),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.Y(n_1775)
);

NAND4xp25_ASAP7_75t_L g1776 ( 
.A(n_1723),
.B(n_1732),
.C(n_1730),
.D(n_1736),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1752),
.B(n_1700),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1752),
.B(n_1709),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1753),
.B(n_1694),
.Y(n_1780)
);

NAND2x1_ASAP7_75t_L g1781 ( 
.A(n_1754),
.B(n_1716),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1753),
.B(n_1708),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1751),
.B(n_1694),
.Y(n_1783)
);

OR2x6_ASAP7_75t_L g1784 ( 
.A(n_1744),
.B(n_1746),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1726),
.B(n_1689),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1751),
.B(n_1731),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1741),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1729),
.B(n_1711),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1731),
.B(n_1708),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1740),
.A2(n_1695),
.B(n_1688),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1731),
.B(n_1710),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1747),
.B(n_1698),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_1727),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1738),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1760),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1760),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1759),
.B(n_1747),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1761),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1762),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1774),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1776),
.B(n_1723),
.C(n_1732),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1759),
.B(n_1747),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1763),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1787),
.B(n_1741),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1763),
.Y(n_1805)
);

NAND2x1_ASAP7_75t_L g1806 ( 
.A(n_1785),
.B(n_1754),
.Y(n_1806)
);

OR2x6_ASAP7_75t_L g1807 ( 
.A(n_1785),
.B(n_1734),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1764),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1761),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1776),
.A2(n_1730),
.B1(n_1736),
.B2(n_1737),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1761),
.Y(n_1811)
);

INVxp67_ASAP7_75t_SL g1812 ( 
.A(n_1774),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1764),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1768),
.B(n_1747),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1770),
.B(n_1782),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1765),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1770),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1741),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1765),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1786),
.A2(n_1733),
.B(n_1734),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1768),
.B(n_1747),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1766),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1766),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1771),
.B(n_1755),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1781),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1769),
.Y(n_1826)
);

INVxp33_ASAP7_75t_L g1827 ( 
.A(n_1788),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1782),
.B(n_1780),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1769),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1780),
.B(n_1721),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1787),
.B(n_1520),
.Y(n_1831)
);

NOR2xp67_ASAP7_75t_SL g1832 ( 
.A(n_1792),
.B(n_1737),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1772),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1766),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1786),
.B(n_1707),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1783),
.B(n_1750),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1772),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1773),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1783),
.B(n_1726),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1789),
.B(n_1726),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1795),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1807),
.B(n_1771),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1817),
.B(n_1779),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1799),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1795),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1796),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1807),
.B(n_1784),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1807),
.B(n_1784),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1807),
.B(n_1784),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1796),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1814),
.B(n_1784),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1814),
.B(n_1784),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1820),
.B(n_1779),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1803),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1801),
.A2(n_1726),
.B1(n_1693),
.B2(n_1742),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_SL g1856 ( 
.A(n_1832),
.B(n_1744),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1815),
.B(n_1789),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1821),
.B(n_1793),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1798),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1798),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1828),
.B(n_1778),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1830),
.B(n_1778),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1800),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1821),
.B(n_1793),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1803),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1806),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1810),
.B(n_1741),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1809),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1836),
.B(n_1791),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1797),
.B(n_1792),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1835),
.B(n_1791),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1812),
.A2(n_1806),
.B(n_1742),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1831),
.B(n_1520),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1805),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1827),
.B(n_1741),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1805),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1832),
.B(n_1520),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1858),
.B(n_1804),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1873),
.B(n_1683),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1858),
.B(n_1804),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1841),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1841),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1844),
.A2(n_1837),
.B1(n_1829),
.B2(n_1833),
.C(n_1826),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1863),
.B(n_1804),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1856),
.A2(n_1839),
.B(n_1840),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1856),
.A2(n_1818),
.B1(n_1797),
.B2(n_1802),
.Y(n_1886)
);

NOR3xp33_ASAP7_75t_L g1887 ( 
.A(n_1867),
.B(n_1833),
.C(n_1829),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1863),
.B(n_1837),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1851),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1853),
.B(n_1767),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1845),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1877),
.B(n_1818),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1845),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1846),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1853),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_SL g1896 ( 
.A1(n_1866),
.A2(n_1875),
.B(n_1855),
.Y(n_1896)
);

INVx5_ASAP7_75t_L g1897 ( 
.A(n_1866),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1869),
.B(n_1816),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1846),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1864),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1864),
.Y(n_1901)
);

NAND2xp33_ASAP7_75t_L g1902 ( 
.A(n_1847),
.B(n_1802),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1862),
.B(n_1767),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1850),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1881),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1895),
.B(n_1869),
.Y(n_1906)
);

O2A1O1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1896),
.A2(n_1872),
.B(n_1866),
.C(n_1849),
.Y(n_1907)
);

NAND2x1_ASAP7_75t_SL g1908 ( 
.A(n_1884),
.B(n_1847),
.Y(n_1908)
);

INVxp67_ASAP7_75t_SL g1909 ( 
.A(n_1900),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1879),
.B(n_1862),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1889),
.B(n_1870),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1901),
.B(n_1888),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1882),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1892),
.B(n_1870),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1878),
.B(n_1880),
.Y(n_1915)
);

OAI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1886),
.A2(n_1855),
.B1(n_1872),
.B2(n_1843),
.Y(n_1916)
);

AOI211xp5_ASAP7_75t_L g1917 ( 
.A1(n_1887),
.A2(n_1848),
.B(n_1849),
.C(n_1851),
.Y(n_1917)
);

O2A1O1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1885),
.A2(n_1848),
.B(n_1839),
.C(n_1842),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1900),
.A2(n_1842),
.B1(n_1852),
.B2(n_1843),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1891),
.Y(n_1920)
);

OAI21xp33_ASAP7_75t_L g1921 ( 
.A1(n_1902),
.A2(n_1852),
.B(n_1871),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1890),
.B(n_1871),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1897),
.Y(n_1923)
);

AND4x1_ASAP7_75t_L g1924 ( 
.A(n_1885),
.B(n_1672),
.C(n_1678),
.D(n_1647),
.Y(n_1924)
);

OAI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1897),
.A2(n_1861),
.B1(n_1818),
.B2(n_1743),
.Y(n_1925)
);

NAND4xp25_ASAP7_75t_SL g1926 ( 
.A(n_1907),
.B(n_1883),
.C(n_1888),
.D(n_1898),
.Y(n_1926)
);

OAI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1916),
.A2(n_1917),
.B1(n_1897),
.B2(n_1906),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1915),
.B(n_1884),
.Y(n_1928)
);

A2O1A1Ixp33_ASAP7_75t_L g1929 ( 
.A1(n_1908),
.A2(n_1918),
.B(n_1883),
.C(n_1921),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1909),
.A2(n_1898),
.B(n_1897),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1912),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1912),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1905),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1913),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1910),
.A2(n_1894),
.B(n_1893),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1911),
.A2(n_1903),
.B1(n_1861),
.B2(n_1857),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1914),
.A2(n_1906),
.B(n_1919),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1923),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1920),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_SL g1940 ( 
.A(n_1929),
.B(n_1927),
.C(n_1924),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1930),
.B(n_1922),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1938),
.Y(n_1942)
);

NAND5xp2_ASAP7_75t_L g1943 ( 
.A(n_1937),
.B(n_1899),
.C(n_1904),
.D(n_1854),
.E(n_1874),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1928),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1927),
.B(n_1925),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1933),
.Y(n_1946)
);

NAND4xp25_ASAP7_75t_L g1947 ( 
.A(n_1935),
.B(n_1932),
.C(n_1931),
.D(n_1936),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1934),
.Y(n_1948)
);

NAND4xp25_ASAP7_75t_SL g1949 ( 
.A(n_1926),
.B(n_1840),
.C(n_1857),
.D(n_1874),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1939),
.B(n_1850),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1949),
.A2(n_1876),
.B1(n_1865),
.B2(n_1854),
.C(n_1860),
.Y(n_1951)
);

NOR2x1_ASAP7_75t_L g1952 ( 
.A(n_1947),
.B(n_1940),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1943),
.A2(n_1876),
.B1(n_1865),
.B2(n_1868),
.C(n_1860),
.Y(n_1953)
);

OAI222xp33_ASAP7_75t_L g1954 ( 
.A1(n_1945),
.A2(n_1944),
.B1(n_1941),
.B2(n_1948),
.C1(n_1942),
.C2(n_1946),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1950),
.A2(n_1868),
.B(n_1860),
.C(n_1859),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1944),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1952),
.B(n_1868),
.C(n_1859),
.Y(n_1957)
);

OAI211xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1956),
.A2(n_1859),
.B(n_1825),
.C(n_1813),
.Y(n_1958)
);

XNOR2xp5_ASAP7_75t_L g1959 ( 
.A(n_1953),
.B(n_1658),
.Y(n_1959)
);

AOI221x1_ASAP7_75t_L g1960 ( 
.A1(n_1955),
.A2(n_1825),
.B1(n_1808),
.B2(n_1813),
.C(n_1819),
.Y(n_1960)
);

OAI211xp5_ASAP7_75t_SL g1961 ( 
.A1(n_1951),
.A2(n_1825),
.B(n_1819),
.C(n_1808),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1954),
.B(n_1781),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1954),
.A2(n_1809),
.B(n_1811),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1957),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1962),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1960),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1959),
.A2(n_1824),
.B1(n_1838),
.B2(n_1822),
.Y(n_1967)
);

INVx2_ASAP7_75t_SL g1968 ( 
.A(n_1958),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1961),
.Y(n_1969)
);

AOI322xp5_ASAP7_75t_L g1970 ( 
.A1(n_1964),
.A2(n_1963),
.A3(n_1824),
.B1(n_1777),
.B2(n_1834),
.C1(n_1822),
.C2(n_1811),
.Y(n_1970)
);

AOI21xp33_ASAP7_75t_L g1971 ( 
.A1(n_1965),
.A2(n_1834),
.B(n_1823),
.Y(n_1971)
);

NAND3x1_ASAP7_75t_L g1972 ( 
.A(n_1967),
.B(n_1838),
.C(n_1777),
.Y(n_1972)
);

NOR3xp33_ASAP7_75t_SL g1973 ( 
.A(n_1971),
.B(n_1968),
.C(n_1966),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1973),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1974),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1974),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1975),
.A2(n_1967),
.B1(n_1969),
.B2(n_1972),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_R g1978 ( 
.A1(n_1976),
.A2(n_1970),
.B1(n_1823),
.B2(n_1749),
.Y(n_1978)
);

AOI21xp33_ASAP7_75t_L g1979 ( 
.A1(n_1977),
.A2(n_1749),
.B(n_1628),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1978),
.A2(n_1790),
.B(n_1775),
.Y(n_1980)
);

OAI21xp33_ASAP7_75t_L g1981 ( 
.A1(n_1979),
.A2(n_1758),
.B(n_1749),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1981),
.A2(n_1980),
.B(n_1790),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1982),
.Y(n_1983)
);

OAI221xp5_ASAP7_75t_R g1984 ( 
.A1(n_1983),
.A2(n_1748),
.B1(n_1755),
.B2(n_1757),
.C(n_1686),
.Y(n_1984)
);

AOI211xp5_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1647),
.B(n_1506),
.C(n_1794),
.Y(n_1985)
);


endmodule