module fake_jpeg_12105_n_169 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVxp33_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_21),
.B(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_27),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_59),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_26),
.C(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_56),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_26),
.C(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_65),
.Y(n_89)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVxp67_ASAP7_75t_SL g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_15),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_46),
.B1(n_48),
.B2(n_34),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_24),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_25),
.B1(n_37),
.B2(n_16),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_37),
.B1(n_20),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_94),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_87),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_49),
.B1(n_54),
.B2(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_91),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_41),
.B1(n_20),
.B2(n_24),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_49),
.B1(n_72),
.B2(n_15),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_106),
.B1(n_82),
.B2(n_96),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_23),
.C(n_68),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_108),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_63),
.B1(n_70),
.B2(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_0),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_85),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_78),
.B(n_91),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_125),
.B(n_128),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_75),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_114),
.Y(n_132)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_39),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_93),
.B(n_63),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_134),
.C(n_141),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_99),
.C(n_102),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_103),
.B(n_98),
.C(n_110),
.D(n_112),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_125),
.B(n_122),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_103),
.B(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_145),
.B(n_148),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_115),
.B1(n_128),
.B2(n_120),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_4),
.B1(n_8),
.B2(n_10),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_131),
.C(n_132),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_139),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_122),
.C(n_10),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_135),
.B(n_123),
.Y(n_153)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_139),
.B1(n_141),
.B2(n_130),
.C(n_136),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_144),
.B(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_144),
.C(n_3),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_148),
.B(n_142),
.Y(n_156)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_11),
.B1(n_13),
.B2(n_2),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_155),
.B(n_151),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_SL g164 ( 
.A(n_162),
.B(n_160),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_154),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_162),
.C(n_156),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_163),
.B1(n_11),
.B2(n_3),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_163),
.Y(n_169)
);


endmodule