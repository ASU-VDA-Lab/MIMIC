module real_aes_82_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_0), .B(n_117), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_1), .A2(n_126), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_2), .B(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_3), .B(n_133), .Y(n_196) );
INVx1_ASAP7_75t_L g124 ( .A(n_4), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_5), .B(n_133), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_6), .B(n_137), .Y(n_466) );
INVx1_ASAP7_75t_L g500 ( .A(n_7), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g789 ( .A(n_8), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_9), .Y(n_538) );
NAND2xp33_ASAP7_75t_L g134 ( .A(n_10), .B(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g114 ( .A(n_11), .Y(n_114) );
AOI221x1_ASAP7_75t_L g212 ( .A1(n_12), .A2(n_24), .B1(n_117), .B2(n_126), .C(n_213), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_13), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_14), .B(n_117), .Y(n_116) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_15), .A2(n_112), .B(n_115), .Y(n_111) );
INVx1_ASAP7_75t_L g475 ( .A(n_16), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_17), .B(n_151), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_18), .B(n_133), .Y(n_160) );
AO21x1_ASAP7_75t_L g191 ( .A1(n_19), .A2(n_117), .B(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g434 ( .A(n_20), .Y(n_434) );
INVx1_ASAP7_75t_L g473 ( .A(n_21), .Y(n_473) );
INVx1_ASAP7_75t_SL g483 ( .A(n_22), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_23), .B(n_118), .Y(n_566) );
NAND2x1_ASAP7_75t_L g182 ( .A(n_25), .B(n_133), .Y(n_182) );
AOI33xp33_ASAP7_75t_L g512 ( .A1(n_26), .A2(n_50), .A3(n_450), .B1(n_455), .B2(n_513), .B3(n_514), .Y(n_512) );
NAND2x1_ASAP7_75t_L g170 ( .A(n_27), .B(n_135), .Y(n_170) );
INVx1_ASAP7_75t_L g532 ( .A(n_28), .Y(n_532) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_29), .A2(n_85), .B(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g138 ( .A(n_29), .B(n_85), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_30), .B(n_458), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_31), .B(n_135), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_32), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_33), .B(n_135), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_34), .A2(n_126), .B(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g123 ( .A(n_35), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g127 ( .A(n_35), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g449 ( .A(n_35), .Y(n_449) );
OR2x6_ASAP7_75t_L g432 ( .A(n_36), .B(n_433), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_37), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_38), .B(n_117), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_39), .B(n_458), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_40), .A2(n_137), .B1(n_144), .B2(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_41), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_42), .B(n_118), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_43), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_44), .B(n_135), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_45), .B(n_112), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_46), .B(n_118), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_47), .A2(n_126), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_48), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_49), .B(n_135), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_51), .B(n_118), .Y(n_524) );
INVx1_ASAP7_75t_L g120 ( .A(n_52), .Y(n_120) );
INVx1_ASAP7_75t_L g130 ( .A(n_52), .Y(n_130) );
AND2x2_ASAP7_75t_L g525 ( .A(n_53), .B(n_151), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_54), .A2(n_71), .B1(n_447), .B2(n_458), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_55), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_56), .B(n_133), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_57), .B(n_144), .Y(n_540) );
AOI21xp5_ASAP7_75t_SL g446 ( .A1(n_58), .A2(n_447), .B(n_452), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_59), .A2(n_126), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g469 ( .A(n_60), .Y(n_469) );
AO21x1_ASAP7_75t_L g193 ( .A1(n_61), .A2(n_126), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_62), .B(n_117), .Y(n_146) );
INVx1_ASAP7_75t_L g523 ( .A(n_63), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_64), .B(n_117), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_65), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_66), .A2(n_447), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g206 ( .A(n_67), .B(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g122 ( .A(n_68), .Y(n_122) );
INVx1_ASAP7_75t_L g128 ( .A(n_68), .Y(n_128) );
AND2x2_ASAP7_75t_L g174 ( .A(n_69), .B(n_143), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_70), .B(n_458), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_72), .A2(n_772), .B1(n_776), .B2(n_778), .Y(n_775) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_73), .A2(n_101), .B1(n_782), .B2(n_793), .C1(n_811), .C2(n_815), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g798 ( .A1(n_73), .A2(n_83), .B1(n_799), .B2(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_73), .Y(n_799) );
AND2x2_ASAP7_75t_L g485 ( .A(n_74), .B(n_143), .Y(n_485) );
INVx1_ASAP7_75t_L g470 ( .A(n_75), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_76), .A2(n_447), .B(n_482), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_77), .A2(n_447), .B(n_507), .C(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g435 ( .A(n_78), .Y(n_435) );
AND2x2_ASAP7_75t_L g142 ( .A(n_79), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_80), .B(n_117), .Y(n_162) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_81), .B(n_143), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_82), .A2(n_447), .B1(n_510), .B2(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g800 ( .A(n_83), .Y(n_800) );
AND2x2_ASAP7_75t_L g192 ( .A(n_84), .B(n_137), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_86), .B(n_135), .Y(n_161) );
AND2x2_ASAP7_75t_L g186 ( .A(n_87), .B(n_143), .Y(n_186) );
INVx1_ASAP7_75t_L g453 ( .A(n_88), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_89), .B(n_133), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_90), .A2(n_126), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_91), .B(n_135), .Y(n_214) );
AND2x2_ASAP7_75t_L g516 ( .A(n_92), .B(n_143), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_93), .A2(n_94), .B1(n_773), .B2(n_774), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_93), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_94), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_95), .B(n_133), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_96), .A2(n_530), .B(n_531), .C(n_533), .Y(n_529) );
BUFx2_ASAP7_75t_L g790 ( .A(n_97), .Y(n_790) );
BUFx2_ASAP7_75t_SL g819 ( .A(n_97), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_98), .A2(n_126), .B(n_131), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_99), .B(n_118), .Y(n_456) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_772), .B(n_775), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_427), .B1(n_436), .B2(n_770), .Y(n_104) );
INVx2_ASAP7_75t_L g777 ( .A(n_105), .Y(n_777) );
INVx1_ASAP7_75t_L g796 ( .A(n_105), .Y(n_796) );
INVx2_ASAP7_75t_L g802 ( .A(n_105), .Y(n_802) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_348), .Y(n_105) );
NOR3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_260), .C(n_300), .Y(n_106) );
OAI221xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_175), .B1(n_224), .B2(n_239), .C(n_242), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_139), .Y(n_109) );
INVx2_ASAP7_75t_L g257 ( .A(n_110), .Y(n_257) );
AND2x2_ASAP7_75t_L g287 ( .A(n_110), .B(n_288), .Y(n_287) );
BUFx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g225 ( .A(n_111), .B(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g232 ( .A(n_111), .B(n_165), .Y(n_232) );
INVx2_ASAP7_75t_L g238 ( .A(n_111), .Y(n_238) );
AND2x2_ASAP7_75t_L g247 ( .A(n_111), .B(n_141), .Y(n_247) );
INVx1_ASAP7_75t_L g263 ( .A(n_111), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_111), .B(n_309), .Y(n_308) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_112), .A2(n_498), .B(n_502), .Y(n_497) );
INVx2_ASAP7_75t_SL g507 ( .A(n_112), .Y(n_507) );
BUFx4f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx3_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
AND2x4_ASAP7_75t_L g137 ( .A(n_114), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_114), .B(n_138), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_125), .B(n_137), .Y(n_115) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_123), .Y(n_117) );
INVx1_ASAP7_75t_L g471 ( .A(n_118), .Y(n_471) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
AND2x6_ASAP7_75t_L g135 ( .A(n_119), .B(n_128), .Y(n_135) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g133 ( .A(n_121), .B(n_130), .Y(n_133) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx5_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_123), .Y(n_533) );
AND2x2_ASAP7_75t_L g129 ( .A(n_124), .B(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_124), .Y(n_460) );
AND2x6_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
BUFx3_ASAP7_75t_L g461 ( .A(n_127), .Y(n_461) );
INVx2_ASAP7_75t_L g451 ( .A(n_128), .Y(n_451) );
AND2x4_ASAP7_75t_L g447 ( .A(n_129), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g455 ( .A(n_130), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_134), .B(n_136), .Y(n_131) );
INVxp67_ASAP7_75t_L g476 ( .A(n_133), .Y(n_476) );
INVxp67_ASAP7_75t_L g474 ( .A(n_135), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_136), .A2(n_149), .B(n_150), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_136), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_136), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_136), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_136), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_136), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_136), .A2(n_214), .B(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_136), .A2(n_453), .B(n_454), .C(n_456), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_136), .B(n_137), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_136), .A2(n_454), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_SL g499 ( .A1(n_136), .A2(n_454), .B(n_500), .C(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g510 ( .A(n_136), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_136), .A2(n_454), .B(n_523), .C(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_136), .A2(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_SL g156 ( .A(n_137), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_137), .B(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_137), .A2(n_446), .B(n_457), .Y(n_445) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_153), .Y(n_139) );
INVx4_ASAP7_75t_L g228 ( .A(n_140), .Y(n_228) );
AND2x2_ASAP7_75t_L g259 ( .A(n_140), .B(n_166), .Y(n_259) );
AND2x2_ASAP7_75t_L g335 ( .A(n_140), .B(n_309), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_140), .B(n_165), .Y(n_377) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_141), .B(n_165), .Y(n_264) );
AND2x2_ASAP7_75t_L g288 ( .A(n_141), .B(n_166), .Y(n_288) );
BUFx2_ASAP7_75t_L g304 ( .A(n_141), .Y(n_304) );
NOR2x1_ASAP7_75t_SL g407 ( .A(n_141), .B(n_309), .Y(n_407) );
OR2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_145), .Y(n_141) );
INVx3_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_143), .A2(n_185), .B1(n_529), .B2(n_534), .Y(n_528) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_144), .B(n_537), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_151), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_151), .Y(n_173) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_151), .A2(n_212), .B(n_216), .Y(n_211) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_151), .A2(n_212), .B(n_216), .Y(n_274) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g284 ( .A(n_153), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_153), .A2(n_351), .B1(n_353), .B2(n_355), .C(n_360), .Y(n_350) );
AND2x2_ASAP7_75t_L g370 ( .A(n_153), .B(n_263), .Y(n_370) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_165), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g226 ( .A(n_155), .Y(n_226) );
INVx1_ASAP7_75t_L g279 ( .A(n_155), .Y(n_279) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_163), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_156), .B(n_164), .Y(n_163) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_156), .A2(n_157), .B(n_163), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_162), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_165), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g248 ( .A(n_165), .B(n_236), .Y(n_248) );
INVx2_ASAP7_75t_L g290 ( .A(n_165), .Y(n_290) );
AND2x2_ASAP7_75t_L g423 ( .A(n_165), .B(n_238), .Y(n_423) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_166), .Y(n_280) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_173), .B(n_174), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_173), .A2(n_479), .B(n_485), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_207), .C(n_222), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_187), .Y(n_176) );
INVx2_ASAP7_75t_L g337 ( .A(n_177), .Y(n_337) );
AND2x2_ASAP7_75t_L g382 ( .A(n_177), .B(n_259), .Y(n_382) );
BUFx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g327 ( .A(n_178), .Y(n_327) );
AND2x4_ASAP7_75t_SL g342 ( .A(n_178), .B(n_254), .Y(n_342) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_185), .B(n_186), .Y(n_178) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_179), .A2(n_185), .B(n_186), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_184), .Y(n_179) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_185), .A2(n_200), .B(n_206), .Y(n_199) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_185), .A2(n_200), .B(n_206), .Y(n_219) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_185), .A2(n_519), .B(n_525), .Y(n_518) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_185), .A2(n_519), .B(n_525), .Y(n_548) );
INVx2_ASAP7_75t_L g296 ( .A(n_187), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_187), .B(n_326), .Y(n_352) );
AND2x4_ASAP7_75t_L g385 ( .A(n_187), .B(n_332), .Y(n_385) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
AND2x2_ASAP7_75t_L g223 ( .A(n_188), .B(n_218), .Y(n_223) );
OR2x2_ASAP7_75t_L g253 ( .A(n_188), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_188), .B(n_274), .Y(n_322) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g267 ( .A(n_189), .Y(n_267) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g241 ( .A(n_190), .Y(n_241) );
OAI21x1_ASAP7_75t_SL g190 ( .A1(n_191), .A2(n_193), .B(n_197), .Y(n_190) );
INVx1_ASAP7_75t_L g198 ( .A(n_192), .Y(n_198) );
INVx2_ASAP7_75t_L g254 ( .A(n_199), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_201), .B(n_205), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_207), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_217), .Y(n_208) );
AND2x2_ASAP7_75t_L g222 ( .A(n_209), .B(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g295 ( .A(n_209), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g380 ( .A(n_209), .Y(n_380) );
BUFx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x4_ASAP7_75t_L g240 ( .A(n_210), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g359 ( .A(n_210), .B(n_219), .Y(n_359) );
AND2x2_ASAP7_75t_L g363 ( .A(n_210), .B(n_229), .Y(n_363) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g332 ( .A(n_211), .Y(n_332) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_211), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_217), .B(n_240), .Y(n_316) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_218), .B(n_241), .Y(n_426) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g230 ( .A(n_219), .B(n_221), .Y(n_230) );
AND2x2_ASAP7_75t_L g312 ( .A(n_219), .B(n_274), .Y(n_312) );
AND2x2_ASAP7_75t_L g331 ( .A(n_219), .B(n_220), .Y(n_331) );
BUFx2_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_220), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
BUFx3_ASAP7_75t_L g229 ( .A(n_221), .Y(n_229) );
INVxp67_ASAP7_75t_L g272 ( .A(n_221), .Y(n_272) );
INVx1_ASAP7_75t_L g245 ( .A(n_223), .Y(n_245) );
AND2x2_ASAP7_75t_L g281 ( .A(n_223), .B(n_252), .Y(n_281) );
NAND2xp33_ASAP7_75t_L g362 ( .A(n_223), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g399 ( .A(n_223), .B(n_400), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_227), .B1(n_230), .B2(n_231), .C(n_233), .Y(n_224) );
AND2x2_ASAP7_75t_L g328 ( .A(n_225), .B(n_228), .Y(n_328) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_225), .B(n_288), .Y(n_347) );
AND2x2_ASAP7_75t_L g365 ( .A(n_225), .B(n_290), .Y(n_365) );
AND2x2_ASAP7_75t_L g420 ( .A(n_225), .B(n_259), .Y(n_420) );
INVx1_ASAP7_75t_L g236 ( .A(n_226), .Y(n_236) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_226), .Y(n_292) );
CKINVDCx16_ASAP7_75t_R g372 ( .A(n_227), .Y(n_372) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_228), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_228), .B(n_279), .Y(n_354) );
AND2x2_ASAP7_75t_L g321 ( .A(n_229), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g357 ( .A(n_229), .Y(n_357) );
AND2x2_ASAP7_75t_L g266 ( .A(n_230), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_230), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g408 ( .A(n_230), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_230), .B(n_332), .Y(n_418) );
AND2x4_ASAP7_75t_L g334 ( .A(n_231), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g405 ( .A(n_232), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
OR2x2_ASAP7_75t_L g276 ( .A(n_237), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g283 ( .A(n_238), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g314 ( .A(n_238), .B(n_288), .Y(n_314) );
AND2x2_ASAP7_75t_L g388 ( .A(n_238), .B(n_309), .Y(n_388) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g336 ( .A(n_240), .B(n_337), .Y(n_336) );
OAI32xp33_ASAP7_75t_L g401 ( .A1(n_240), .A2(n_402), .A3(n_404), .B1(n_405), .B2(n_408), .Y(n_401) );
AND2x4_ASAP7_75t_L g273 ( .A(n_241), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g371 ( .A(n_241), .B(n_274), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_246), .B1(n_249), .B2(n_255), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g360 ( .A1(n_244), .A2(n_258), .B(n_361), .C(n_362), .Y(n_360) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g344 ( .A(n_245), .B(n_272), .Y(n_344) );
INVx1_ASAP7_75t_SL g415 ( .A(n_246), .Y(n_415) );
AND2x4_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x4_ASAP7_75t_L g318 ( .A(n_248), .B(n_257), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_248), .A2(n_397), .B1(n_398), .B2(n_399), .C(n_401), .Y(n_396) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_253), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_256), .A2(n_286), .B1(n_339), .B2(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_257), .A2(n_375), .B(n_383), .C(n_396), .Y(n_374) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g294 ( .A(n_259), .B(n_263), .Y(n_294) );
OAI211xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_265), .B(n_268), .C(n_297), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g291 ( .A(n_263), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g411 ( .A(n_263), .B(n_407), .Y(n_411) );
OAI32xp33_ASAP7_75t_L g368 ( .A1(n_264), .A2(n_369), .A3(n_371), .B1(n_372), .B2(n_373), .Y(n_368) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_SL g358 ( .A(n_267), .B(n_359), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_275), .B1(n_281), .B2(n_282), .C(n_285), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g425 ( .A(n_272), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_273), .B(n_337), .Y(n_339) );
A2O1A1O1Ixp25_ASAP7_75t_L g410 ( .A1(n_273), .A2(n_342), .B(n_358), .C(n_404), .D(n_411), .Y(n_410) );
AOI31xp33_ASAP7_75t_L g412 ( .A1(n_273), .A2(n_294), .A3(n_404), .B(n_411), .Y(n_412) );
AND2x2_ASAP7_75t_L g326 ( .A(n_274), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_276), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx2_ASAP7_75t_L g403 ( .A(n_278), .Y(n_403) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g398 ( .A(n_279), .B(n_290), .Y(n_398) );
INVx1_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
AND2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AOI31xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .A3(n_293), .B(n_295), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_288), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g421 ( .A(n_288), .B(n_367), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g366 ( .A(n_290), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g392 ( .A(n_290), .Y(n_392) );
INVxp67_ASAP7_75t_L g361 ( .A(n_291), .Y(n_361) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g299 ( .A(n_295), .Y(n_299) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND3xp33_ASAP7_75t_SL g300 ( .A(n_301), .B(n_317), .C(n_333), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_310), .B1(n_314), .B2(n_315), .Y(n_301) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx2_ASAP7_75t_L g387 ( .A(n_304), .Y(n_387) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_308), .Y(n_367) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_308), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_308), .B(n_377), .Y(n_394) );
NAND2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_328), .B2(n_329), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_326), .A2(n_331), .B1(n_365), .B2(n_366), .C(n_368), .Y(n_364) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g404 ( .A(n_331), .Y(n_404) );
AND2x2_ASAP7_75t_L g341 ( .A(n_332), .B(n_342), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_SL g389 ( .A1(n_332), .A2(n_390), .B(n_394), .C(n_395), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_338), .C(n_343), .Y(n_333) );
AND2x2_ASAP7_75t_L g384 ( .A(n_337), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
AOI21xp33_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_345), .B(n_346), .Y(n_343) );
INVx2_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NOR3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_374), .C(n_409), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_350), .B(n_364), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g373 ( .A(n_358), .Y(n_373) );
INVxp67_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g381 ( .A(n_371), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B1(n_381), .B2(n_382), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B(n_389), .Y(n_383) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g422 ( .A(n_407), .B(n_423), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_413), .B2(n_416), .C(n_419), .Y(n_409) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI31xp33_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .A3(n_422), .B(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx4_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx3_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_429), .A2(n_437), .B1(n_770), .B2(n_777), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
AND2x6_ASAP7_75t_SL g430 ( .A(n_431), .B(n_432), .Y(n_430) );
OR2x6_ASAP7_75t_SL g770 ( .A(n_431), .B(n_771), .Y(n_770) );
OR2x2_ASAP7_75t_L g781 ( .A(n_431), .B(n_432), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_431), .B(n_771), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_432), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_657), .C(n_734), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_609), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_440), .B(n_549), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_486), .B1(n_493), .B2(n_542), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_462), .Y(n_441) );
NOR2xp67_ASAP7_75t_SL g592 ( .A(n_442), .B(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g607 ( .A(n_442), .B(n_608), .Y(n_607) );
NOR2x1_ASAP7_75t_L g624 ( .A(n_442), .B(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_SL g664 ( .A(n_442), .B(n_665), .Y(n_664) );
INVx4_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_443), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_443), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g599 ( .A(n_443), .Y(n_599) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_443), .Y(n_604) );
AND2x2_ASAP7_75t_L g633 ( .A(n_443), .B(n_573), .Y(n_633) );
OR2x2_ASAP7_75t_L g637 ( .A(n_443), .B(n_478), .Y(n_637) );
AND2x4_ASAP7_75t_L g650 ( .A(n_443), .B(n_608), .Y(n_650) );
NOR2x1_ASAP7_75t_SL g652 ( .A(n_443), .B(n_465), .Y(n_652) );
AND2x2_ASAP7_75t_L g680 ( .A(n_443), .B(n_558), .Y(n_680) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVxp67_ASAP7_75t_L g539 ( .A(n_447), .Y(n_539) );
NOR2x1p5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x6_ASAP7_75t_L g454 ( .A(n_451), .B(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_454), .A2(n_469), .B1(n_470), .B2(n_471), .Y(n_468) );
INVxp67_ASAP7_75t_L g530 ( .A(n_454), .Y(n_530) );
INVx2_ASAP7_75t_L g568 ( .A(n_454), .Y(n_568) );
AND2x2_ASAP7_75t_L g459 ( .A(n_455), .B(n_460), .Y(n_459) );
INVxp33_ASAP7_75t_L g513 ( .A(n_455), .Y(n_513) );
INVx1_ASAP7_75t_L g541 ( .A(n_458), .Y(n_541) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g561 ( .A(n_459), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_461), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_462), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_463), .A2(n_738), .B1(n_740), .B2(n_743), .Y(n_737) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_478), .Y(n_463) );
INVx1_ASAP7_75t_L g492 ( .A(n_464), .Y(n_492) );
AND2x2_ASAP7_75t_L g595 ( .A(n_464), .B(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g600 ( .A(n_464), .B(n_558), .Y(n_600) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g557 ( .A(n_465), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g573 ( .A(n_465), .Y(n_573) );
AND2x2_ASAP7_75t_L g606 ( .A(n_465), .B(n_478), .Y(n_606) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_472), .B(n_477), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_471), .B(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_472) );
INVx2_ASAP7_75t_L g490 ( .A(n_478), .Y(n_490) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_478), .Y(n_575) );
INVx1_ASAP7_75t_L g594 ( .A(n_478), .Y(n_594) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_478), .Y(n_663) );
INVx1_ASAP7_75t_L g675 ( .A(n_478), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI31xp33_ASAP7_75t_SL g729 ( .A1(n_487), .A2(n_730), .A3(n_731), .B(n_732), .Y(n_729) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_488), .B(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g654 ( .A(n_489), .B(n_556), .Y(n_654) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g570 ( .A(n_490), .Y(n_570) );
AND2x4_ASAP7_75t_SL g690 ( .A(n_492), .B(n_594), .Y(n_690) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_493), .A2(n_611), .B(n_614), .Y(n_610) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
INVx2_ASAP7_75t_L g583 ( .A(n_494), .Y(n_583) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g710 ( .A(n_495), .B(n_618), .Y(n_710) );
BUFx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g620 ( .A(n_496), .B(n_526), .Y(n_620) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVxp67_ASAP7_75t_L g545 ( .A(n_497), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_497), .B(n_506), .Y(n_580) );
AND2x4_ASAP7_75t_L g590 ( .A(n_497), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g635 ( .A(n_497), .B(n_527), .Y(n_635) );
INVx2_ASAP7_75t_L g643 ( .A(n_497), .Y(n_643) );
INVx1_ASAP7_75t_L g742 ( .A(n_497), .Y(n_742) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_497), .Y(n_751) );
INVx1_ASAP7_75t_L g688 ( .A(n_503), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_504), .B(n_517), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g544 ( .A(n_505), .B(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g683 ( .A(n_505), .B(n_618), .Y(n_683) );
AND2x2_ASAP7_75t_L g700 ( .A(n_505), .B(n_518), .Y(n_700) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_506), .B(n_548), .Y(n_723) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_516), .Y(n_506) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_507), .A2(n_508), .B(n_516), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g646 ( .A(n_517), .B(n_544), .Y(n_646) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_526), .Y(n_517) );
INVx2_ASAP7_75t_L g552 ( .A(n_518), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g733 ( .A(n_518), .B(n_526), .Y(n_733) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_518), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AND2x2_ASAP7_75t_L g649 ( .A(n_526), .B(n_553), .Y(n_649) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_527), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g578 ( .A(n_527), .Y(n_578) );
AND2x4_ASAP7_75t_L g642 ( .A(n_527), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g672 ( .A(n_527), .Y(n_672) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_535), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_539), .B1(n_540), .B2(n_541), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_543), .A2(n_556), .B1(n_694), .B2(n_695), .C(n_696), .Y(n_693) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g670 ( .A(n_544), .B(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g713 ( .A(n_544), .Y(n_713) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g656 ( .A(n_547), .B(n_580), .Y(n_656) );
INVx3_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
AND2x2_ASAP7_75t_L g750 ( .A(n_548), .B(n_751), .Y(n_750) );
NAND3xp33_ASAP7_75t_SL g549 ( .A(n_550), .B(n_581), .C(n_597), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_554), .B1(n_571), .B2(n_576), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_551), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g681 ( .A(n_551), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g692 ( .A(n_551), .B(n_587), .Y(n_692) );
AND2x2_ASAP7_75t_L g762 ( .A(n_551), .B(n_635), .Y(n_762) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g591 ( .A(n_553), .Y(n_591) );
INVx1_ASAP7_75t_L g640 ( .A(n_553), .Y(n_640) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI222xp33_ASAP7_75t_L g707 ( .A1(n_555), .A2(n_708), .B1(n_709), .B2(n_711), .C1(n_712), .C2(n_714), .Y(n_707) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_569), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_556), .B(n_583), .Y(n_582) );
NOR2x1_ASAP7_75t_L g715 ( .A(n_556), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g674 ( .A(n_557), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g730 ( .A(n_557), .B(n_604), .Y(n_730) );
INVx2_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
INVx1_ASAP7_75t_L g608 ( .A(n_558), .Y(n_608) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_558), .Y(n_665) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_564), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_563), .Y(n_560) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_570), .Y(n_613) );
INVx3_ASAP7_75t_L g632 ( .A(n_570), .Y(n_632) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g698 ( .A(n_572), .Y(n_698) );
NAND2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g685 ( .A(n_574), .Y(n_685) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g686 ( .A(n_577), .Y(n_686) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g587 ( .A(n_578), .Y(n_587) );
AND2x2_ASAP7_75t_L g705 ( .A(n_578), .B(n_590), .Y(n_705) );
AND2x2_ASAP7_75t_L g768 ( .A(n_578), .B(n_700), .Y(n_768) );
AND2x2_ASAP7_75t_L g697 ( .A(n_579), .B(n_617), .Y(n_697) );
INVx1_ASAP7_75t_L g708 ( .A(n_579), .Y(n_708) );
AND2x2_ASAP7_75t_L g725 ( .A(n_579), .B(n_672), .Y(n_725) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B1(n_588), .B2(n_592), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g597 ( .A1(n_584), .A2(n_598), .B(n_601), .Y(n_597) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g629 ( .A(n_587), .B(n_590), .Y(n_629) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g732 ( .A(n_590), .B(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g695 ( .A(n_593), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
AND2x2_ASAP7_75t_SL g603 ( .A(n_595), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g668 ( .A(n_595), .Y(n_668) );
AND2x2_ASAP7_75t_L g766 ( .A(n_595), .B(n_663), .Y(n_766) );
INVx1_ASAP7_75t_L g721 ( .A(n_596), .Y(n_721) );
INVx1_ASAP7_75t_L g627 ( .A(n_598), .Y(n_627) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g716 ( .A(n_599), .Y(n_716) );
INVx4_ASAP7_75t_L g625 ( .A(n_600), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI32xp33_ASAP7_75t_L g696 ( .A1(n_603), .A2(n_697), .A3(n_698), .B1(n_699), .B2(n_700), .Y(n_696) );
AND2x2_ASAP7_75t_L g691 ( .A(n_604), .B(n_606), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_SL g754 ( .A1(n_604), .A2(n_755), .B(n_756), .C(n_758), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_SL g719 ( .A(n_606), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g758 ( .A(n_606), .Y(n_758) );
AND2x2_ASAP7_75t_L g612 ( .A(n_607), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g739 ( .A(n_607), .Y(n_739) );
AND2x2_ASAP7_75t_L g745 ( .A(n_607), .B(n_632), .Y(n_745) );
NOR3x1_ASAP7_75t_L g609 ( .A(n_610), .B(n_626), .C(n_644), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_621), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AND2x2_ASAP7_75t_L g634 ( .A(n_617), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g677 ( .A(n_617), .B(n_642), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_617), .B(n_663), .Y(n_704) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_625), .B(n_632), .Y(n_731) );
INVx2_ASAP7_75t_L g753 ( .A(n_625), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B(n_630), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_627), .A2(n_718), .B1(n_722), .B2(n_724), .C(n_729), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_628), .A2(n_748), .B1(n_749), .B2(n_752), .Y(n_747) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B1(n_636), .B2(n_638), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x2_ASAP7_75t_L g676 ( .A(n_632), .B(n_652), .Y(n_676) );
INVx1_ASAP7_75t_L g682 ( .A(n_632), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_632), .B(n_650), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_635), .B(n_703), .Y(n_769) );
NAND2x1_ASAP7_75t_L g752 ( .A(n_636), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
NOR2x1_ASAP7_75t_L g667 ( .A(n_637), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2x1_ASAP7_75t_SL g755 ( .A(n_640), .B(n_642), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_640), .B(n_740), .Y(n_761) );
OR2x2_ASAP7_75t_L g722 ( .A(n_641), .B(n_723), .Y(n_722) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g757 ( .A(n_642), .B(n_683), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_645), .B(n_651), .Y(n_644) );
OAI21xp33_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_647), .B(n_650), .Y(n_645) );
OR2x2_ASAP7_75t_L g709 ( .A(n_648), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g743 ( .A(n_649), .B(n_741), .Y(n_743) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_650), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g699 ( .A(n_650), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_655), .Y(n_651) );
AND2x2_ASAP7_75t_L g684 ( .A(n_652), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_701), .Y(n_658) );
NOR3xp33_ASAP7_75t_SL g659 ( .A(n_660), .B(n_678), .C(n_693), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_666), .B(n_669), .C(n_673), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g727 ( .A(n_672), .Y(n_727) );
AND2x2_ASAP7_75t_L g740 ( .A(n_672), .B(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g748 ( .A(n_674), .Y(n_748) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_686), .B(n_687), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B1(n_683), .B2(n_684), .Y(n_679) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_680), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_691), .B2(n_692), .Y(n_687) );
INVx1_ASAP7_75t_SL g694 ( .A(n_692), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_698), .B(n_739), .Y(n_738) );
OAI22xp33_ASAP7_75t_SL g764 ( .A1(n_699), .A2(n_765), .B1(n_767), .B2(n_769), .Y(n_764) );
AOI211x1_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_706), .B(n_707), .C(n_717), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_719), .A2(n_760), .B(n_762), .Y(n_759) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g728 ( .A(n_723), .Y(n_728) );
NOR2xp67_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_726), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND4xp25_ASAP7_75t_L g735 ( .A(n_736), .B(n_746), .C(n_759), .D(n_763), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_744), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_754), .Y(n_746) );
INVxp67_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_791), .Y(n_784) );
INVxp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g786 ( .A(n_787), .B(n_790), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OR2x2_ASAP7_75t_SL g814 ( .A(n_788), .B(n_790), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_788), .A2(n_817), .B(n_820), .Y(n_816) );
INVx1_ASAP7_75t_SL g804 ( .A(n_791), .Y(n_804) );
BUFx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx3_ASAP7_75t_L g809 ( .A(n_792), .Y(n_809) );
BUFx2_ASAP7_75t_L g821 ( .A(n_792), .Y(n_821) );
INVxp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_803), .B(n_805), .Y(n_794) );
OAI22xp5_ASAP7_75t_SL g795 ( .A1(n_796), .A2(n_797), .B1(n_798), .B2(n_801), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_SL g805 ( .A(n_806), .B(n_810), .Y(n_805) );
INVx1_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
CKINVDCx11_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
CKINVDCx8_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
endmodule