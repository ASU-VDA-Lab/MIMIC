module fake_jpeg_2667_n_228 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_228);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_11),
.B(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_63),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_99),
.Y(n_109)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_55),
.B1(n_56),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_74),
.B1(n_76),
.B2(n_58),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_56),
.B1(n_68),
.B2(n_79),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_74),
.C(n_58),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_90),
.B1(n_96),
.B2(n_89),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_106),
.B1(n_118),
.B2(n_70),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_64),
.B(n_76),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_107),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_67),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_96),
.B1(n_89),
.B2(n_93),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_54),
.B1(n_88),
.B2(n_73),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_62),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_116),
.Y(n_128)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_60),
.B1(n_77),
.B2(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_139),
.B1(n_131),
.B2(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_79),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_115),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_64),
.B1(n_72),
.B2(n_61),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_130),
.B(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_134),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_61),
.B1(n_72),
.B2(n_71),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_60),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_1),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_65),
.B(n_57),
.C(n_70),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_43),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_65),
.B1(n_57),
.B2(n_2),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_104),
.B1(n_57),
.B2(n_2),
.Y(n_148)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_152),
.Y(n_180)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_150),
.B1(n_157),
.B2(n_164),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_158),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_159),
.B1(n_13),
.B2(n_14),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_4),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_165),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_50),
.B1(n_45),
.B2(n_44),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_8),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_128),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_9),
.B(n_10),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_10),
.B(n_12),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_9),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_173),
.Y(n_187)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_168),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_129),
.B1(n_136),
.B2(n_121),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_148),
.B(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_186),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_176),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_183),
.B(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_35),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_185),
.B(n_34),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_26),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_146),
.B(n_155),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_188),
.A2(n_197),
.B(n_172),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_142),
.C(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_178),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_196),
.B1(n_173),
.B2(n_176),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_175),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_33),
.B(n_32),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_199),
.B(n_200),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_166),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_204),
.B1(n_195),
.B2(n_194),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_174),
.B1(n_180),
.B2(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_170),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_207),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_206),
.A2(n_208),
.B1(n_193),
.B2(n_180),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_212),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_211),
.C(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_R g217 ( 
.A(n_213),
.B(n_204),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_177),
.C(n_30),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_210),
.C(n_214),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_186),
.B(n_29),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_28),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_19),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_219),
.B(n_168),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_20),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_24),
.C2(n_25),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_24),
.B(n_25),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_227),
.Y(n_228)
);


endmodule