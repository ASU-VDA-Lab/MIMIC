module real_jpeg_20534_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_267, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_267;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_202;
wire n_213;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_0),
.A2(n_3),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_0),
.A2(n_26),
.B1(n_29),
.B2(n_38),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_0),
.A2(n_5),
.B1(n_38),
.B2(n_62),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_1),
.A2(n_19),
.B1(n_26),
.B2(n_29),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_1),
.A2(n_5),
.B1(n_19),
.B2(n_62),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_3),
.B1(n_37),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_49),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_26),
.B1(n_29),
.B2(n_49),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_5),
.B1(n_49),
.B2(n_62),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_7),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_3),
.A2(n_35),
.B(n_42),
.C(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_4),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_5),
.A2(n_10),
.B1(n_60),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_5),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_7),
.B1(n_42),
.B2(n_62),
.Y(n_146)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_5),
.A2(n_7),
.B(n_10),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_7),
.A2(n_20),
.B1(n_21),
.B2(n_42),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_7),
.A2(n_26),
.B1(n_29),
.B2(n_42),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_7),
.A2(n_20),
.B(n_45),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_7),
.B(n_52),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_7),
.A2(n_27),
.B(n_29),
.Y(n_207)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_35),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_34),
.B(n_37),
.C(n_44),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_26),
.B1(n_29),
.B2(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_10),
.Y(n_60)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_82),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_81),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_64),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_16),
.B(n_64),
.Y(n_81)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_16),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_33),
.CI(n_46),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_18),
.A2(n_24),
.B1(n_30),
.B2(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_20),
.A2(n_28),
.B(n_42),
.C(n_207),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_25),
.B(n_27),
.C(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_27),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_23),
.B(n_80),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_24),
.A2(n_79),
.B(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_25),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_25),
.A2(n_31),
.B1(n_80),
.B2(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_25),
.B(n_42),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_29),
.A2(n_42),
.B(n_60),
.C(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_34),
.B(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_48),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_42),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_42),
.B(n_61),
.Y(n_190)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.C(n_55),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_47),
.B(n_111),
.C(n_118),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_47),
.A2(n_67),
.B1(n_104),
.B2(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_47),
.B(n_152),
.C(n_153),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_47),
.A2(n_67),
.B1(n_118),
.B2(n_163),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_55),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_57),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_61),
.B1(n_63),
.B2(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_61),
.B1(n_102),
.B2(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_62),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_72),
.C(n_74),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.C(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_73),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_72),
.A2(n_73),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_72),
.A2(n_73),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_118),
.C(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_73),
.B(n_238),
.C(n_240),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_127),
.A3(n_131),
.B1(n_263),
.B2(n_264),
.C(n_267),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_119),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_84),
.B(n_119),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_103),
.C(n_109),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_85),
.B(n_103),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_97),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_94),
.B2(n_96),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_87),
.A2(n_88),
.B1(n_98),
.B2(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_94),
.B(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_90),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_93),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_91),
.A2(n_92),
.B1(n_146),
.B2(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_98),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_102),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B(n_108),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_107),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_168),
.C(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_104),
.A2(n_152),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_121),
.C(n_124),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_109),
.A2(n_110),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_111),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_112),
.A2(n_116),
.B1(n_199),
.B2(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_112),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_114),
.B(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_145),
.B(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_116),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_157),
.C(n_198),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_116),
.A2(n_199),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_116),
.B(n_217),
.C(n_222),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_148),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_118),
.A2(n_138),
.B1(n_139),
.B2(n_163),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_118),
.B(n_139),
.C(n_205),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_128),
.B(n_129),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_257),
.B(n_262),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_245),
.B(n_256),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_173),
.B(n_230),
.C(n_244),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_159),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_135),
.B(n_159),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_150),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_137),
.B(n_147),
.C(n_150),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_139),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_138),
.B(n_143),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_139),
.B(n_182),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

NOR2x1_ASAP7_75t_R g189 ( 
.A(n_157),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_190),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_157),
.A2(n_166),
.B1(n_196),
.B2(n_200),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.C(n_167),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_167),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_229),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_224),
.B(n_228),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_214),
.B(n_223),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_202),
.B(n_213),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_193),
.B(n_201),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_192),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_191),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_204),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_211),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_221),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_242),
.B2(n_243),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_237),
.C(n_243),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_247),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_253),
.C(n_255),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_259),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);


endmodule