module fake_jpeg_28416_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_10),
.B1(n_12),
.B2(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_10),
.B1(n_12),
.B2(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_25),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_41),
.B(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_43),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_23),
.B(n_26),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_45),
.B1(n_27),
.B2(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_21),
.B1(n_36),
.B2(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_37),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_34),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_35),
.C(n_25),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_56),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_43),
.B(n_41),
.C(n_37),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_57),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_72),
.C(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_76),
.Y(n_83)
);

AOI21x1_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_51),
.B(n_28),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_73),
.B(n_75),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_35),
.C(n_25),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_27),
.B(n_2),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_27),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_74),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

A2O1A1O1Ixp25_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_63),
.B(n_65),
.C(n_59),
.D(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_67),
.B(n_27),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_82),
.B1(n_75),
.B2(n_29),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_68),
.C(n_72),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_20),
.B(n_19),
.C(n_16),
.D(n_13),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_29),
.B1(n_33),
.B2(n_19),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_90),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_33),
.C(n_29),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_33),
.B1(n_16),
.B2(n_4),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_83),
.B(n_89),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_95),
.B(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_3),
.B(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

AOI31xp33_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_3),
.A3(n_6),
.B(n_7),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_6),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_6),
.B(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_9),
.Y(n_101)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_102),
.B(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_8),
.Y(n_104)
);


endmodule