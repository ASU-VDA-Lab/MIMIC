module fake_jpeg_9266_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_41),
.CON(n_74),
.SN(n_74)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_46),
.Y(n_64)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_62),
.B(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_30),
.B(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_76),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_17),
.B(n_33),
.Y(n_69)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_72),
.C(n_31),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_30),
.B1(n_32),
.B2(n_31),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_75),
.B1(n_24),
.B2(n_23),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_22),
.B(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_22),
.B1(n_27),
.B2(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_79),
.B(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_87),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g132 ( 
.A(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_95),
.Y(n_129)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_63),
.Y(n_89)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_90),
.A2(n_96),
.B1(n_100),
.B2(n_16),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_40),
.C(n_39),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_53),
.Y(n_117)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_98),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_64),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_58),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_61),
.Y(n_133)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_76),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_122),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_90),
.B(n_93),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_97),
.B(n_26),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_34),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_128),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_85),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_82),
.B(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_34),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_99),
.B1(n_61),
.B2(n_113),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_96),
.B1(n_78),
.B2(n_84),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_115),
.B1(n_77),
.B2(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_34),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_142),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_25),
.B1(n_19),
.B2(n_37),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_34),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_82),
.A2(n_29),
.B(n_26),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_28),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_147),
.A2(n_151),
.B(n_155),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_148),
.A2(n_176),
.B1(n_116),
.B2(n_132),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_158),
.B1(n_126),
.B2(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_150),
.B(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_86),
.B1(n_77),
.B2(n_103),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_140),
.B1(n_135),
.B2(n_119),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_111),
.C(n_45),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_162),
.C(n_164),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_16),
.B(n_35),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_45),
.B1(n_95),
.B2(n_37),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_94),
.B1(n_45),
.B2(n_35),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_166),
.B1(n_116),
.B2(n_176),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_141),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_127),
.C(n_124),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_0),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_180),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_48),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_109),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_94),
.B1(n_25),
.B2(n_19),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_12),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_12),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_172),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_38),
.C(n_37),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_174),
.C(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_11),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_48),
.Y(n_174)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_179),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_123),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_178),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_11),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_11),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_181),
.B(n_183),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_182),
.A2(n_186),
.B(n_199),
.Y(n_221)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_184),
.B(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_194),
.C(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_119),
.C(n_140),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_155),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_136),
.B1(n_132),
.B2(n_143),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_201),
.A2(n_209),
.B1(n_212),
.B2(n_48),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_143),
.C(n_144),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_144),
.C(n_38),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_209),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_211),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_145),
.B1(n_104),
.B2(n_38),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_151),
.B1(n_147),
.B2(n_163),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_180),
.B(n_177),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_214),
.B(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_230),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_173),
.B(n_174),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_173),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_223),
.Y(n_259)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_157),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_188),
.C(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_145),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_211),
.B(n_201),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_207),
.B1(n_206),
.B2(n_193),
.Y(n_250)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_236),
.B(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_185),
.A2(n_1),
.B(n_2),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_213),
.B1(n_183),
.B2(n_181),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_10),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_186),
.B(n_10),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_38),
.B1(n_37),
.B2(n_89),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_256),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_188),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_245),
.C(n_260),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_237),
.A2(n_194),
.B1(n_210),
.B2(n_203),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_262),
.B1(n_240),
.B2(n_223),
.Y(n_273)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_248),
.B(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_1),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_235),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_89),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_217),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_265),
.B(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_271),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_228),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_274),
.C(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_227),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_216),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_217),
.B1(n_218),
.B2(n_215),
.Y(n_277)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_280),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_257),
.B(n_236),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_219),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_283),
.C(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_226),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_266),
.A2(n_247),
.B(n_249),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

AO221x1_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_232),
.B1(n_229),
.B2(n_251),
.C(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_274),
.B(n_230),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_224),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_290),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_295),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_267),
.B(n_214),
.Y(n_295)
);

XNOR2x2_ASAP7_75t_SL g297 ( 
.A(n_265),
.B(n_264),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_298),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_5),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_260),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_304),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_283),
.C(n_281),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_311),
.C(n_287),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_275),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_234),
.C(n_253),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_306),
.C(n_309),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_262),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_244),
.C(n_238),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_320),
.B1(n_15),
.B2(n_7),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_321),
.B(n_316),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_284),
.B(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_308),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_319),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_289),
.B1(n_297),
.B2(n_8),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_6),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_6),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_7),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_312),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_8),
.B(n_9),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_302),
.C(n_312),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_328),
.C(n_9),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_7),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_6),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_331),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_332),
.C(n_326),
.Y(n_335)
);

O2A1O1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_322),
.B(n_325),
.C(n_332),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.C(n_328),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_13),
.C(n_14),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);


endmodule