module fake_jpeg_15427_n_358 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_9),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_50),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_17),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_48),
.C(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_42),
.Y(n_88)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_29),
.B1(n_21),
.B2(n_34),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_29),
.B1(n_21),
.B2(n_34),
.Y(n_80)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_80),
.A2(n_84),
.B1(n_30),
.B2(n_38),
.Y(n_140)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_29),
.B1(n_21),
.B2(n_34),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_41),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_35),
.C(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g131 ( 
.A(n_91),
.Y(n_131)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

BUFx6f_ASAP7_75t_SL g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_105),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_107),
.Y(n_124)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_40),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_35),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_111),
.B1(n_68),
.B2(n_32),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_35),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_30),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_53),
.B1(n_55),
.B2(n_33),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_118),
.B1(n_137),
.B2(n_123),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_53),
.B1(n_55),
.B2(n_76),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_140),
.B1(n_86),
.B2(n_23),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_33),
.B1(n_76),
.B2(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_133),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_54),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_31),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_135),
.B(n_142),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_94),
.B1(n_82),
.B2(n_25),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_24),
.B1(n_39),
.B2(n_28),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_31),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_143),
.A2(n_159),
.B1(n_165),
.B2(n_126),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_92),
.B1(n_93),
.B2(n_68),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_127),
.B1(n_121),
.B2(n_129),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_15),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_38),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_0),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_155),
.B(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_32),
.B(n_93),
.C(n_56),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_25),
.B1(n_26),
.B2(n_23),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_125),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_91),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_54),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_37),
.B1(n_26),
.B2(n_22),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_0),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_37),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_168),
.B(n_10),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_45),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_27),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_133),
.C(n_142),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_174),
.C(n_176),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_51),
.C(n_118),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_135),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_184),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_179),
.B(n_182),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_148),
.B(n_169),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_183),
.A2(n_160),
.B1(n_167),
.B2(n_131),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_51),
.C(n_127),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_90),
.B(n_108),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_155),
.B(n_170),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_191),
.B(n_198),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_125),
.C(n_141),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_203),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_200),
.B(n_159),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_202),
.B(n_165),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_125),
.C(n_56),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_201),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_207),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_154),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_143),
.B1(n_146),
.B2(n_156),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_216),
.A2(n_191),
.B1(n_175),
.B2(n_39),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_150),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_217),
.Y(n_260)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_170),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_218),
.A2(n_222),
.B(n_225),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_182),
.B(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_228),
.B1(n_231),
.B2(n_183),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_181),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_224),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_177),
.B(n_192),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_187),
.Y(n_225)
);

NOR2x1_ASAP7_75t_R g226 ( 
.A(n_186),
.B(n_153),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_226),
.A2(n_190),
.B1(n_188),
.B2(n_176),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_171),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_233),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_180),
.B(n_122),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_232),
.C(n_233),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_131),
.B1(n_171),
.B2(n_122),
.Y(n_231)
);

NOR4xp25_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_90),
.C(n_122),
.D(n_108),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_39),
.Y(n_233)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_173),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_50),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_240),
.A2(n_255),
.B1(n_231),
.B2(n_222),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_242),
.A2(n_245),
.B1(n_251),
.B2(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_249),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_203),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_228),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_199),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_200),
.C(n_178),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.C(n_213),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_204),
.A2(n_175),
.B1(n_0),
.B2(n_103),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_90),
.C(n_95),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_39),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_36),
.Y(n_280)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_208),
.B1(n_226),
.B2(n_218),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_263),
.A2(n_276),
.B1(n_282),
.B2(n_260),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_208),
.B(n_219),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_272),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_273),
.C(n_277),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_SL g268 ( 
.A(n_245),
.B(n_210),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_251),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_210),
.B(n_220),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_216),
.C(n_215),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_227),
.B1(n_211),
.B2(n_3),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_99),
.C(n_95),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_257),
.C(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_27),
.C(n_36),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_248),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_275),
.B1(n_265),
.B2(n_278),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_291),
.B1(n_292),
.B2(n_238),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_259),
.B1(n_247),
.B2(n_256),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_263),
.A2(n_259),
.B1(n_256),
.B2(n_241),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_247),
.B1(n_246),
.B2(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_281),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_282),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_2),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_235),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_252),
.Y(n_300)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_305),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_273),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_267),
.C(n_277),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_306),
.C(n_312),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_254),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_313),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_246),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_315),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_271),
.C(n_266),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_258),
.C(n_36),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_312),
.C(n_288),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_316),
.A2(n_287),
.B1(n_296),
.B2(n_292),
.Y(n_320)
);

OR2x2_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_297),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_329),
.Y(n_335)
);

XNOR2x1_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_28),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_28),
.C(n_24),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_289),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_309),
.A2(n_293),
.B1(n_297),
.B2(n_36),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_28),
.B1(n_24),
.B2(n_9),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_310),
.B(n_4),
.Y(n_327)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_327),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_303),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_314),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_27),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_325),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_331),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_316),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_332),
.B(n_333),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_339),
.C(n_317),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_321),
.A2(n_6),
.B(n_8),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_6),
.B(n_8),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_319),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_19),
.C(n_50),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_342),
.B(n_343),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_335),
.A2(n_326),
.B(n_320),
.Y(n_344)
);

AOI322xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_346),
.A3(n_333),
.B1(n_334),
.B2(n_338),
.C1(n_24),
.C2(n_19),
.Y(n_347)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_347),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_349),
.B(n_350),
.Y(n_352)
);

AOI322xp5_ASAP7_75t_L g349 ( 
.A1(n_345),
.A2(n_19),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_16),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_340),
.C(n_10),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_340),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_351),
.B1(n_11),
.B2(n_16),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_6),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_11),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_357),
.B(n_17),
.CI(n_50),
.CON(n_358),
.SN(n_358)
);


endmodule