module real_aes_4375_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_92;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_98;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g206 ( .A(n_0), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_1), .B(n_100), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_2), .B(n_134), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_3), .A2(n_28), .B1(n_149), .B2(n_255), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_4), .A2(n_30), .B1(n_168), .B2(n_233), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_5), .A2(n_49), .B1(n_214), .B2(n_216), .Y(n_224) );
INVx1_ASAP7_75t_L g200 ( .A(n_6), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_7), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_8), .A2(n_16), .B1(n_561), .B2(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g544 ( .A(n_9), .Y(n_544) );
INVxp67_ASAP7_75t_L g571 ( .A(n_9), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_9), .B(n_59), .Y(n_603) );
INVx1_ASAP7_75t_L g204 ( .A(n_10), .Y(n_204) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_10), .Y(n_640) );
OA21x2_ASAP7_75t_L g91 ( .A1(n_11), .A2(n_53), .B(n_92), .Y(n_91) );
OA21x2_ASAP7_75t_L g193 ( .A1(n_11), .A2(n_53), .B(n_92), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_12), .B(n_529), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_13), .A2(n_51), .B1(n_214), .B2(n_216), .Y(n_213) );
NAND2xp33_ASAP7_75t_L g523 ( .A(n_14), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g197 ( .A(n_15), .Y(n_197) );
BUFx3_ASAP7_75t_L g627 ( .A(n_17), .Y(n_627) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_18), .Y(n_529) );
AO22x1_ASAP7_75t_L g125 ( .A1(n_19), .A2(n_62), .B1(n_126), .B2(n_130), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_20), .Y(n_152) );
AND2x2_ASAP7_75t_L g167 ( .A(n_21), .B(n_168), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_22), .A2(n_54), .B1(n_548), .B2(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g597 ( .A(n_23), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_24), .B(n_130), .Y(n_161) );
AOI22x1_ASAP7_75t_L g238 ( .A1(n_25), .A2(n_74), .B1(n_214), .B2(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g530 ( .A(n_26), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_26), .B(n_58), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_27), .B(n_241), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_29), .B(n_96), .Y(n_177) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_31), .Y(n_611) );
INVx1_ASAP7_75t_SL g620 ( .A(n_32), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_33), .B(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_33), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_34), .B(n_159), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_35), .A2(n_57), .B1(n_580), .B2(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g92 ( .A(n_36), .Y(n_92) );
AND2x4_ASAP7_75t_L g114 ( .A(n_37), .B(n_115), .Y(n_114) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_37), .Y(n_637) );
INVx2_ASAP7_75t_L g615 ( .A(n_38), .Y(n_615) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_39), .Y(n_103) );
INVx2_ASAP7_75t_L g219 ( .A(n_40), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_41), .A2(n_43), .B1(n_574), .B2(n_578), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_42), .A2(n_60), .B1(n_149), .B2(n_239), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g137 ( .A(n_44), .Y(n_137) );
AND2x2_ASAP7_75t_L g175 ( .A(n_45), .B(n_130), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_46), .A2(n_520), .B1(n_608), .B2(n_646), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_46), .Y(n_646) );
OA22x2_ASAP7_75t_L g534 ( .A1(n_47), .A2(n_59), .B1(n_529), .B2(n_533), .Y(n_534) );
INVx1_ASAP7_75t_L g557 ( .A(n_47), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_48), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_50), .B(n_89), .Y(n_88) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_52), .B(n_121), .Y(n_178) );
CKINVDCx14_ASAP7_75t_R g244 ( .A(n_55), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_56), .A2(n_63), .B1(n_586), .B2(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g546 ( .A(n_58), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_58), .B(n_555), .Y(n_606) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_58), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g558 ( .A1(n_59), .A2(n_65), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_61), .B(n_100), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_64), .A2(n_75), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g532 ( .A(n_65), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_65), .B(n_73), .Y(n_604) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_66), .Y(n_98) );
BUFx5_ASAP7_75t_L g101 ( .A(n_66), .Y(n_101) );
INVx1_ASAP7_75t_L g129 ( .A(n_66), .Y(n_129) );
INVx2_ASAP7_75t_L g208 ( .A(n_67), .Y(n_208) );
AOI21xp33_ASAP7_75t_SL g594 ( .A1(n_68), .A2(n_595), .B(n_596), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_69), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_SL g115 ( .A(n_70), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_71), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g95 ( .A(n_72), .B(n_96), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_73), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_76), .B(n_119), .Y(n_164) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_509), .B1(n_516), .B2(n_622), .C(n_638), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
OR2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_413), .Y(n_81) );
NAND4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_308), .C(n_349), .D(n_384), .Y(n_82) );
AOI211xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_140), .B(n_257), .C(n_279), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
OR2x2_ASAP7_75t_L g377 ( .A(n_85), .B(n_286), .Y(n_377) );
OR2x2_ASAP7_75t_L g398 ( .A(n_85), .B(n_277), .Y(n_398) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g259 ( .A(n_86), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g446 ( .A(n_86), .B(n_277), .Y(n_446) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_116), .Y(n_86) );
AND2x2_ASAP7_75t_L g274 ( .A(n_87), .B(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g294 ( .A(n_87), .Y(n_294) );
INVx2_ASAP7_75t_L g298 ( .A(n_87), .Y(n_298) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
NOR2x1_ASAP7_75t_L g112 ( .A(n_89), .B(n_113), .Y(n_112) );
INVx3_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_90), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx4_ASAP7_75t_L g122 ( .A(n_91), .Y(n_122) );
BUFx3_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
OAI21x1_ASAP7_75t_L g93 ( .A1(n_94), .A2(n_104), .B(n_112), .Y(n_93) );
AOI21xp5_ASAP7_75t_L g94 ( .A1(n_95), .A2(n_99), .B(n_102), .Y(n_94) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g169 ( .A(n_97), .Y(n_169) );
INVx1_ASAP7_75t_L g172 ( .A(n_97), .Y(n_172) );
INVx6_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx3_ASAP7_75t_L g107 ( .A(n_98), .Y(n_107) );
INVx2_ASAP7_75t_L g156 ( .A(n_98), .Y(n_156) );
INVx2_ASAP7_75t_L g160 ( .A(n_98), .Y(n_160) );
INVx2_ASAP7_75t_L g149 ( .A(n_100), .Y(n_149) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g109 ( .A(n_101), .Y(n_109) );
INVx2_ASAP7_75t_L g130 ( .A(n_101), .Y(n_130) );
INVx2_ASAP7_75t_L g215 ( .A(n_101), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_102), .A2(n_149), .B1(n_150), .B2(n_154), .Y(n_148) );
INVx4_ASAP7_75t_L g153 ( .A(n_102), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_102), .B(n_249), .Y(n_248) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_103), .Y(n_111) );
INVxp67_ASAP7_75t_L g173 ( .A(n_103), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_103), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_103), .B(n_200), .Y(n_199) );
INVx4_ASAP7_75t_L g203 ( .A(n_103), .Y(n_203) );
INVx3_ASAP7_75t_L g223 ( .A(n_103), .Y(n_223) );
INVx1_ASAP7_75t_L g237 ( .A(n_103), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_108), .B(n_110), .Y(n_104) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
INVx2_ASAP7_75t_L g217 ( .A(n_107), .Y(n_217) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g124 ( .A(n_111), .Y(n_124) );
INVx2_ASAP7_75t_SL g135 ( .A(n_111), .Y(n_135) );
INVxp67_ASAP7_75t_L g162 ( .A(n_111), .Y(n_162) );
INVx2_ASAP7_75t_L g183 ( .A(n_113), .Y(n_183) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g118 ( .A(n_114), .Y(n_118) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
INVx3_ASAP7_75t_L g250 ( .A(n_114), .Y(n_250) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_115), .Y(n_635) );
INVx2_ASAP7_75t_SL g275 ( .A(n_116), .Y(n_275) );
AND2x2_ASAP7_75t_L g401 ( .A(n_116), .B(n_294), .Y(n_401) );
OAI21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_123), .B(n_136), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_117), .A2(n_123), .B(n_136), .Y(n_347) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_118), .B(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g218 ( .A(n_120), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g182 ( .A(n_122), .Y(n_182) );
AOI21x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B(n_131), .Y(n_123) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g235 ( .A(n_129), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_130), .A2(n_159), .B1(n_202), .B2(n_205), .Y(n_201) );
AOI21x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_135), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_135), .B(n_178), .Y(n_179) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
NOR2xp67_ASAP7_75t_SL g243 ( .A(n_138), .B(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_139), .A2(n_147), .B(n_164), .Y(n_146) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_139), .A2(n_147), .B(n_164), .Y(n_271) );
AO21x1_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_185), .B(n_225), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_141), .A2(n_421), .B1(n_426), .B2(n_429), .Y(n_420) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g226 ( .A(n_144), .Y(n_226) );
INVx1_ASAP7_75t_L g375 ( .A(n_144), .Y(n_375) );
OR2x2_ASAP7_75t_L g459 ( .A(n_144), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g333 ( .A(n_145), .B(n_268), .Y(n_333) );
AND2x2_ASAP7_75t_L g475 ( .A(n_145), .B(n_460), .Y(n_475) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_165), .Y(n_145) );
AND2x2_ASAP7_75t_L g369 ( .A(n_146), .B(n_246), .Y(n_369) );
AND2x2_ASAP7_75t_L g383 ( .A(n_146), .B(n_262), .Y(n_383) );
OAI21x1_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_157), .B(n_163), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI22x1_ASAP7_75t_L g231 ( .A1(n_153), .A2(n_232), .B1(n_236), .B2(n_238), .Y(n_231) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_153), .Y(n_515) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_162), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_159), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g514 ( .A(n_160), .Y(n_514) );
AO31x2_ASAP7_75t_L g230 ( .A1(n_163), .A2(n_231), .A3(n_240), .B(n_243), .Y(n_230) );
AO31x2_ASAP7_75t_L g265 ( .A1(n_163), .A2(n_231), .A3(n_240), .B(n_243), .Y(n_265) );
AND2x2_ASAP7_75t_L g510 ( .A(n_163), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g264 ( .A(n_165), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g322 ( .A(n_165), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g329 ( .A(n_165), .B(n_265), .Y(n_329) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_174), .B(n_180), .Y(n_165) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_166), .A2(n_174), .B(n_180), .Y(n_284) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_173), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_168), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g239 ( .A(n_172), .Y(n_239) );
OAI21x1_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_179), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g184 ( .A(n_178), .Y(n_184) );
AOI21xp33_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_183), .B(n_184), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND3xp33_ASAP7_75t_SL g212 ( .A(n_183), .B(n_192), .C(n_203), .Y(n_212) );
NAND3xp33_ASAP7_75t_L g221 ( .A(n_183), .B(n_192), .C(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g395 ( .A(n_186), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g326 ( .A(n_187), .B(n_311), .Y(n_326) );
AND2x2_ASAP7_75t_L g379 ( .A(n_187), .B(n_274), .Y(n_379) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_209), .Y(n_187) );
AND2x2_ASAP7_75t_L g287 ( .A(n_188), .B(n_210), .Y(n_287) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g300 ( .A(n_189), .Y(n_300) );
INVx1_ASAP7_75t_L g315 ( .A(n_189), .Y(n_315) );
AND2x2_ASAP7_75t_L g336 ( .A(n_189), .B(n_275), .Y(n_336) );
AND2x2_ASAP7_75t_L g348 ( .A(n_189), .B(n_210), .Y(n_348) );
OR2x2_ASAP7_75t_L g358 ( .A(n_189), .B(n_347), .Y(n_358) );
INVxp67_ASAP7_75t_L g506 ( .A(n_189), .Y(n_506) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_194), .B(n_207), .Y(n_189) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_193), .B(n_250), .Y(n_249) );
NAND3xp33_ASAP7_75t_SL g194 ( .A(n_195), .B(n_198), .C(n_201), .Y(n_194) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_203), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
NOR2x1_ASAP7_75t_L g314 ( .A(n_210), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g340 ( .A(n_210), .Y(n_340) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_210), .Y(n_364) );
INVx1_ASAP7_75t_L g412 ( .A(n_210), .Y(n_412) );
AND2x2_ASAP7_75t_L g430 ( .A(n_210), .B(n_294), .Y(n_430) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_220), .Y(n_210) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_218), .Y(n_211) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g220 ( .A(n_221), .B(n_224), .Y(n_220) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g465 ( .A(n_225), .Y(n_465) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_245), .Y(n_227) );
INVx2_ASAP7_75t_L g268 ( .A(n_228), .Y(n_268) );
INVx1_ASAP7_75t_L g367 ( .A(n_228), .Y(n_367) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g321 ( .A(n_229), .Y(n_321) );
AND2x2_ASAP7_75t_L g342 ( .A(n_229), .B(n_305), .Y(n_342) );
AND2x2_ASAP7_75t_L g407 ( .A(n_229), .B(n_284), .Y(n_407) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g356 ( .A(n_230), .B(n_270), .Y(n_356) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_237), .B(n_249), .Y(n_253) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g460 ( .A(n_245), .Y(n_460) );
INVx2_ASAP7_75t_L g483 ( .A(n_245), .Y(n_483) );
INVx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_252), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_247), .B(n_252), .Y(n_262) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_256), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_263), .B(n_266), .C(n_276), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g477 ( .A(n_260), .B(n_462), .Y(n_477) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g269 ( .A(n_262), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g291 ( .A(n_262), .Y(n_291) );
INVx2_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_262), .B(n_425), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_263), .A2(n_416), .B(n_420), .Y(n_415) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g282 ( .A(n_265), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g390 ( .A(n_265), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_272), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g374 ( .A(n_268), .Y(n_374) );
AND2x2_ASAP7_75t_L g403 ( .A(n_268), .B(n_322), .Y(n_403) );
INVx1_ASAP7_75t_L g437 ( .A(n_269), .Y(n_437) );
INVx2_ASAP7_75t_L g496 ( .A(n_269), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_270), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g423 ( .A(n_270), .Y(n_423) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g323 ( .A(n_271), .Y(n_323) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_271), .Y(n_410) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2x1_ASAP7_75t_SL g453 ( .A(n_274), .B(n_348), .Y(n_453) );
INVx1_ASAP7_75t_L g301 ( .A(n_275), .Y(n_301) );
INVx1_ASAP7_75t_L g397 ( .A(n_275), .Y(n_397) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g427 ( .A(n_277), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_SL g498 ( .A(n_277), .B(n_400), .Y(n_498) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g418 ( .A(n_278), .B(n_419), .Y(n_418) );
OAI32xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_285), .A3(n_288), .B1(n_295), .B2(n_306), .Y(n_279) );
OAI22xp33_ASAP7_75t_SL g337 ( .A1(n_280), .A2(n_338), .B1(n_341), .B2(n_343), .Y(n_337) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx3_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
AND2x4_ASAP7_75t_L g500 ( .A(n_282), .B(n_369), .Y(n_500) );
AND2x2_ASAP7_75t_L g507 ( .A(n_282), .B(n_483), .Y(n_507) );
INVx1_ASAP7_75t_L g355 ( .A(n_283), .Y(n_355) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVxp67_ASAP7_75t_L g382 ( .A(n_284), .Y(n_382) );
INVx1_ASAP7_75t_L g425 ( .A(n_284), .Y(n_425) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_287), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g463 ( .A(n_287), .B(n_401), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_287), .B(n_301), .Y(n_489) );
INVx2_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g417 ( .A(n_289), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g479 ( .A(n_292), .Y(n_479) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g428 ( .A(n_293), .B(n_397), .Y(n_428) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_302), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g311 ( .A(n_298), .Y(n_311) );
AND2x2_ASAP7_75t_L g339 ( .A(n_298), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g361 ( .A(n_298), .B(n_358), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_298), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g466 ( .A(n_299), .Y(n_466) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g472 ( .A(n_300), .Y(n_472) );
AND2x2_ASAP7_75t_L g494 ( .A(n_300), .B(n_311), .Y(n_494) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVxp67_ASAP7_75t_L g388 ( .A(n_304), .Y(n_388) );
OR2x2_ASAP7_75t_L g444 ( .A(n_304), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g406 ( .A(n_305), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_306), .A2(n_491), .B(n_493), .C(n_495), .Y(n_490) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_316), .B(n_324), .C(n_337), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g393 ( .A(n_311), .Y(n_393) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g439 ( .A(n_314), .B(n_401), .Y(n_439) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp67_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_318), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_319), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g441 ( .A(n_319), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g451 ( .A(n_321), .Y(n_451) );
AND2x2_ASAP7_75t_L g508 ( .A(n_321), .B(n_383), .Y(n_508) );
BUFx3_ASAP7_75t_L g371 ( .A(n_322), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_322), .B(n_342), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_323), .B(n_390), .Y(n_462) );
OAI32xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .A3(n_330), .B1(n_332), .B2(n_334), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2x1_ASAP7_75t_L g482 ( .A(n_328), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g442 ( .A(n_329), .Y(n_442) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g487 ( .A(n_331), .Y(n_487) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
NAND2x2_ASAP7_75t_L g338 ( .A(n_335), .B(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_336), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g429 ( .A(n_336), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g399 ( .A(n_340), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_342), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_348), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g492 ( .A(n_346), .B(n_412), .Y(n_492) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g450 ( .A(n_348), .B(n_396), .Y(n_450) );
INVx1_ASAP7_75t_L g456 ( .A(n_348), .Y(n_456) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_348), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_357), .B1(n_359), .B2(n_365), .C(n_376), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g467 ( .A(n_352), .Y(n_467) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g501 ( .A(n_353), .B(n_502), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_355), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g419 ( .A(n_358), .Y(n_419) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g470 ( .A(n_364), .B(n_419), .Y(n_470) );
NAND3xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_370), .C(n_372), .Y(n_365) );
INVx2_ASAP7_75t_L g433 ( .A(n_366), .Y(n_433) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OR2x2_ASAP7_75t_L g436 ( .A(n_367), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_380), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_380), .A2(n_449), .B1(n_454), .B2(n_455), .C(n_457), .Y(n_448) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g454 ( .A(n_383), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_383), .B(n_442), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_391), .B1(n_394), .B2(n_402), .C(n_404), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .C(n_399), .Y(n_394) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_SL g497 ( .A1(n_398), .A2(n_498), .B1(n_499), .B2(n_501), .C(n_503), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g481 ( .A1(n_399), .A2(n_482), .B(n_484), .C(n_490), .Y(n_481) );
OR2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_403), .B(n_470), .Y(n_469) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_408), .B(n_411), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_447), .C(n_480), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_431), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g445 ( .A(n_425), .Y(n_445) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_429), .B(n_439), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B(n_438), .C(n_440), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_439), .A2(n_441), .B1(n_443), .B2(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_446), .A2(n_504), .B1(n_507), .B2(n_508), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_464), .C(n_471), .Y(n_447) );
AOI21xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_452), .Y(n_449) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .B(n_463), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_467), .B2(n_468), .C(n_469), .Y(n_464) );
INVx2_ASAP7_75t_L g486 ( .A(n_470), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_474), .C(n_479), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_478), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_475), .A2(n_485), .B1(n_487), .B2(n_488), .Y(n_484) );
INVxp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_497), .Y(n_480) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g493 ( .A(n_492), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g504 ( .A(n_492), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OA21x2_ASAP7_75t_L g650 ( .A1(n_511), .A2(n_651), .B(n_652), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
XOR2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_609), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_520), .B1(n_607), .B2(n_608), .Y(n_517) );
INVx1_ASAP7_75t_L g607 ( .A(n_518), .Y(n_607) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g608 ( .A(n_520), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_520), .A2(n_608), .B1(n_640), .B2(n_641), .Y(n_639) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2x1_ASAP7_75t_L g521 ( .A(n_522), .B(n_572), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_547), .C(n_560), .Y(n_522) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_535), .Y(n_525) );
AND2x4_ASAP7_75t_L g548 ( .A(n_526), .B(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g574 ( .A(n_526), .B(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g580 ( .A(n_526), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_534), .Y(n_526) );
INVx1_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_531), .Y(n_527) );
NAND2xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g533 ( .A(n_529), .Y(n_533) );
INVx3_ASAP7_75t_L g539 ( .A(n_529), .Y(n_539) );
NAND2xp33_ASAP7_75t_L g545 ( .A(n_529), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g559 ( .A(n_529), .Y(n_559) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_529), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_530), .B(n_557), .Y(n_556) );
INVxp67_ASAP7_75t_L g631 ( .A(n_530), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g570 ( .A1(n_532), .A2(n_559), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g562 ( .A(n_534), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g569 ( .A(n_534), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g588 ( .A(n_534), .Y(n_588) );
AND2x4_ASAP7_75t_L g552 ( .A(n_535), .B(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g589 ( .A(n_535), .B(n_587), .Y(n_589) );
AND2x2_ASAP7_75t_L g595 ( .A(n_535), .B(n_562), .Y(n_595) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g549 ( .A(n_537), .B(n_541), .Y(n_549) );
AND2x2_ASAP7_75t_L g565 ( .A(n_537), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g576 ( .A(n_537), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g581 ( .A(n_537), .B(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_539), .B(n_544), .Y(n_543) );
INVxp67_ASAP7_75t_L g555 ( .A(n_539), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g605 ( .A(n_540), .B(n_554), .C(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g577 ( .A(n_542), .Y(n_577) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AND2x4_ASAP7_75t_L g561 ( .A(n_549), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g586 ( .A(n_549), .B(n_587), .Y(n_586) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g578 ( .A(n_553), .B(n_575), .Y(n_578) );
AND2x4_ASAP7_75t_L g583 ( .A(n_553), .B(n_581), .Y(n_583) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_558), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_557), .Y(n_632) );
AND2x4_ASAP7_75t_L g587 ( .A(n_563), .B(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g601 ( .A(n_567), .Y(n_601) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_568), .Y(n_628) );
NAND4xp25_ASAP7_75t_SL g572 ( .A(n_573), .B(n_579), .C(n_584), .D(n_594), .Y(n_572) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g593 ( .A(n_576), .Y(n_593) );
INVx1_ASAP7_75t_L g582 ( .A(n_577), .Y(n_582) );
AND2x4_ASAP7_75t_L g591 ( .A(n_581), .B(n_587), .Y(n_591) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
AND2x4_ASAP7_75t_L g592 ( .A(n_587), .B(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AO21x2_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_605), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
XOR2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_616), .B2(n_617), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_620), .B2(n_621), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_620), .Y(n_621) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_633), .Y(n_624) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g643 ( .A(n_626), .B(n_633), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B(n_629), .C(n_632), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
OR2x2_ASAP7_75t_L g648 ( .A(n_634), .B(n_637), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_634), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_634), .B(n_636), .Y(n_652) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B1(n_642), .B2(n_644), .C1(n_647), .C2(n_649), .Y(n_638) );
INVx1_ASAP7_75t_L g641 ( .A(n_640), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
endmodule