module real_aes_7532_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_884;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_468;
wire n_746;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_756;
wire n_404;
wire n_598;
wire n_288;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_741;
wire n_314;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_SL g701 ( .A1(n_0), .A2(n_239), .B1(n_650), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_1), .A2(n_14), .B1(n_711), .B2(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g640 ( .A(n_2), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_3), .A2(n_120), .B1(n_509), .B2(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_4), .A2(n_57), .B1(n_422), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_5), .A2(n_15), .B1(n_566), .B2(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_6), .Y(n_860) );
INVx1_ASAP7_75t_L g871 ( .A(n_7), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_8), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_9), .A2(n_132), .B1(n_436), .B2(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_10), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_11), .A2(n_139), .B1(n_649), .B2(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_12), .A2(n_151), .B1(n_428), .B2(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_13), .A2(n_222), .B1(n_739), .B2(n_741), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_16), .A2(n_75), .B1(n_472), .B2(n_473), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_17), .Y(n_610) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_18), .A2(n_172), .B1(n_432), .B2(n_433), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_19), .Y(n_706) );
AOI222xp33_ASAP7_75t_L g822 ( .A1(n_20), .A2(n_92), .B1(n_146), .B2(n_585), .C1(n_678), .C2(n_756), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_21), .A2(n_108), .B1(n_388), .B2(n_391), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_22), .Y(n_857) );
INVxp67_ASAP7_75t_L g881 ( .A(n_23), .Y(n_881) );
XOR2x2_ASAP7_75t_L g883 ( .A(n_23), .B(n_884), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_24), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_25), .B(n_418), .Y(n_417) );
AO22x2_ASAP7_75t_L g311 ( .A1(n_26), .A2(n_93), .B1(n_312), .B2(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g839 ( .A(n_26), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_27), .A2(n_162), .B1(n_457), .B2(n_459), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_28), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_29), .Y(n_455) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_30), .A2(n_137), .B1(n_649), .B2(n_650), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_31), .A2(n_213), .B1(n_338), .B2(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_32), .A2(n_166), .B1(n_441), .B2(n_538), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_33), .A2(n_260), .B1(n_493), .B2(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_34), .A2(n_606), .B1(n_636), .B2(n_637), .Y(n_605) );
INVx1_ASAP7_75t_L g636 ( .A(n_34), .Y(n_636) );
INVx1_ASAP7_75t_L g528 ( .A(n_35), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_36), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_37), .A2(n_181), .B1(n_422), .B2(n_424), .Y(n_421) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_38), .A2(n_97), .B1(n_312), .B2(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g840 ( .A(n_38), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_39), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_40), .A2(n_134), .B1(n_348), .B2(n_425), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_41), .A2(n_269), .B1(n_415), .B2(n_560), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_42), .A2(n_168), .B1(n_501), .B2(n_538), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_43), .A2(n_287), .B(n_295), .C(n_841), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_44), .A2(n_90), .B1(n_388), .B2(n_815), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_45), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_46), .A2(n_116), .B1(n_399), .B2(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_47), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_48), .A2(n_96), .B1(n_399), .B2(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_49), .B(n_346), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_50), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_51), .A2(n_71), .B1(n_565), .B2(n_566), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_52), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_53), .A2(n_165), .B1(n_459), .B2(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_54), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_55), .A2(n_122), .B1(n_395), .B2(n_399), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g504 ( .A1(n_56), .A2(n_192), .B1(n_262), .B2(n_338), .C1(n_505), .C2(n_507), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_58), .A2(n_60), .B1(n_372), .B2(n_392), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_59), .A2(n_242), .B1(n_501), .B2(n_741), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_61), .Y(n_609) );
AOI22xp5_ASAP7_75t_SL g698 ( .A1(n_62), .A2(n_167), .B1(n_441), .B2(n_699), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_63), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_63), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_64), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_65), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_66), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_67), .A2(n_276), .B1(n_430), .B2(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_68), .B(n_893), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_69), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_70), .A2(n_196), .B1(n_432), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_72), .A2(n_185), .B1(n_428), .B2(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_73), .A2(n_200), .B1(n_428), .B2(n_430), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_74), .B(n_560), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_76), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_77), .A2(n_173), .B1(n_383), .B2(n_686), .Y(n_746) );
AOI22xp5_ASAP7_75t_SL g697 ( .A1(n_78), .A2(n_145), .B1(n_439), .B2(n_533), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_79), .Y(n_583) );
INVx1_ASAP7_75t_L g334 ( .A(n_80), .Y(n_334) );
AO22x2_ASAP7_75t_L g575 ( .A1(n_81), .A2(n_576), .B1(n_598), .B2(n_599), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_81), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_82), .A2(n_237), .B1(n_433), .B2(n_503), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_83), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_84), .A2(n_227), .B1(n_416), .B2(n_560), .Y(n_712) );
AOI211xp5_ASAP7_75t_L g776 ( .A1(n_85), .A2(n_585), .B(n_777), .C(n_781), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_86), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_87), .A2(n_228), .B1(n_819), .B2(n_820), .Y(n_818) );
AOI22xp5_ASAP7_75t_SL g643 ( .A1(n_88), .A2(n_152), .B1(n_533), .B2(n_538), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_89), .A2(n_153), .B1(n_436), .B2(n_437), .Y(n_760) );
INVx1_ASAP7_75t_L g541 ( .A(n_91), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_94), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_95), .Y(n_451) );
INVx1_ASAP7_75t_L g322 ( .A(n_98), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_99), .A2(n_205), .B1(n_393), .B2(n_400), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_100), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_101), .Y(n_627) );
INVx1_ASAP7_75t_L g293 ( .A(n_102), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_103), .B(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_104), .A2(n_155), .B1(n_366), .B2(n_437), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_105), .A2(n_135), .B1(n_383), .B2(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_106), .A2(n_204), .B1(n_428), .B2(n_537), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_107), .A2(n_141), .B1(n_540), .B2(n_789), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_109), .A2(n_189), .B1(n_461), .B2(n_554), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_110), .A2(n_142), .B1(n_366), .B2(n_372), .Y(n_365) );
INVx1_ASAP7_75t_L g290 ( .A(n_111), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_112), .A2(n_150), .B1(n_338), .B2(n_348), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_113), .A2(n_174), .B1(n_383), .B2(n_396), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_114), .A2(n_206), .B1(n_540), .B2(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_115), .B(n_415), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g887 ( .A(n_117), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_118), .A2(n_194), .B1(n_481), .B2(n_736), .Y(n_897) );
INVx1_ASAP7_75t_L g849 ( .A(n_119), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_121), .A2(n_161), .B1(n_424), .B2(n_498), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_123), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_124), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_125), .A2(n_177), .B1(n_385), .B2(n_596), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_126), .A2(n_258), .B1(n_366), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_127), .A2(n_211), .B1(n_392), .B2(n_479), .Y(n_690) );
XNOR2xp5_ASAP7_75t_L g547 ( .A(n_128), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_129), .B(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_130), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_131), .A2(n_247), .B1(n_479), .B2(n_482), .Y(n_478) );
AOI22xp5_ASAP7_75t_SL g302 ( .A1(n_133), .A2(n_303), .B1(n_403), .B2(n_404), .Y(n_302) );
INVx1_ASAP7_75t_L g404 ( .A(n_133), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_136), .A2(n_843), .B1(n_872), .B2(n_873), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_136), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_138), .A2(n_190), .B1(n_425), .B2(n_509), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_140), .A2(n_216), .B1(n_459), .B2(n_562), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_143), .A2(n_261), .B1(n_464), .B2(n_498), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_144), .A2(n_198), .B1(n_428), .B2(n_702), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_147), .B(n_496), .Y(n_779) );
INVx2_ASAP7_75t_L g294 ( .A(n_148), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_149), .A2(n_249), .B1(n_347), .B2(n_459), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_154), .A2(n_225), .B1(n_336), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_156), .A2(n_235), .B1(n_425), .B2(n_562), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_157), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_158), .A2(n_223), .B1(n_493), .B2(n_901), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_159), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_160), .A2(n_209), .B1(n_399), .B2(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g289 ( .A(n_163), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_163), .Y(n_833) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_164), .A2(n_234), .B1(n_312), .B2(n_316), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g774 ( .A(n_169), .Y(n_774) );
INVx1_ASAP7_75t_L g306 ( .A(n_170), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_171), .A2(n_203), .B1(n_439), .B2(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_175), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_176), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_178), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_179), .A2(n_263), .B1(n_537), .B2(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_180), .B(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_182), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_183), .Y(n_765) );
INVx1_ASAP7_75t_L g356 ( .A(n_184), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_186), .A2(n_208), .B1(n_379), .B2(n_383), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_187), .A2(n_264), .B1(n_481), .B2(n_491), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_188), .A2(n_254), .B1(n_436), .B2(n_437), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_191), .Y(n_442) );
AO22x2_ASAP7_75t_L g319 ( .A1(n_193), .A2(n_250), .B1(n_312), .B2(n_313), .Y(n_319) );
INVx1_ASAP7_75t_L g344 ( .A(n_195), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_197), .A2(n_256), .B1(n_507), .B2(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g800 ( .A(n_199), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_201), .A2(n_218), .B1(n_569), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g846 ( .A(n_202), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_207), .A2(n_277), .B1(n_347), .B2(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g869 ( .A(n_210), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_212), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_214), .A2(n_255), .B1(n_439), .B2(n_441), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_215), .A2(n_233), .B1(n_388), .B2(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_217), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g858 ( .A(n_219), .B(n_650), .Y(n_858) );
INVx1_ASAP7_75t_L g732 ( .A(n_220), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_221), .A2(n_251), .B1(n_400), .B2(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_224), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_226), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_229), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_230), .A2(n_238), .B1(n_392), .B2(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_231), .Y(n_680) );
INVx1_ASAP7_75t_L g728 ( .A(n_232), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_234), .B(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_236), .B(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_240), .A2(n_280), .B1(n_686), .B2(n_687), .Y(n_685) );
AOI22xp5_ASAP7_75t_SL g646 ( .A1(n_241), .A2(n_284), .B1(n_437), .B2(n_647), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_243), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_244), .A2(n_259), .B1(n_415), .B2(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_245), .Y(n_580) );
INVx1_ASAP7_75t_L g351 ( .A(n_246), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_248), .A2(n_266), .B1(n_476), .B2(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g836 ( .A(n_250), .Y(n_836) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_252), .A2(n_253), .B1(n_736), .B2(n_737), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_257), .Y(n_468) );
OA22x2_ASAP7_75t_L g666 ( .A1(n_265), .A2(n_667), .B1(n_668), .B2(n_693), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_265), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_267), .Y(n_654) );
INVx1_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_270), .Y(n_552) );
INVx1_ASAP7_75t_L g725 ( .A(n_271), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_272), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_273), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_274), .A2(n_285), .B1(n_338), .B2(n_554), .Y(n_729) );
INVx1_ASAP7_75t_L g724 ( .A(n_275), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_278), .Y(n_751) );
INVx1_ASAP7_75t_L g731 ( .A(n_279), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_281), .A2(n_446), .B1(n_485), .B2(n_486), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_281), .Y(n_485) );
OA22x2_ASAP7_75t_L g805 ( .A1(n_282), .A2(n_806), .B1(n_807), .B2(n_823), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_282), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_283), .Y(n_672) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_290), .Y(n_832) );
OA21x2_ASAP7_75t_L g879 ( .A1(n_291), .A2(n_831), .B(n_880), .Y(n_879) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_513), .B1(n_826), .B2(n_827), .C(n_828), .Y(n_295) );
INVx1_ASAP7_75t_L g826 ( .A(n_296), .Y(n_826) );
AOI22xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_487), .B1(n_511), .B2(n_512), .Y(n_296) );
INVx1_ASAP7_75t_L g511 ( .A(n_297), .Y(n_511) );
BUFx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI22xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_301), .B1(n_444), .B2(n_445), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OA22x2_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_405), .B1(n_406), .B2(n_443), .Y(n_301) );
INVx1_ASAP7_75t_L g443 ( .A(n_302), .Y(n_443) );
INVx2_ASAP7_75t_SL g403 ( .A(n_303), .Y(n_403) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_363), .Y(n_303) );
NOR3xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_327), .C(n_350), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_322), .B2(n_323), .Y(n_305) );
OAI21xp5_ASAP7_75t_SL g655 ( .A1(n_307), .A2(n_656), .B(n_657), .Y(n_655) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g450 ( .A(n_308), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g845 ( .A1(n_308), .A2(n_846), .B(n_847), .Y(n_845) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .Y(n_308) );
INVx2_ASAP7_75t_L g382 ( .A(n_309), .Y(n_382) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_315), .Y(n_309) );
AND2x2_ASAP7_75t_L g326 ( .A(n_310), .B(n_315), .Y(n_326) );
AND2x2_ASAP7_75t_L g371 ( .A(n_310), .B(n_342), .Y(n_371) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g331 ( .A(n_311), .B(n_315), .Y(n_331) );
AND2x2_ASAP7_75t_L g343 ( .A(n_311), .B(n_321), .Y(n_343) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_314), .Y(n_316) );
INVx2_ASAP7_75t_L g342 ( .A(n_315), .Y(n_342) );
INVx1_ASAP7_75t_L g402 ( .A(n_315), .Y(n_402) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_318), .B(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g393 ( .A(n_318), .B(n_371), .Y(n_393) );
AND2x6_ASAP7_75t_L g416 ( .A(n_318), .B(n_326), .Y(n_416) );
AND2x4_ASAP7_75t_L g420 ( .A(n_318), .B(n_382), .Y(n_420) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g333 ( .A(n_319), .Y(n_333) );
INVx1_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_319), .B(n_321), .Y(n_377) );
AND2x2_ASAP7_75t_L g332 ( .A(n_320), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g370 ( .A(n_321), .B(n_362), .Y(n_370) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g581 ( .A(n_324), .Y(n_581) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g454 ( .A(n_325), .Y(n_454) );
AND2x4_ASAP7_75t_L g385 ( .A(n_326), .B(n_332), .Y(n_385) );
AND2x2_ASAP7_75t_L g398 ( .A(n_326), .B(n_370), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g867 ( .A(n_326), .B(n_370), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_334), .B1(n_335), .B2(n_344), .C(n_345), .Y(n_327) );
OAI21xp33_ASAP7_75t_SL g727 ( .A1(n_328), .A2(n_728), .B(n_729), .Y(n_727) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g551 ( .A(n_329), .Y(n_551) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g410 ( .A(n_330), .Y(n_410) );
INVx4_ASAP7_75t_L g506 ( .A(n_330), .Y(n_506) );
BUFx3_ASAP7_75t_L g585 ( .A(n_330), .Y(n_585) );
INVx2_ASAP7_75t_L g707 ( .A(n_330), .Y(n_707) );
INVx2_ASAP7_75t_SL g853 ( .A(n_330), .Y(n_853) );
AND2x6_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g359 ( .A(n_331), .Y(n_359) );
AND2x4_ASAP7_75t_L g425 ( .A(n_331), .B(n_361), .Y(n_425) );
AND2x6_ASAP7_75t_L g381 ( .A(n_332), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g390 ( .A(n_332), .B(n_371), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g673 ( .A1(n_335), .A2(n_674), .B1(n_675), .B2(n_676), .C(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_337), .A2(n_852), .B1(n_853), .B2(n_854), .Y(n_851) );
INVx4_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g660 ( .A(n_338), .Y(n_660) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_339), .Y(n_464) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_339), .Y(n_526) );
BUFx2_ASAP7_75t_L g587 ( .A(n_339), .Y(n_587) );
BUFx4f_ASAP7_75t_SL g756 ( .A(n_339), .Y(n_756) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g349 ( .A(n_341), .Y(n_349) );
INVx1_ASAP7_75t_L g355 ( .A(n_342), .Y(n_355) );
AND2x4_ASAP7_75t_L g348 ( .A(n_343), .B(n_349), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_343), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g422 ( .A(n_343), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g467 ( .A(n_346), .Y(n_467) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx12f_ASAP7_75t_L g509 ( .A(n_348), .Y(n_509) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_348), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_356), .B2(n_357), .Y(n_350) );
OAI22xp5_ASAP7_75t_SL g652 ( .A1(n_352), .A2(n_581), .B1(n_653), .B2(n_654), .Y(n_652) );
INVx3_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g590 ( .A(n_353), .Y(n_590) );
INVx4_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g632 ( .A(n_354), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_354), .A2(n_357), .B1(n_731), .B2(n_732), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_354), .A2(n_454), .B1(n_849), .B2(n_850), .Y(n_848) );
AND2x2_ASAP7_75t_L g650 ( .A(n_355), .B(n_376), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_357), .A2(n_632), .B1(n_680), .B2(n_681), .Y(n_679) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_358), .A2(n_589), .B1(n_590), .B2(n_591), .Y(n_588) );
CKINVDCx16_ASAP7_75t_R g635 ( .A(n_358), .Y(n_635) );
OR2x6_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_386), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_378), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx4f_ASAP7_75t_SL g736 ( .A(n_368), .Y(n_736) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g436 ( .A(n_369), .Y(n_436) );
BUFx3_ASAP7_75t_L g538 ( .A(n_369), .Y(n_538) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_370), .B(n_371), .Y(n_803) );
AND2x4_ASAP7_75t_L g375 ( .A(n_371), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g608 ( .A1(n_373), .A2(n_440), .B1(n_609), .B2(n_610), .C(n_611), .Y(n_608) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx3_ASAP7_75t_L g437 ( .A(n_375), .Y(n_437) );
BUFx3_ASAP7_75t_L g491 ( .A(n_375), .Y(n_491) );
BUFx2_ASAP7_75t_L g540 ( .A(n_375), .Y(n_540) );
BUFx3_ASAP7_75t_L g702 ( .A(n_375), .Y(n_702) );
BUFx2_ASAP7_75t_SL g737 ( .A(n_375), .Y(n_737) );
INVx1_ASAP7_75t_L g865 ( .A(n_375), .Y(n_865) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x6_ASAP7_75t_L g401 ( .A(n_377), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_SL g481 ( .A(n_380), .Y(n_481) );
INVx5_ASAP7_75t_SL g537 ( .A(n_380), .Y(n_537) );
INVx4_ASAP7_75t_L g572 ( .A(n_380), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_380), .B(n_871), .Y(n_870) );
INVx11_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx11_ASAP7_75t_L g440 ( .A(n_381), .Y(n_440) );
INVx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g482 ( .A(n_384), .Y(n_482) );
INVx2_ASAP7_75t_L g493 ( .A(n_384), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_384), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_793) );
INVx2_ASAP7_75t_L g810 ( .A(n_384), .Y(n_810) );
OAI22xp5_ASAP7_75t_SL g859 ( .A1(n_384), .A2(n_429), .B1(n_860), .B2(n_861), .Y(n_859) );
INVx6_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g441 ( .A(n_385), .Y(n_441) );
BUFx3_ASAP7_75t_L g565 ( .A(n_385), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_394), .Y(n_386) );
BUFx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx3_ASAP7_75t_L g472 ( .A(n_389), .Y(n_472) );
INVx3_ASAP7_75t_L g614 ( .A(n_389), .Y(n_614) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_389), .Y(n_686) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
BUFx2_ASAP7_75t_SL g699 ( .A(n_390), .Y(n_699) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
INVx2_ASAP7_75t_L g474 ( .A(n_393), .Y(n_474) );
BUFx3_ASAP7_75t_L g501 ( .A(n_393), .Y(n_501) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_393), .Y(n_649) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx2_ASAP7_75t_L g476 ( .A(n_396), .Y(n_476) );
INVx5_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
INVx2_ASAP7_75t_L g503 ( .A(n_397), .Y(n_503) );
INVx3_ASAP7_75t_L g533 ( .A(n_397), .Y(n_533) );
INVx4_ASAP7_75t_L g570 ( .A(n_397), .Y(n_570) );
BUFx3_ASAP7_75t_L g902 ( .A(n_397), .Y(n_902) );
INVx8_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx4f_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
BUFx2_ASAP7_75t_L g741 ( .A(n_400), .Y(n_741) );
BUFx2_ASAP7_75t_L g812 ( .A(n_400), .Y(n_812) );
INVx6_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g535 ( .A(n_401), .Y(n_535) );
INVx1_ASAP7_75t_L g692 ( .A(n_401), .Y(n_692) );
INVx1_ASAP7_75t_SL g792 ( .A(n_401), .Y(n_792) );
INVx1_ASAP7_75t_L g423 ( .A(n_402), .Y(n_423) );
INVx4_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
XOR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_442), .Y(n_406) );
NAND3x1_ASAP7_75t_L g407 ( .A(n_408), .B(n_426), .C(n_434), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_413), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_411), .B(n_412), .Y(n_409) );
OAI222xp33_ASAP7_75t_L g462 ( .A1(n_410), .A2(n_463), .B1(n_465), .B2(n_466), .C1(n_467), .C2(n_468), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_410), .A2(n_528), .B(n_529), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_410), .A2(n_751), .B(n_752), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .C(n_421), .Y(n_413) );
INVx1_ASAP7_75t_L g558 ( .A(n_415), .Y(n_558) );
BUFx4f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g820 ( .A(n_416), .Y(n_820) );
BUFx2_ASAP7_75t_L g893 ( .A(n_416), .Y(n_893) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g496 ( .A(n_419), .Y(n_496) );
INVx2_ASAP7_75t_L g523 ( .A(n_419), .Y(n_523) );
INVx5_ASAP7_75t_L g560 ( .A(n_419), .Y(n_560) );
INVx4_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g458 ( .A(n_422), .Y(n_458) );
BUFx2_ASAP7_75t_L g498 ( .A(n_422), .Y(n_498) );
BUFx2_ASAP7_75t_L g562 ( .A(n_422), .Y(n_562) );
BUFx3_ASAP7_75t_L g711 ( .A(n_422), .Y(n_711) );
BUFx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_425), .Y(n_461) );
BUFx2_ASAP7_75t_SL g530 ( .A(n_425), .Y(n_530) );
BUFx2_ASAP7_75t_SL g753 ( .A(n_425), .Y(n_753) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_431), .Y(n_426) );
INVx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g596 ( .A(n_429), .Y(n_596) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
BUFx2_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
INVx1_ASAP7_75t_L g795 ( .A(n_439), .Y(n_795) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx4_ASAP7_75t_L g647 ( .A(n_440), .Y(n_647) );
INVx2_ASAP7_75t_SL g815 ( .A(n_440), .Y(n_815) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g486 ( .A(n_446), .Y(n_486) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_469), .Y(n_446) );
NOR2xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_462), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_451), .B1(n_452), .B2(n_455), .C(n_456), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_449), .A2(n_579), .B1(n_580), .B2(n_581), .Y(n_578) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g624 ( .A(n_450), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_452), .A2(n_624), .B1(n_671), .B2(n_672), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g777 ( .A1(n_452), .A2(n_778), .B(n_779), .C(n_780), .Y(n_777) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g726 ( .A(n_454), .Y(n_726) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
OAI222xp33_ASAP7_75t_L g626 ( .A1(n_463), .A2(n_467), .B1(n_551), .B2(n_627), .C1(n_628), .C2(n_629), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI21xp5_ASAP7_75t_SL g856 ( .A1(n_474), .A2(n_857), .B(n_858), .Y(n_856) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_478), .B(n_483), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g512 ( .A(n_487), .Y(n_512) );
XOR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_510), .Y(n_487) );
NAND4xp75_ASAP7_75t_L g488 ( .A(n_489), .B(n_494), .C(n_499), .D(n_504), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
AND2x2_ASAP7_75t_SL g494 ( .A(n_495), .B(n_497), .Y(n_494) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_501), .Y(n_617) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_503), .Y(n_612) );
INVx4_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI22xp5_ASAP7_75t_SL g658 ( .A1(n_506), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_658) );
BUFx2_ASAP7_75t_L g674 ( .A(n_506), .Y(n_674) );
INVx1_ASAP7_75t_L g785 ( .A(n_507), .Y(n_785) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx4f_ASAP7_75t_SL g678 ( .A(n_509), .Y(n_678) );
INVx1_ASAP7_75t_L g827 ( .A(n_513), .Y(n_827) );
AOI22xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_769), .B1(n_770), .B2(n_825), .Y(n_513) );
INVx1_ASAP7_75t_L g825 ( .A(n_514), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_600), .B2(n_768), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_542), .B2(n_543), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
XOR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_541), .Y(n_518) );
NAND4xp75_ASAP7_75t_SL g519 ( .A(n_520), .B(n_531), .C(n_536), .D(n_539), .Y(n_519) );
NOR2xp67_ASAP7_75t_SL g520 ( .A(n_521), .B(n_527), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .C(n_525), .Y(n_521) );
INVx1_ASAP7_75t_L g783 ( .A(n_526), .Y(n_783) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g745 ( .A(n_537), .Y(n_745) );
INVx1_ASAP7_75t_L g567 ( .A(n_538), .Y(n_567) );
BUFx2_ASAP7_75t_L g620 ( .A(n_538), .Y(n_620) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AO22x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_574), .B2(n_575), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND4xp75_ASAP7_75t_SL g548 ( .A(n_549), .B(n_563), .C(n_571), .D(n_573), .Y(n_548) );
NOR2xp67_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .Y(n_549) );
OAI21xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_552), .B(n_553), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .C(n_561), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_560), .Y(n_819) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_560), .Y(n_891) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
INVx1_ASAP7_75t_L g688 ( .A(n_565), .Y(n_688) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g740 ( .A(n_570), .Y(n_740) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g598 ( .A(n_576), .Y(n_598) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_577), .B(n_592), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_582), .C(n_588), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_581), .A2(n_623), .B1(n_624), .B2(n_625), .Y(n_622) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_586), .Y(n_582) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND4x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .C(n_595), .D(n_597), .Y(n_592) );
INVx1_ASAP7_75t_L g768 ( .A(n_600), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_663), .B2(n_767), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_604), .B1(n_638), .B2(n_662), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g637 ( .A(n_606), .Y(n_637) );
AND2x2_ASAP7_75t_SL g606 ( .A(n_607), .B(n_621), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_613), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_615), .B1(n_616), .B2(n_618), .C(n_619), .Y(n_613) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .C(n_630), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_624), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g662 ( .A(n_638), .Y(n_662) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
XNOR2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND3x1_ASAP7_75t_SL g641 ( .A(n_642), .B(n_645), .C(n_651), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx4_ASAP7_75t_L g790 ( .A(n_649), .Y(n_790) );
NOR3xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .C(n_658), .Y(n_651) );
INVx1_ASAP7_75t_L g767 ( .A(n_663), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_715), .B2(n_716), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_694), .B1(n_695), .B2(n_714), .Y(n_665) );
INVx1_ASAP7_75t_L g714 ( .A(n_666), .Y(n_714) );
INVx1_ASAP7_75t_L g693 ( .A(n_668), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_682), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .C(n_679), .Y(n_669) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_683), .B(n_689), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_SL g799 ( .A(n_686), .Y(n_799) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
XOR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_713), .Y(n_695) );
NAND4xp75_ASAP7_75t_SL g696 ( .A(n_697), .B(n_698), .C(n_700), .D(n_704), .Y(n_696) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_709), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B(n_708), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AO22x1_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_747), .B2(n_766), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_733), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .C(n_730), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_742), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_738), .Y(n_734) );
INVx3_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_746), .Y(n_742) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_SL g766 ( .A(n_747), .Y(n_766) );
XOR2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_765), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_749), .B(n_758), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_754), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_804), .B1(n_805), .B2(n_824), .Y(n_770) );
INVx1_ASAP7_75t_SL g824 ( .A(n_771), .Y(n_824) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
XNOR2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
AND2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_786), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B1(n_784), .B2(n_785), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_793), .C(n_797), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
INVx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_803), .B(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_SL g823 ( .A(n_807), .Y(n_823) );
NAND4xp75_ASAP7_75t_L g807 ( .A(n_808), .B(n_813), .C(n_817), .D(n_822), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_811), .Y(n_808) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
AND2x2_ASAP7_75t_SL g817 ( .A(n_818), .B(n_821), .Y(n_817) );
INVx1_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
NOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_834), .Y(n_829) );
OR2x2_ASAP7_75t_SL g906 ( .A(n_830), .B(n_835), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_831), .Y(n_875) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_832), .B(n_878), .Y(n_880) );
CKINVDCx16_ASAP7_75t_R g878 ( .A(n_833), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
OAI322xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_874), .A3(n_876), .B1(n_879), .B2(n_881), .C1(n_882), .C2(n_904), .Y(n_841) );
INVx1_ASAP7_75t_L g873 ( .A(n_843), .Y(n_873) );
AND3x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_855), .C(n_862), .Y(n_843) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .C(n_851), .Y(n_844) );
OAI21xp5_ASAP7_75t_SL g886 ( .A1(n_853), .A2(n_887), .B(n_888), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_859), .Y(n_855) );
NOR3xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_868), .C(n_870), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_863) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_SL g884 ( .A(n_885), .B(n_895), .Y(n_884) );
NOR2xp33_ASAP7_75t_SL g885 ( .A(n_886), .B(n_889), .Y(n_885) );
NAND3xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .C(n_894), .Y(n_889) );
NOR2x1_ASAP7_75t_L g895 ( .A(n_896), .B(n_899), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_903), .Y(n_899) );
INVx3_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_905), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_906), .Y(n_905) );
endmodule