module fake_jpeg_3576_n_245 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_13),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_62),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_44),
.B(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_46),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_0),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_29),
.Y(n_55)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_25),
.B(n_10),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_18),
.A2(n_32),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_61),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_10),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_13),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_70),
.Y(n_116)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_76),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_73),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_49),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_25),
.B1(n_33),
.B2(n_27),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_106),
.B1(n_116),
.B2(n_115),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_39),
.B1(n_33),
.B2(n_27),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_42),
.A2(n_39),
.B1(n_30),
.B2(n_7),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_2),
.B1(n_6),
.B2(n_8),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_41),
.A2(n_6),
.B1(n_80),
.B2(n_78),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_111),
.B1(n_113),
.B2(n_81),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_117),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_47),
.B1(n_38),
.B2(n_46),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_47),
.A2(n_38),
.B1(n_46),
.B2(n_21),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_41),
.B(n_45),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_116),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_127),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_122),
.B(n_138),
.Y(n_162)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_132),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_134),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_137),
.B1(n_106),
.B2(n_149),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_136),
.Y(n_175)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_87),
.B1(n_117),
.B2(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_83),
.B(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_143),
.Y(n_159)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_110),
.C(n_99),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_146),
.B(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_150),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_84),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_107),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_127),
.C(n_121),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_177),
.B1(n_179),
.B2(n_175),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_102),
.B1(n_103),
.B2(n_94),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_140),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_102),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_169),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_123),
.B1(n_131),
.B2(n_147),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_174),
.B1(n_168),
.B2(n_158),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_145),
.B(n_148),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_166),
.B(n_177),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_125),
.B(n_147),
.C(n_150),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_193),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_126),
.B(n_143),
.C(n_144),
.D(n_161),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_190),
.B(n_196),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_158),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_166),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_168),
.B1(n_174),
.B2(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_170),
.CI(n_174),
.CON(n_191),
.SN(n_191)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_192),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_159),
.B(n_165),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_195),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_168),
.B1(n_174),
.B2(n_158),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_190),
.B1(n_181),
.B2(n_182),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_189),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_197),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_212),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_R g213 ( 
.A(n_201),
.B(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_214),
.Y(n_223)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_196),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_207),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_186),
.C(n_188),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_227),
.B(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_232),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_208),
.B1(n_211),
.B2(n_219),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_218),
.B1(n_211),
.B2(n_216),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_231),
.A2(n_203),
.B1(n_204),
.B2(n_182),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_236),
.B(n_225),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_226),
.B(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_225),
.C(n_222),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_239),
.B(n_236),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.C(n_224),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_238),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_243),
.B(n_184),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_235),
.Y(n_245)
);


endmodule