module fake_jpeg_20902_n_301 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx12f_ASAP7_75t_SL g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_44),
.Y(n_50)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_59),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_58),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_44),
.B(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_15),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_30),
.B1(n_22),
.B2(n_18),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_55),
.B1(n_51),
.B2(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_62),
.B(n_76),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_65),
.Y(n_104)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_42),
.B1(n_14),
.B2(n_26),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_73),
.B1(n_82),
.B2(n_87),
.Y(n_113)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g127 ( 
.A(n_70),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_44),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_23),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_14),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_84),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_16),
.B1(n_20),
.B2(n_25),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_31),
.B1(n_25),
.B2(n_27),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_91),
.B1(n_0),
.B2(n_1),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_43),
.B1(n_36),
.B2(n_39),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_36),
.C(n_39),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_0),
.C(n_1),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_20),
.B(n_27),
.C(n_28),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_24),
.B(n_22),
.C(n_11),
.Y(n_111)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_37),
.B1(n_28),
.B2(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_48),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_38),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_22),
.B(n_23),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_37),
.B1(n_32),
.B2(n_18),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_24),
.B1(n_19),
.B2(n_32),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_29),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_24),
.B1(n_19),
.B2(n_32),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_99),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_24),
.B1(n_32),
.B2(n_21),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_100),
.B1(n_102),
.B2(n_2),
.Y(n_135)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_24),
.B1(n_21),
.B2(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_40),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_103),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_24),
.B1(n_21),
.B2(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_40),
.B1(n_22),
.B2(n_23),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_129),
.B1(n_82),
.B2(n_87),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_29),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_122),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_22),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_118),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_72),
.B1(n_74),
.B2(n_99),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_63),
.B(n_0),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_73),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_137),
.A2(n_129),
.B1(n_100),
.B2(n_107),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_147),
.Y(n_177)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_142),
.Y(n_194)
);

AO21x2_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_113),
.B(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_143),
.B(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_75),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_106),
.B(n_71),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_150),
.B(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_76),
.B1(n_86),
.B2(n_61),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_68),
.B1(n_134),
.B2(n_119),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_153),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_85),
.B(n_76),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_156),
.A2(n_160),
.B(n_118),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_80),
.B1(n_83),
.B2(n_88),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_163),
.B1(n_122),
.B2(n_115),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_124),
.B1(n_66),
.B2(n_103),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_62),
.B(n_90),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_89),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_162),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_123),
.B1(n_113),
.B2(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_109),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_136),
.B1(n_142),
.B2(n_133),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_106),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_169),
.A2(n_185),
.B(n_186),
.Y(n_215)
);

AOI21x1_ASAP7_75t_SL g171 ( 
.A1(n_165),
.A2(n_62),
.B(n_135),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_157),
.B(n_154),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_182),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_181),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_183),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_118),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_147),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_144),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_188),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_125),
.B(n_90),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_192),
.B1(n_157),
.B2(n_139),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_193),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_97),
.B1(n_64),
.B2(n_65),
.Y(n_192)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_116),
.B(n_70),
.Y(n_193)
);

NAND2x1p5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_143),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_139),
.B1(n_143),
.B2(n_151),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_202),
.B1(n_205),
.B2(n_210),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_158),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_208),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_167),
.A2(n_143),
.B1(n_156),
.B2(n_155),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_189),
.B1(n_190),
.B2(n_170),
.Y(n_226)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_219),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_157),
.B1(n_161),
.B2(n_149),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_207),
.B1(n_174),
.B2(n_127),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_127),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_167),
.B1(n_169),
.B2(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_133),
.B1(n_127),
.B2(n_134),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_174),
.B1(n_193),
.B2(n_94),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_136),
.Y(n_214)
);

OAI221xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_172),
.B1(n_218),
.B2(n_175),
.C(n_184),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_127),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_153),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_193),
.B(n_172),
.Y(n_220)
);

OAI322xp33_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_2),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_181),
.B(n_186),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_229),
.Y(n_254)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_226),
.A2(n_228),
.B1(n_236),
.B2(n_239),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_190),
.B1(n_170),
.B2(n_173),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_180),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_218),
.B1(n_216),
.B2(n_207),
.Y(n_247)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_208),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_119),
.B1(n_117),
.B2(n_153),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_201),
.C(n_200),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_200),
.C(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_215),
.C(n_210),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_248),
.B1(n_256),
.B2(n_257),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_78),
.C(n_204),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_78),
.C(n_117),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_117),
.B1(n_11),
.B2(n_4),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_252),
.B1(n_242),
.B2(n_237),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_260),
.A2(n_269),
.B1(n_255),
.B2(n_239),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_261),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_233),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_264),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_254),
.A2(n_229),
.B(n_221),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_225),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_224),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_267),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_229),
.B1(n_231),
.B2(n_230),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_243),
.C(n_244),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_268),
.C(n_241),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_258),
.Y(n_286)
);

OAI321xp33_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_252),
.A3(n_247),
.B1(n_231),
.B2(n_253),
.C(n_236),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_279),
.B(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_270),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_SL g280 ( 
.A(n_278),
.B(n_264),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_284),
.B(n_273),
.Y(n_291)
);

AO21x2_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_260),
.B(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_282),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_268),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_274),
.B(n_95),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_286),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_295),
.A2(n_289),
.B(n_274),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_290),
.B(n_281),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_296),
.B(n_283),
.Y(n_299)
);

AOI321xp33_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_7),
.Y(n_301)
);


endmodule