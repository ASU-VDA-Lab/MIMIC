module fake_aes_4632_n_570 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_570);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_570;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_517;
wire n_560;
wire n_479;
wire n_554;
wire n_447;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_198;
wire n_424;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_43), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_31), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_91), .Y(n_180) );
BUFx10_ASAP7_75t_L g181 ( .A(n_92), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_157), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_62), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_116), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_13), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_56), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_75), .Y(n_189) );
INVx1_ASAP7_75t_SL g190 ( .A(n_60), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_13), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_153), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_61), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_144), .Y(n_194) );
INVx1_ASAP7_75t_SL g195 ( .A(n_16), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_148), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_107), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_73), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_131), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_145), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_147), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_97), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_89), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_19), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_52), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_11), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_105), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_81), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_167), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_117), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_161), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_152), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_27), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_55), .Y(n_214) );
INVx1_ASAP7_75t_SL g215 ( .A(n_57), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_42), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_135), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_7), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_9), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_68), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_29), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_15), .Y(n_222) );
NOR2xp67_ASAP7_75t_L g223 ( .A(n_136), .B(n_58), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_7), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_63), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_99), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_98), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_143), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_118), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_93), .Y(n_230) );
INVxp33_ASAP7_75t_R g231 ( .A(n_102), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_142), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_6), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_33), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_159), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_138), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_156), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_119), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_51), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_100), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_39), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_165), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_23), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_110), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_0), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_112), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_53), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_133), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_134), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_124), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_9), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_155), .Y(n_252) );
BUFx5_ASAP7_75t_L g253 ( .A(n_96), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_72), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_88), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_125), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_163), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_127), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_5), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_78), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_126), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_154), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_70), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_34), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_120), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_77), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_166), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_164), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_158), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_90), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_5), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_160), .Y(n_272) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_172), .A2(n_179), .B(n_173), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_181), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_235), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_181), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_240), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_247), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_255), .B(n_0), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_224), .Y(n_281) );
INVx4_ASAP7_75t_L g282 ( .A(n_178), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_185), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_191), .B(n_1), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_184), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_177), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_253), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_218), .Y(n_289) );
OAI22x1_ASAP7_75t_L g290 ( .A1(n_259), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_176), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_177), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_271), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_177), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_253), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_291), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_275), .B(n_214), .Y(n_298) );
NOR2xp33_ASAP7_75t_R g299 ( .A(n_275), .B(n_196), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_288), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_284), .Y(n_301) );
NAND2xp33_ASAP7_75t_R g302 ( .A(n_281), .B(n_233), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_293), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_287), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_282), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_277), .B(n_229), .Y(n_307) );
NOR2xp33_ASAP7_75t_R g308 ( .A(n_276), .B(n_193), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_283), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_282), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_278), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_279), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_274), .B(n_175), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_313), .B(n_280), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_306), .B(n_280), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g316 ( .A1(n_309), .A2(n_285), .B(n_274), .C(n_294), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_300), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_313), .B(n_303), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_303), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_310), .B(n_285), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_301), .B(n_289), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_304), .B(n_273), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_298), .B(n_273), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_307), .B(n_311), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_312), .Y(n_325) );
AND2x6_ASAP7_75t_SL g326 ( .A(n_297), .B(n_231), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_305), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_299), .B(n_186), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_308), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
NOR3xp33_ASAP7_75t_L g331 ( .A(n_311), .B(n_219), .C(n_245), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_306), .B(n_180), .Y(n_332) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_305), .B(n_194), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_318), .A2(n_321), .B1(n_323), .B2(n_314), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_319), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_317), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_322), .B(n_296), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_330), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_325), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_331), .A2(n_290), .B1(n_187), .B2(n_202), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_316), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_326), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_320), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_329), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_324), .B(n_251), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_328), .B(n_217), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_333), .B(n_2), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_331), .B(n_182), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_329), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_327), .B(n_200), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_332), .B(n_3), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_337), .A2(n_210), .B(n_207), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_334), .A2(n_195), .B1(n_215), .B2(n_190), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_344), .B(n_226), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_346), .B(n_192), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_335), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_339), .B(n_197), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_337), .A2(n_241), .B(n_239), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_336), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_343), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_341), .A2(n_243), .B(n_248), .C(n_246), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g363 ( .A1(n_351), .A2(n_254), .B(n_256), .C(n_252), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_345), .A2(n_261), .B(n_258), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_350), .B(n_199), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_203), .B1(n_204), .B2(n_201), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_348), .B(n_262), .Y(n_367) );
BUFx8_ASAP7_75t_L g368 ( .A(n_347), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_351), .A2(n_270), .B(n_265), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_349), .B(n_205), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_338), .A2(n_188), .B(n_174), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_340), .B(n_208), .Y(n_372) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_352), .A2(n_244), .B(n_257), .C(n_189), .Y(n_373) );
AOI22x1_ASAP7_75t_L g374 ( .A1(n_353), .A2(n_338), .B1(n_286), .B2(n_295), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_357), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_371), .A2(n_223), .B(n_253), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_368), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_361), .B(n_342), .Y(n_378) );
INVx8_ASAP7_75t_L g379 ( .A(n_368), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_372), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_367), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_362), .A2(n_253), .B(n_286), .Y(n_382) );
INVx4_ASAP7_75t_L g383 ( .A(n_358), .Y(n_383) );
INVx5_ASAP7_75t_L g384 ( .A(n_363), .Y(n_384) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_365), .B(n_356), .Y(n_385) );
OA21x2_ASAP7_75t_L g386 ( .A1(n_359), .A2(n_211), .B(n_209), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_354), .B(n_366), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_369), .A2(n_253), .B(n_286), .Y(n_388) );
BUFx12f_ASAP7_75t_L g389 ( .A(n_373), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_370), .B(n_198), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_371), .A2(n_249), .B(n_295), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_371), .A2(n_249), .B(n_295), .Y(n_393) );
BUFx10_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_371), .A2(n_249), .B(n_292), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_360), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_355), .Y(n_398) );
INVx8_ASAP7_75t_L g399 ( .A(n_355), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_355), .B(n_4), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_371), .A2(n_292), .B(n_14), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_357), .B(n_220), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g404 ( .A1(n_364), .A2(n_213), .B(n_212), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_368), .Y(n_405) );
NAND2x1p5_ASAP7_75t_L g406 ( .A(n_357), .B(n_242), .Y(n_406) );
CKINVDCx11_ASAP7_75t_R g407 ( .A(n_357), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_397), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_397), .Y(n_409) );
INVx3_ASAP7_75t_SL g410 ( .A(n_379), .Y(n_410) );
CKINVDCx6p67_ASAP7_75t_R g411 ( .A(n_379), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_399), .A2(n_268), .B1(n_263), .B2(n_216), .Y(n_412) );
INVx8_ASAP7_75t_L g413 ( .A(n_405), .Y(n_413) );
INVx5_ASAP7_75t_L g414 ( .A(n_377), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
BUFx12f_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_394), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_383), .B(n_6), .Y(n_420) );
BUFx12f_ASAP7_75t_L g421 ( .A(n_403), .Y(n_421) );
INVx4_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_380), .B(n_8), .Y(n_423) );
AOI21x1_ASAP7_75t_L g424 ( .A1(n_390), .A2(n_222), .B(n_221), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_396), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_396), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_388), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
INVx2_ASAP7_75t_SL g430 ( .A(n_385), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_393), .A2(n_227), .B(n_225), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_387), .A2(n_230), .B1(n_232), .B2(n_228), .Y(n_432) );
CKINVDCx6p67_ASAP7_75t_R g433 ( .A(n_384), .Y(n_433) );
BUFx4f_ASAP7_75t_SL g434 ( .A(n_391), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_382), .Y(n_436) );
AO21x1_ASAP7_75t_SL g437 ( .A1(n_374), .A2(n_18), .B(n_17), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_395), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_386), .A2(n_404), .B1(n_374), .B2(n_401), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_375), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_400), .B(n_8), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_389), .A2(n_272), .B1(n_269), .B2(n_267), .Y(n_442) );
OAI21x1_ASAP7_75t_L g443 ( .A1(n_392), .A2(n_21), .B(n_20), .Y(n_443) );
BUFx3_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_375), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_389), .A2(n_266), .B1(n_264), .B2(n_260), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_376), .A2(n_236), .B(n_234), .Y(n_447) );
CKINVDCx11_ASAP7_75t_R g448 ( .A(n_410), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_421), .Y(n_449) );
NAND2xp33_ASAP7_75t_R g450 ( .A(n_420), .B(n_10), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_444), .Y(n_451) );
NOR2xp33_ASAP7_75t_R g452 ( .A(n_411), .B(n_10), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_416), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_413), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_441), .B(n_12), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_430), .A2(n_22), .B(n_24), .C(n_25), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_408), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_423), .A2(n_250), .B1(n_238), .B2(n_237), .Y(n_458) );
NOR2xp33_ASAP7_75t_R g459 ( .A(n_413), .B(n_26), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_422), .B(n_28), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_409), .B(n_440), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_419), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_445), .B(n_30), .Y(n_463) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_412), .A2(n_32), .B(n_35), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_417), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_466) );
NOR2xp33_ASAP7_75t_R g467 ( .A(n_414), .B(n_40), .Y(n_467) );
NAND2xp33_ASAP7_75t_R g468 ( .A(n_418), .B(n_41), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_426), .Y(n_469) );
AO31x2_ASAP7_75t_L g470 ( .A1(n_436), .A2(n_44), .A3(n_45), .B(n_46), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_425), .Y(n_471) );
AND2x4_ASAP7_75t_SL g472 ( .A(n_433), .B(n_47), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_427), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_429), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_432), .B(n_170), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_429), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_435), .B(n_54), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_447), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_424), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_437), .A2(n_59), .B(n_64), .C(n_65), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_442), .B(n_66), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_446), .B(n_169), .Y(n_483) );
AO31x2_ASAP7_75t_L g484 ( .A1(n_428), .A2(n_67), .A3(n_69), .B(n_71), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_431), .Y(n_485) );
NOR3xp33_ASAP7_75t_SL g486 ( .A(n_439), .B(n_74), .C(n_76), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_443), .Y(n_487) );
NAND3xp33_ASAP7_75t_SL g488 ( .A(n_438), .B(n_79), .C(n_80), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_415), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_425), .B(n_82), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_460), .B(n_83), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_474), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_457), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_455), .B(n_84), .Y(n_495) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_472), .B(n_85), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_461), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_490), .B(n_86), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_477), .B(n_87), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_469), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_471), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_473), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_487), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_489), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_478), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_479), .B(n_94), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_451), .B(n_95), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_491), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_463), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_465), .B(n_101), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_459), .B(n_491), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_485), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_467), .Y(n_513) );
INVx5_ASAP7_75t_L g514 ( .A(n_449), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_484), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_480), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_452), .A2(n_103), .B1(n_104), .B2(n_106), .C(n_108), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_470), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_497), .B(n_486), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_494), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_501), .B(n_504), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_493), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_493), .B(n_454), .Y(n_524) );
NAND4xp25_ASAP7_75t_L g525 ( .A(n_511), .B(n_450), .C(n_468), .D(n_458), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_500), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_496), .A2(n_464), .B(n_476), .Y(n_527) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_492), .A2(n_475), .B1(n_483), .B2(n_482), .C(n_448), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_492), .A2(n_481), .B(n_488), .Y(n_529) );
OAI221xp5_ASAP7_75t_SL g530 ( .A1(n_507), .A2(n_462), .B1(n_456), .B2(n_466), .C(n_453), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_516), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_508), .B(n_109), .Y(n_532) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_515), .A2(n_111), .B(n_113), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_503), .B(n_114), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_503), .B(n_115), .Y(n_535) );
BUFx3_ASAP7_75t_L g536 ( .A(n_514), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_521), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_522), .B(n_502), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_523), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_526), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_531), .B(n_512), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_524), .B(n_505), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_536), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_524), .B(n_513), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_540), .Y(n_545) );
OAI32xp33_ASAP7_75t_L g546 ( .A1(n_539), .A2(n_525), .A3(n_527), .B1(n_520), .B2(n_532), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_541), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_537), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_543), .A2(n_530), .B(n_529), .C(n_528), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_544), .Y(n_550) );
AOI21xp33_ASAP7_75t_L g551 ( .A1(n_546), .A2(n_509), .B(n_510), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_549), .A2(n_514), .B(n_538), .C(n_542), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_547), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_545), .Y(n_554) );
OAI311xp33_ASAP7_75t_L g555 ( .A1(n_552), .A2(n_550), .A3(n_517), .B1(n_495), .C1(n_499), .Y(n_555) );
AOI21xp33_ASAP7_75t_SL g556 ( .A1(n_551), .A2(n_533), .B(n_548), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_556), .Y(n_557) );
AOI211x1_ASAP7_75t_L g558 ( .A1(n_557), .A2(n_554), .B(n_553), .C(n_555), .Y(n_558) );
NOR3x1_ASAP7_75t_L g559 ( .A(n_558), .B(n_498), .C(n_535), .Y(n_559) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_559), .B(n_534), .Y(n_560) );
AND4x2_ASAP7_75t_L g561 ( .A(n_560), .B(n_506), .C(n_121), .D(n_122), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_561), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_562), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_563), .A2(n_515), .B1(n_518), .B2(n_519), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_564), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_565), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_566), .B(n_123), .Y(n_567) );
AOI22xp5_ASAP7_75t_SL g568 ( .A1(n_567), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_568) );
OR2x6_ASAP7_75t_L g569 ( .A(n_568), .B(n_132), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_569), .A2(n_137), .B1(n_139), .B2(n_140), .Y(n_570) );
endmodule