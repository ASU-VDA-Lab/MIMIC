module real_aes_17282_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_853, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_853;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
AND2x4_ASAP7_75t_L g113 ( .A(n_0), .B(n_114), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_1), .A2(n_4), .B1(n_270), .B2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_2), .A2(n_43), .B1(n_151), .B2(n_243), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_3), .A2(n_23), .B1(n_211), .B2(n_243), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_5), .A2(n_16), .B1(n_183), .B2(n_185), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_6), .A2(n_61), .B1(n_147), .B2(n_213), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_7), .A2(n_17), .B1(n_151), .B2(n_156), .Y(n_509) );
INVx1_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_9), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_10), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_11), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_12), .A2(n_18), .B1(n_146), .B2(n_150), .Y(n_145) );
BUFx2_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
OR2x2_ASAP7_75t_L g132 ( .A(n_13), .B(n_38), .Y(n_132) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_14), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_15), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_19), .A2(n_101), .B1(n_183), .B2(n_270), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_20), .A2(n_39), .B1(n_175), .B2(n_177), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_21), .B(n_184), .Y(n_232) );
OAI21x1_ASAP7_75t_L g162 ( .A1(n_22), .A2(n_58), .B(n_163), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_24), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_25), .A2(n_54), .B1(n_135), .B2(n_136), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_25), .Y(n_135) );
INVx4_ASAP7_75t_R g534 ( .A(n_26), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_27), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_28), .B(n_154), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_29), .A2(n_47), .B1(n_196), .B2(n_199), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_30), .A2(n_53), .B1(n_183), .B2(n_199), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_31), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_32), .B(n_175), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_33), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_34), .B(n_243), .Y(n_577) );
INVx1_ASAP7_75t_L g616 ( .A(n_35), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_SL g552 ( .A1(n_36), .A2(n_151), .B(n_153), .C(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_37), .A2(n_55), .B1(n_151), .B2(n_199), .Y(n_561) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_38), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_40), .A2(n_87), .B1(n_151), .B2(n_210), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_41), .A2(n_80), .B1(n_835), .B2(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_41), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_42), .A2(n_46), .B1(n_151), .B2(n_156), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_44), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_45), .A2(n_59), .B1(n_183), .B2(n_197), .Y(n_272) );
INVx1_ASAP7_75t_L g574 ( .A(n_48), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_49), .B(n_151), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_50), .Y(n_593) );
INVx2_ASAP7_75t_L g124 ( .A(n_51), .Y(n_124) );
INVx1_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
BUFx3_ASAP7_75t_L g830 ( .A(n_52), .Y(n_830) );
INVx1_ASAP7_75t_L g136 ( .A(n_54), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_56), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_57), .A2(n_88), .B1(n_151), .B2(n_199), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g832 ( .A1(n_60), .A2(n_833), .B1(n_834), .B2(n_837), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_60), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_62), .A2(n_75), .B1(n_196), .B2(n_197), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_63), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_64), .A2(n_77), .B1(n_151), .B2(n_156), .Y(n_220) );
AOI21xp33_ASAP7_75t_R g841 ( .A1(n_65), .A2(n_486), .B(n_842), .Y(n_841) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_66), .A2(n_99), .B1(n_150), .B2(n_183), .Y(n_219) );
INVx1_ASAP7_75t_L g163 ( .A(n_67), .Y(n_163) );
AND2x4_ASAP7_75t_L g165 ( .A(n_68), .B(n_166), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_69), .A2(n_91), .B1(n_196), .B2(n_199), .Y(n_612) );
AO22x1_ASAP7_75t_L g521 ( .A1(n_70), .A2(n_76), .B1(n_177), .B2(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g166 ( .A(n_71), .Y(n_166) );
AND2x2_ASAP7_75t_L g555 ( .A(n_72), .B(n_238), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_73), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_74), .B(n_213), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_78), .B(n_243), .Y(n_594) );
INVx2_ASAP7_75t_L g154 ( .A(n_79), .Y(n_154) );
INVx1_ASAP7_75t_L g836 ( .A(n_80), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_81), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_82), .B(n_238), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_83), .A2(n_98), .B1(n_199), .B2(n_213), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_84), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_85), .B(n_161), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_86), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_89), .B(n_238), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_90), .A2(n_104), .B1(n_120), .B2(n_849), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_92), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_93), .B(n_238), .Y(n_590) );
INVx1_ASAP7_75t_L g112 ( .A(n_94), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_94), .B(n_492), .Y(n_491) );
NAND2xp33_ASAP7_75t_L g235 ( .A(n_95), .B(n_184), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_96), .A2(n_158), .B(n_213), .C(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g536 ( .A(n_97), .B(n_537), .Y(n_536) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_100), .A2(n_126), .B(n_482), .Y(n_125) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_100), .Y(n_484) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_102), .B(n_176), .Y(n_598) );
INVx5_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_115), .Y(n_105) );
OR2x6_ASAP7_75t_L g851 ( .A(n_106), .B(n_115), .Y(n_851) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NOR2x1p5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND3x2_ASAP7_75t_L g130 ( .A(n_108), .B(n_111), .C(n_131), .Y(n_130) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g492 ( .A(n_109), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g822 ( .A(n_112), .Y(n_822) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_125), .B(n_494), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
BUFx8_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g827 ( .A(n_124), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_124), .B(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_133), .Y(n_127) );
BUFx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_130), .B(n_484), .Y(n_483) );
AND2x6_ASAP7_75t_SL g490 ( .A(n_131), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_131), .B(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2x1_ASAP7_75t_L g848 ( .A(n_132), .B(n_830), .Y(n_848) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_133), .Y(n_485) );
XNOR2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_137), .Y(n_133) );
NAND4xp25_ASAP7_75t_L g137 ( .A(n_138), .B(n_357), .C(n_411), .D(n_450), .Y(n_137) );
NAND4xp75_ASAP7_75t_L g823 ( .A(n_138), .B(n_357), .C(n_411), .D(n_450), .Y(n_823) );
NOR2x1_ASAP7_75t_L g138 ( .A(n_139), .B(n_315), .Y(n_138) );
NAND3xp33_ASAP7_75t_SL g139 ( .A(n_140), .B(n_258), .C(n_297), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_205), .B1(n_248), .B2(n_253), .Y(n_140) );
INVx1_ASAP7_75t_L g421 ( .A(n_141), .Y(n_421) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_170), .Y(n_141) );
INVx1_ASAP7_75t_L g284 ( .A(n_142), .Y(n_284) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_SL g250 ( .A(n_143), .Y(n_250) );
AND2x2_ASAP7_75t_L g302 ( .A(n_143), .B(n_191), .Y(n_302) );
AND2x2_ASAP7_75t_L g341 ( .A(n_143), .B(n_172), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_143), .B(n_278), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_143), .B(n_477), .Y(n_476) );
AO31x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_159), .A3(n_164), .B(n_167), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_152), .B1(n_155), .B2(n_157), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_148), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g151 ( .A(n_149), .Y(n_151) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
INVx2_ASAP7_75t_L g211 ( .A(n_149), .Y(n_211) );
INVx1_ASAP7_75t_L g213 ( .A(n_149), .Y(n_213) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_149), .Y(n_243) );
INVx1_ASAP7_75t_L g271 ( .A(n_149), .Y(n_271) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g156 ( .A(n_151), .Y(n_156) );
INVx1_ASAP7_75t_L g197 ( .A(n_151), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_152), .A2(n_174), .B1(n_179), .B2(n_182), .Y(n_173) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_152), .A2(n_179), .B1(n_195), .B2(n_198), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_152), .A2(n_209), .B1(n_212), .B2(n_214), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_152), .A2(n_157), .B1(n_219), .B2(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_152), .A2(n_234), .B(n_235), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_152), .A2(n_179), .B1(n_242), .B2(n_244), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_152), .A2(n_179), .B1(n_269), .B2(n_272), .Y(n_268) );
OAI22x1_ASAP7_75t_L g508 ( .A1(n_152), .A2(n_214), .B1(n_509), .B2(n_510), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_152), .A2(n_517), .B1(n_560), .B2(n_561), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_152), .A2(n_214), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx6_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
O2A1O1Ixp5_ASAP7_75t_L g230 ( .A1(n_153), .A2(n_156), .B(n_231), .C(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_153), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_153), .A2(n_598), .B(n_599), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_153), .A2(n_516), .B(n_521), .C(n_524), .Y(n_637) );
BUFx8_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g158 ( .A(n_154), .Y(n_158) );
INVx2_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
INVx1_ASAP7_75t_L g551 ( .A(n_154), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_156), .A2(n_593), .B(n_594), .C(n_595), .Y(n_592) );
INVx1_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_159), .A2(n_218), .A3(n_221), .B(n_223), .Y(n_217) );
AOI21x1_ASAP7_75t_L g543 ( .A1(n_159), .A2(n_544), .B(n_555), .Y(n_543) );
AO31x2_ASAP7_75t_L g610 ( .A1(n_159), .A2(n_200), .A3(n_611), .B(n_615), .Y(n_610) );
BUFx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_160), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g537 ( .A(n_160), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_160), .B(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_160), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
INVx2_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
OAI21xp33_ASAP7_75t_L g524 ( .A1(n_161), .A2(n_519), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
AO31x2_ASAP7_75t_L g172 ( .A1(n_164), .A2(n_173), .A3(n_187), .B(n_189), .Y(n_172) );
INVx2_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_164), .A2(n_241), .A3(n_245), .B(n_246), .Y(n_240) );
AO31x2_ASAP7_75t_L g507 ( .A1(n_164), .A2(n_204), .A3(n_508), .B(n_511), .Y(n_507) );
BUFx10_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
INVx1_ASAP7_75t_L g525 ( .A(n_165), .Y(n_525) );
BUFx10_ASAP7_75t_L g562 ( .A(n_165), .Y(n_562) );
NOR2xp33_ASAP7_75t_SL g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx2_ASAP7_75t_L g193 ( .A(n_168), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_168), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OR2x2_ASAP7_75t_L g325 ( .A(n_171), .B(n_300), .Y(n_325) );
OR2x2_ASAP7_75t_L g367 ( .A(n_171), .B(n_347), .Y(n_367) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_191), .Y(n_171) );
INVx2_ASAP7_75t_L g252 ( .A(n_172), .Y(n_252) );
INVx1_ASAP7_75t_L g278 ( .A(n_172), .Y(n_278) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_172), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_172), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g432 ( .A(n_172), .Y(n_432) );
AND2x2_ASAP7_75t_L g437 ( .A(n_172), .B(n_266), .Y(n_437) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_176), .A2(n_186), .B1(n_534), .B2(n_535), .Y(n_533) );
OAI21xp33_ASAP7_75t_SL g570 ( .A1(n_177), .A2(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g517 ( .A(n_180), .Y(n_517) );
BUFx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g596 ( .A(n_181), .Y(n_596) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_184), .Y(n_522) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AO31x2_ASAP7_75t_L g207 ( .A1(n_187), .A2(n_200), .A3(n_208), .B(n_215), .Y(n_207) );
BUFx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_188), .B(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_188), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_SL g228 ( .A(n_188), .Y(n_228) );
INVx4_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_188), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g578 ( .A(n_188), .B(n_562), .Y(n_578) );
AND2x4_ASAP7_75t_L g251 ( .A(n_191), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g275 ( .A(n_191), .Y(n_275) );
INVx2_ASAP7_75t_L g324 ( .A(n_191), .Y(n_324) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_191), .Y(n_340) );
INVx1_ASAP7_75t_L g477 ( .A(n_191), .Y(n_477) );
AO31x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .A3(n_200), .B(n_202), .Y(n_191) );
AO31x2_ASAP7_75t_L g267 ( .A1(n_192), .A2(n_221), .A3(n_268), .B(n_273), .Y(n_267) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_192), .A2(n_528), .B(n_536), .Y(n_527) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_199), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g614 ( .A(n_199), .Y(n_614) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_SL g236 ( .A(n_201), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_204), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_225), .Y(n_205) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_206), .Y(n_305) );
AND2x2_ASAP7_75t_L g312 ( .A(n_206), .B(n_308), .Y(n_312) );
AND2x2_ASAP7_75t_L g369 ( .A(n_206), .B(n_356), .Y(n_369) );
AND2x4_ASAP7_75t_SL g478 ( .A(n_206), .B(n_280), .Y(n_478) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
BUFx2_ASAP7_75t_L g259 ( .A(n_207), .Y(n_259) );
OR2x2_ASAP7_75t_L g296 ( .A(n_207), .B(n_282), .Y(n_296) );
AND2x4_ASAP7_75t_L g309 ( .A(n_207), .B(n_257), .Y(n_309) );
INVx2_ASAP7_75t_L g337 ( .A(n_207), .Y(n_337) );
OR2x2_ASAP7_75t_L g363 ( .A(n_207), .B(n_240), .Y(n_363) );
INVx1_ASAP7_75t_L g416 ( .A(n_207), .Y(n_416) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_211), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_214), .B(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g257 ( .A(n_217), .Y(n_257) );
BUFx2_ASAP7_75t_L g335 ( .A(n_217), .Y(n_335) );
AND2x2_ASAP7_75t_L g423 ( .A(n_217), .B(n_337), .Y(n_423) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_222), .A2(n_529), .B(n_532), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_225), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
AND2x4_ASAP7_75t_L g336 ( .A(n_226), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g410 ( .A(n_226), .B(n_257), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_226), .B(n_259), .Y(n_428) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
BUFx2_ASAP7_75t_L g361 ( .A(n_227), .Y(n_361) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_263) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_233), .B(n_236), .Y(n_229) );
INVx2_ASAP7_75t_L g245 ( .A(n_238), .Y(n_245) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_238), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_239), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g281 ( .A(n_239), .Y(n_281) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_240), .Y(n_295) );
INVx1_ASAP7_75t_L g331 ( .A(n_240), .Y(n_331) );
AND2x2_ASAP7_75t_L g356 ( .A(n_240), .B(n_263), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_243), .B(n_547), .Y(n_546) );
AO31x2_ASAP7_75t_L g558 ( .A1(n_245), .A2(n_559), .A3(n_562), .B(n_563), .Y(n_558) );
AND2x2_ASAP7_75t_L g448 ( .A(n_248), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g481 ( .A(n_248), .B(n_346), .Y(n_481) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
INVx1_ASAP7_75t_L g444 ( .A(n_249), .Y(n_444) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x4_ASAP7_75t_L g276 ( .A(n_250), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g311 ( .A(n_250), .B(n_266), .Y(n_311) );
INVx1_ASAP7_75t_L g321 ( .A(n_250), .Y(n_321) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_250), .Y(n_328) );
INVx2_ASAP7_75t_L g353 ( .A(n_250), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_250), .B(n_275), .Y(n_366) );
OR2x2_ASAP7_75t_L g375 ( .A(n_250), .B(n_329), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_250), .B(n_323), .Y(n_385) );
AND2x2_ASAP7_75t_L g454 ( .A(n_250), .B(n_432), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_251), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g310 ( .A(n_251), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_251), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_251), .B(n_287), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_251), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g466 ( .A(n_251), .B(n_352), .Y(n_466) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_254), .A2(n_320), .B1(n_404), .B2(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_255), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g460 ( .A(n_256), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g480 ( .A(n_256), .B(n_356), .Y(n_480) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g292 ( .A(n_257), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_257), .B(n_281), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_257), .B(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_257), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B1(n_286), .B2(n_290), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_259), .B(n_261), .Y(n_348) );
NAND2x1_ASAP7_75t_L g409 ( .A(n_259), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g463 ( .A(n_259), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .B1(n_279), .B2(n_283), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_262), .Y(n_419) );
INVx1_ASAP7_75t_L g461 ( .A(n_262), .Y(n_461) );
INVx1_ASAP7_75t_L g282 ( .A(n_263), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_276), .Y(n_264) );
AOI211xp5_ASAP7_75t_L g349 ( .A1(n_265), .A2(n_350), .B(n_354), .C(n_355), .Y(n_349) );
INVx1_ASAP7_75t_L g387 ( .A(n_265), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_265), .B(n_341), .Y(n_425) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_275), .Y(n_265) );
INVx3_ASAP7_75t_L g347 ( .A(n_266), .Y(n_347) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g285 ( .A(n_267), .B(n_275), .Y(n_285) );
INVx2_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_271), .B(n_549), .Y(n_548) );
NAND2x1_ASAP7_75t_L g368 ( .A(n_276), .B(n_346), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_276), .B(n_339), .Y(n_378) );
INVx1_ASAP7_75t_L g407 ( .A(n_276), .Y(n_407) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_279), .A2(n_465), .B(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_280), .A2(n_299), .B(n_303), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_280), .B(n_434), .Y(n_470) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx3_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
AND2x4_ASAP7_75t_L g447 ( .A(n_285), .B(n_314), .Y(n_447) );
AND2x2_ASAP7_75t_L g453 ( .A(n_285), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g384 ( .A(n_287), .Y(n_384) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g304 ( .A(n_288), .B(n_295), .Y(n_304) );
AND2x2_ASAP7_75t_L g430 ( .A(n_288), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g301 ( .A(n_289), .Y(n_301) );
OR2x2_ASAP7_75t_L g351 ( .A(n_289), .B(n_324), .Y(n_351) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2x1p5_ASAP7_75t_L g362 ( .A(n_292), .B(n_363), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_292), .B(n_296), .Y(n_449) );
INVx1_ASAP7_75t_L g318 ( .A(n_293), .Y(n_318) );
NOR2x1_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp67_ASAP7_75t_SL g379 ( .A(n_296), .B(n_380), .Y(n_379) );
AOI222xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_305), .B1(n_306), .B2(n_310), .C1(n_312), .C2(n_313), .Y(n_297) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_299), .A2(n_343), .B(n_348), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_300), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g467 ( .A(n_300), .Y(n_467) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_301), .Y(n_473) );
AND2x4_ASAP7_75t_L g313 ( .A(n_302), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_302), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g457 ( .A(n_302), .Y(n_457) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
AND2x2_ASAP7_75t_L g398 ( .A(n_307), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g391 ( .A(n_308), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g330 ( .A(n_309), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_332), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B1(n_326), .B2(n_330), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_325), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g344 ( .A(n_322), .Y(n_344) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g380 ( .A(n_331), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_331), .B(n_336), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_331), .B(n_434), .Y(n_433) );
AOI211x1_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_338), .B(n_342), .C(n_349), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_333), .A2(n_447), .B(n_448), .Y(n_446) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g399 ( .A(n_335), .B(n_336), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_336), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_336), .Y(n_392) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g456 ( .A(n_339), .B(n_437), .Y(n_456) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g354 ( .A(n_341), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_341), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx4_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g374 ( .A(n_347), .B(n_366), .Y(n_374) );
OR2x2_ASAP7_75t_L g475 ( .A(n_347), .B(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_351), .Y(n_408) );
INVx2_ASAP7_75t_L g445 ( .A(n_351), .Y(n_445) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND5xp2_ASAP7_75t_L g451 ( .A(n_354), .B(n_404), .C(n_452), .D(n_455), .E(n_457), .Y(n_451) );
AND2x2_ASAP7_75t_L g422 ( .A(n_356), .B(n_423), .Y(n_422) );
NOR2x1_ASAP7_75t_L g357 ( .A(n_358), .B(n_395), .Y(n_357) );
NAND2xp67_ASAP7_75t_SL g358 ( .A(n_359), .B(n_376), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .B1(n_369), .B2(n_370), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NAND3xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .C(n_368), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
NAND3xp33_ASAP7_75t_SL g370 ( .A(n_371), .B(n_374), .C(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_SL g406 ( .A1(n_374), .A2(n_407), .B(n_408), .C(n_409), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B1(n_381), .B2(n_382), .C(n_386), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_383), .B(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_391), .B2(n_393), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g438 ( .A1(n_387), .A2(n_413), .B(n_439), .C(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g402 ( .A(n_388), .Y(n_402) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g427 ( .A(n_390), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g405 ( .A(n_399), .Y(n_405) );
AOI211xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_403), .C(n_406), .Y(n_400) );
AND3x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_438), .C(n_446), .Y(n_411) );
AOI221x1_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_420), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_433), .B2(n_436), .Y(n_426) );
INVx1_ASAP7_75t_L g440 ( .A(n_431), .Y(n_440) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
AOI211x1_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_458), .B(n_464), .C(n_479), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B1(n_474), .B2(n_478), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_486), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
CKINVDCx8_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
OAI331xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_824), .A3(n_831), .B1(n_838), .B2(n_839), .B3(n_841), .C1(n_853), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g840 ( .A(n_496), .Y(n_840) );
AO22x2_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_819), .B1(n_820), .B2(n_823), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
NOR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_733), .Y(n_498) );
NAND4xp75_ASAP7_75t_L g499 ( .A(n_500), .B(n_638), .C(n_680), .D(n_704), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI211xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_538), .B(n_579), .C(n_617), .Y(n_501) );
INVxp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g724 ( .A(n_504), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g818 ( .A(n_504), .B(n_755), .Y(n_818) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_513), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g633 ( .A(n_506), .B(n_589), .Y(n_633) );
AND2x2_ASAP7_75t_L g674 ( .A(n_506), .B(n_635), .Y(n_674) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g585 ( .A(n_507), .B(n_527), .Y(n_585) );
OR2x2_ASAP7_75t_L g603 ( .A(n_507), .B(n_527), .Y(n_603) );
INVx2_ASAP7_75t_L g625 ( .A(n_507), .Y(n_625) );
AND2x2_ASAP7_75t_L g655 ( .A(n_507), .B(n_589), .Y(n_655) );
AND2x2_ASAP7_75t_L g684 ( .A(n_507), .B(n_526), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_507), .B(n_636), .Y(n_720) );
AND2x2_ASAP7_75t_L g697 ( .A(n_513), .B(n_626), .Y(n_697) );
INVx2_ASAP7_75t_L g792 ( .A(n_513), .Y(n_792) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_526), .Y(n_513) );
INVx2_ASAP7_75t_L g584 ( .A(n_514), .Y(n_584) );
AND2x4_ASAP7_75t_L g623 ( .A(n_514), .B(n_527), .Y(n_623) );
AOI21x1_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_520), .B(n_523), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_517), .A2(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_525), .A2(n_545), .B(n_552), .Y(n_544) );
AND2x2_ASAP7_75t_L g782 ( .A(n_526), .B(n_584), .Y(n_782) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g646 ( .A(n_527), .Y(n_646) );
AND2x2_ASAP7_75t_L g703 ( .A(n_527), .B(n_589), .Y(n_703) );
AND2x2_ASAP7_75t_L g718 ( .A(n_527), .B(n_626), .Y(n_718) );
AND2x2_ASAP7_75t_L g740 ( .A(n_527), .B(n_584), .Y(n_740) );
OAI211xp5_ASAP7_75t_SL g787 ( .A1(n_538), .A2(n_788), .B(n_790), .C(n_797), .Y(n_787) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_565), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g774 ( .A(n_541), .B(n_710), .Y(n_774) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_556), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_542), .B(n_567), .Y(n_673) );
INVxp67_ASAP7_75t_L g687 ( .A(n_542), .Y(n_687) );
AND2x2_ASAP7_75t_L g707 ( .A(n_542), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_542), .B(n_620), .Y(n_714) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_548), .B(n_550), .Y(n_545) );
BUFx4f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_551), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g648 ( .A(n_556), .B(n_630), .Y(n_648) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g696 ( .A(n_557), .B(n_607), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_557), .B(n_610), .Y(n_702) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g606 ( .A(n_558), .B(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g671 ( .A(n_558), .B(n_610), .Y(n_671) );
BUFx2_ASAP7_75t_L g678 ( .A(n_558), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_558), .B(n_610), .Y(n_758) );
INVx1_ASAP7_75t_L g601 ( .A(n_562), .Y(n_601) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g688 ( .A(n_566), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g817 ( .A(n_566), .B(n_606), .Y(n_817) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g620 ( .A(n_567), .Y(n_620) );
AND2x2_ASAP7_75t_L g631 ( .A(n_567), .B(n_610), .Y(n_631) );
AND2x2_ASAP7_75t_L g677 ( .A(n_567), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g710 ( .A(n_567), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_567), .B(n_621), .Y(n_727) );
AND2x2_ASAP7_75t_L g766 ( .A(n_567), .B(n_767), .Y(n_766) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_575), .B(n_578), .Y(n_569) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_586), .B(n_604), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_581), .A2(n_745), .B1(n_746), .B2(n_748), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
AND2x2_ASAP7_75t_L g742 ( .A(n_582), .B(n_633), .Y(n_742) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g657 ( .A(n_583), .Y(n_657) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g806 ( .A(n_584), .B(n_626), .Y(n_806) );
AND2x2_ASAP7_75t_L g770 ( .A(n_585), .B(n_665), .Y(n_770) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_602), .Y(n_586) );
OR2x2_ASAP7_75t_L g667 ( .A(n_587), .B(n_644), .Y(n_667) );
OR2x2_ASAP7_75t_L g779 ( .A(n_587), .B(n_603), .Y(n_779) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g642 ( .A(n_588), .Y(n_642) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g626 ( .A(n_589), .Y(n_626) );
BUFx3_ASAP7_75t_L g708 ( .A(n_589), .Y(n_708) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_597), .B(n_600), .Y(n_591) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g776 ( .A(n_603), .B(n_635), .Y(n_776) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
AND2x2_ASAP7_75t_L g618 ( .A(n_606), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g659 ( .A(n_606), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g796 ( .A(n_606), .Y(n_796) );
INVx1_ASAP7_75t_L g815 ( .A(n_606), .Y(n_815) );
INVx2_ASAP7_75t_L g630 ( .A(n_607), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_607), .B(n_610), .Y(n_679) );
INVx1_ASAP7_75t_L g743 ( .A(n_608), .Y(n_743) );
BUFx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g804 ( .A(n_609), .Y(n_804) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g621 ( .A(n_610), .Y(n_621) );
INVx1_ASAP7_75t_L g711 ( .A(n_610), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_622), .B1(n_627), .B2(n_632), .Y(n_617) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g660 ( .A(n_620), .Y(n_660) );
AND2x2_ASAP7_75t_L g662 ( .A(n_620), .B(n_647), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_620), .B(n_630), .Y(n_722) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx3_ASAP7_75t_L g653 ( .A(n_623), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_623), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g747 ( .A(n_623), .B(n_731), .Y(n_747) );
INVx1_ASAP7_75t_L g651 ( .A(n_624), .Y(n_651) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_624), .A2(n_662), .B1(n_663), .B2(n_668), .C1(n_674), .C2(n_675), .Y(n_661) );
OAI21xp33_ASAP7_75t_SL g691 ( .A1(n_624), .A2(n_692), .B(n_693), .Y(n_691) );
AND2x2_ASAP7_75t_L g715 ( .A(n_624), .B(n_634), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_624), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
OR2x2_ASAP7_75t_L g644 ( .A(n_625), .B(n_636), .Y(n_644) );
INVx1_ASAP7_75t_L g732 ( .A(n_625), .Y(n_732) );
BUFx2_ASAP7_75t_L g666 ( .A(n_626), .Y(n_666) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_629), .B(n_670), .Y(n_699) );
OR2x2_ASAP7_75t_L g811 ( .A(n_629), .B(n_671), .Y(n_811) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g694 ( .A(n_631), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g809 ( .A(n_631), .Y(n_809) );
OAI31xp33_ASAP7_75t_L g790 ( .A1(n_632), .A2(n_791), .A3(n_793), .B(n_794), .Y(n_790) );
AND2x4_ASAP7_75t_SL g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_633), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_661), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_647), .B(n_649), .Y(n_639) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x6_ASAP7_75t_L g760 ( .A(n_642), .B(n_761), .Y(n_760) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g692 ( .A(n_645), .Y(n_692) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g783 ( .A(n_646), .B(n_720), .Y(n_783) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_648), .A2(n_737), .B1(n_739), .B2(n_741), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_648), .A2(n_709), .B(n_771), .C(n_798), .Y(n_797) );
AOI21xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_654), .B(n_658), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g750 ( .A(n_653), .B(n_751), .C(n_752), .D(n_754), .Y(n_750) );
NAND2x1_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_655), .B(n_657), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_655), .B(n_740), .Y(n_763) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g729 ( .A(n_660), .B(n_689), .Y(n_729) );
NAND2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_667), .A2(n_811), .B1(n_812), .B2(n_814), .Y(n_810) );
AOI221x1_ASAP7_75t_L g749 ( .A1(n_668), .A2(n_750), .B1(n_756), .B2(n_759), .C(n_762), .Y(n_749) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g689 ( .A(n_671), .Y(n_689) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g701 ( .A(n_673), .B(n_702), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g764 ( .A(n_674), .B(n_755), .Y(n_764) );
O2A1O1Ixp5_ASAP7_75t_L g777 ( .A1(n_675), .A2(n_759), .B(n_778), .C(n_780), .Y(n_777) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx2_ASAP7_75t_L g726 ( .A(n_678), .Y(n_726) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_690), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g769 ( .A1(n_682), .A2(n_700), .B1(n_770), .B2(n_771), .C(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g706 ( .A(n_684), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_684), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g805 ( .A(n_684), .B(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
NAND2x1_ASAP7_75t_L g784 ( .A(n_687), .B(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g808 ( .A(n_687), .B(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g748 ( .A(n_688), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_694), .B1(n_697), .B2(n_698), .C1(n_700), .C2(n_703), .Y(n_690) );
INVx1_ASAP7_75t_L g775 ( .A(n_694), .Y(n_775) );
INVx1_ASAP7_75t_L g738 ( .A(n_695), .Y(n_738) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g772 ( .A(n_696), .Y(n_772) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g713 ( .A(n_702), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g767 ( .A(n_702), .Y(n_767) );
AND2x2_ASAP7_75t_L g730 ( .A(n_703), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_723), .Y(n_704) );
AOI222xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B1(n_712), .B2(n_715), .C1(n_716), .C2(n_721), .Y(n_705) );
INVx3_ASAP7_75t_L g755 ( .A(n_708), .Y(n_755) );
BUFx2_ASAP7_75t_L g813 ( .A(n_708), .Y(n_813) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g785 ( .A(n_710), .Y(n_785) );
OR2x2_ASAP7_75t_L g795 ( .A(n_710), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx2_ASAP7_75t_SL g753 ( .A(n_718), .Y(n_753) );
AND2x2_ASAP7_75t_L g798 ( .A(n_719), .B(n_755), .Y(n_798) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_720), .Y(n_751) );
INVxp67_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g757 ( .A(n_722), .B(n_758), .Y(n_757) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_728), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
OR2x2_ASAP7_75t_L g814 ( .A(n_727), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g745 ( .A(n_729), .Y(n_745) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g752 ( .A(n_732), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g802 ( .A(n_732), .Y(n_802) );
NAND4xp75_ASAP7_75t_L g733 ( .A(n_734), .B(n_768), .C(n_786), .D(n_799), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_749), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_743), .B(n_744), .Y(n_735) );
INVxp33_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_738), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g761 ( .A(n_740), .Y(n_761) );
AND2x2_ASAP7_75t_L g801 ( .A(n_740), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g771 ( .A(n_743), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g789 ( .A(n_754), .Y(n_789) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OAI22xp33_ASAP7_75t_SL g780 ( .A1(n_757), .A2(n_781), .B1(n_783), .B2(n_784), .Y(n_780) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI21xp33_ASAP7_75t_SL g762 ( .A1(n_763), .A2(n_764), .B(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g793 ( .A(n_764), .Y(n_793) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_777), .Y(n_768) );
AOI21xp5_ASAP7_75t_SL g773 ( .A1(n_774), .A2(n_775), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_816), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_803), .B1(n_805), .B2(n_807), .C(n_810), .Y(n_800) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx12f_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
AND2x2_ASAP7_75t_L g847 ( .A(n_822), .B(n_848), .Y(n_847) );
CKINVDCx16_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
BUFx12f_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND2x6_ASAP7_75t_SL g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
CKINVDCx6p67_ASAP7_75t_R g838 ( .A(n_831), .Y(n_838) );
BUFx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
BUFx10_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
CKINVDCx8_ASAP7_75t_R g849 ( .A(n_850), .Y(n_849) );
CKINVDCx10_ASAP7_75t_R g850 ( .A(n_851), .Y(n_850) );
endmodule