module real_jpeg_18860_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_578;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_313;
wire n_42;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_625;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_625),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_0),
.B(n_626),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_2),
.Y(n_159)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_2),
.Y(n_198)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_3),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_4),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_4),
.A2(n_152),
.B1(n_236),
.B2(n_240),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_4),
.A2(n_152),
.B1(n_354),
.B2(n_357),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_4),
.A2(n_152),
.B1(n_174),
.B2(n_571),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_5),
.A2(n_57),
.B1(n_187),
.B2(n_191),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_5),
.A2(n_57),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_5),
.A2(n_57),
.B1(n_135),
.B2(n_562),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_6),
.B(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_6),
.A2(n_132),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_6),
.B(n_120),
.Y(n_427)
);

OAI32xp33_ASAP7_75t_L g430 ( 
.A1(n_6),
.A2(n_431),
.A3(n_433),
.B1(n_436),
.B2(n_438),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_6),
.A2(n_321),
.B1(n_354),
.B2(n_450),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_6),
.A2(n_139),
.B1(n_516),
.B2(n_521),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_7),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_7),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g472 ( 
.A(n_7),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_7),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_8),
.A2(n_81),
.B1(n_258),
.B2(n_261),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_8),
.A2(n_81),
.B1(n_317),
.B2(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_8),
.A2(n_81),
.B1(n_216),
.B2(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_9),
.A2(n_172),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_9),
.A2(n_180),
.B1(n_279),
.B2(n_284),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_9),
.A2(n_180),
.B1(n_408),
.B2(n_411),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_9),
.A2(n_180),
.B1(n_499),
.B2(n_501),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_10),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

BUFx4f_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_11),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_11),
.A2(n_175),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_11),
.A2(n_175),
.B1(n_402),
.B2(n_405),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_11),
.A2(n_175),
.B1(n_517),
.B2(n_519),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_12),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_12),
.A2(n_63),
.B1(n_191),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_12),
.A2(n_63),
.B1(n_376),
.B2(n_379),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_12),
.A2(n_63),
.B1(n_308),
.B2(n_584),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_13),
.A2(n_217),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_13),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_13),
.A2(n_248),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_13),
.A2(n_248),
.B1(n_313),
.B2(n_317),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_13),
.A2(n_248),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_14),
.Y(n_626)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_16),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_16),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_16),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_16),
.Y(n_404)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_16),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_16),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_17),
.A2(n_150),
.B1(n_161),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_17),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_17),
.A2(n_166),
.B1(n_216),
.B2(n_221),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_17),
.A2(n_166),
.B1(n_266),
.B2(n_372),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_17),
.A2(n_166),
.B1(n_347),
.B2(n_580),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_18),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_18),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_18),
.A2(n_116),
.B1(n_240),
.B2(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_18),
.A2(n_116),
.B1(n_347),
.B2(n_350),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_18),
.A2(n_116),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g179 ( 
.A(n_19),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_69),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_68),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_64),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_24),
.B(n_617),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_24),
.B(n_617),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_46),
.B1(n_58),
.B2(n_59),
.Y(n_24)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_25),
.A2(n_58),
.B1(n_169),
.B2(n_176),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_58),
.B1(n_176),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_25),
.A2(n_58),
.B1(n_169),
.B2(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_25),
.A2(n_58),
.B1(n_257),
.B2(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_25),
.A2(n_58),
.B1(n_346),
.B2(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_25),
.A2(n_58),
.B1(n_387),
.B2(n_570),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_25),
.A2(n_46),
.B1(n_58),
.B2(n_610),
.Y(n_609)
);

AO21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B(n_37),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_32),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_32),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_33),
.A2(n_124),
.B1(n_131),
.B2(n_134),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_34),
.Y(n_133)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_37),
.A2(n_65),
.B1(n_578),
.B2(n_579),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_39),
.Y(n_286)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_40),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_41),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_43),
.Y(n_137)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_43),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_52),
.Y(n_351)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_53),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_53),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_54),
.Y(n_173)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_58),
.B(n_321),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_554),
.B(n_618),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_394),
.B(n_549),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_324),
.C(n_363),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_270),
.B(n_299),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_73),
.B(n_270),
.C(n_551),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_181),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_74),
.B(n_182),
.C(n_243),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_122),
.C(n_167),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_75),
.A2(n_167),
.B1(n_168),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_75),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_85),
.B1(n_111),
.B2(n_120),
.Y(n_75)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_76),
.Y(n_287)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_78),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_79),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_84),
.Y(n_452)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_85),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_85),
.A2(n_120),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_SL g607 ( 
.A1(n_85),
.A2(n_120),
.B(n_608),
.Y(n_607)
);

OA21x2_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_94),
.B(n_100),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_93),
.Y(n_309)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_93),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_94),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_98),
.Y(n_372)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_105),
.B2(n_108),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_104),
.Y(n_334)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_107),
.Y(n_220)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_107),
.Y(n_413)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_111),
.Y(n_263)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_118),
.Y(n_432)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_119),
.Y(n_269)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_121),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_121),
.A2(n_264),
.B1(n_278),
.B2(n_287),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_121),
.A2(n_264),
.B1(n_278),
.B2(n_306),
.Y(n_305)
);

OAI22x1_ASAP7_75t_L g352 ( 
.A1(n_121),
.A2(n_264),
.B1(n_265),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_121),
.A2(n_264),
.B1(n_306),
.B2(n_449),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_121),
.A2(n_264),
.B1(n_371),
.B2(n_561),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_121),
.A2(n_264),
.B1(n_561),
.B2(n_583),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_122),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_138),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_123),
.B(n_138),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_146),
.B1(n_156),
.B2(n_160),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_139),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_139),
.A2(n_160),
.B1(n_186),
.B2(n_252),
.Y(n_251)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_139),
.A2(n_200),
.B(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_139),
.A2(n_194),
.B1(n_415),
.B2(n_421),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_139),
.A2(n_442),
.B1(n_498),
.B2(n_516),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_141),
.Y(n_443)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_144),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_145),
.Y(n_316)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_145),
.Y(n_486)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_147),
.A2(n_184),
.B1(n_312),
.B2(n_319),
.Y(n_311)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_150),
.Y(n_425)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_151),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_151),
.Y(n_423)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_151),
.Y(n_518)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_158),
.Y(n_319)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_159),
.Y(n_340)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_179),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_243),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_203),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_183),
.A2(n_204),
.B(n_224),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_193),
.B2(n_199),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_184),
.A2(n_312),
.B1(n_422),
.B2(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_184),
.A2(n_497),
.B1(n_505),
.B2(n_507),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_189),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_189),
.Y(n_520)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_190),
.Y(n_504)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_194),
.B(n_321),
.Y(n_514)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_195),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_224),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_214),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_205),
.A2(n_225),
.B1(n_235),
.B2(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_R g373 ( 
.A1(n_205),
.A2(n_225),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_205),
.A2(n_225),
.B1(n_401),
.B2(n_407),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_205),
.A2(n_225),
.B1(n_407),
.B2(n_455),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_205),
.A2(n_225),
.B1(n_401),
.B2(n_489),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_205),
.A2(n_225),
.B(n_375),
.Y(n_574)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_206),
.A2(n_294),
.B1(n_295),
.B2(n_298),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_206),
.A2(n_215),
.B1(n_294),
.B2(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_206),
.B(n_321),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_206),
.A2(n_294),
.B1(n_295),
.B2(n_540),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_207),
.B(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_211),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_211),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_227),
.B1(n_229),
.B2(n_232),
.Y(n_226)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_220),
.Y(n_410)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_225),
.Y(n_294)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_239),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_239),
.Y(n_464)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_241),
.Y(n_437)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_242),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_242),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_255),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_245),
.A2(n_246),
.B1(n_251),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_256),
.B(n_262),
.C(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_261),
.Y(n_388)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.C(n_276),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_271),
.B(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_276),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_288),
.C(n_293),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_293),
.Y(n_302)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_322),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_300),
.B(n_322),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_301),
.B(n_546),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_303),
.B(n_304),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.C(n_320),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_305),
.B(n_534),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_310),
.A2(n_311),
.B1(n_320),
.B2(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_319),
.Y(n_521)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_320),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_321),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_321),
.B(n_474),
.Y(n_473)
);

OAI21xp33_ASAP7_75t_SL g489 ( 
.A1(n_321),
.A2(n_473),
.B(n_490),
.Y(n_489)
);

A2O1A1O1Ixp25_ASAP7_75t_L g549 ( 
.A1(n_324),
.A2(n_363),
.B(n_550),
.C(n_552),
.D(n_553),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_362),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_325),
.B(n_362),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_343),
.B1(n_360),
.B2(n_361),
.Y(n_328)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_329),
.B(n_361),
.C(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_342),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_334),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_338),
.B(n_386),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_338),
.A2(n_386),
.B(n_391),
.Y(n_596)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_359),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_352),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_345),
.B(n_352),
.C(n_359),
.Y(n_365)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_392),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_364),
.B(n_392),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_365),
.B(n_599),
.C(n_600),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_382),
.Y(n_366)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_367),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_373),
.B(n_381),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_373),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_381),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_381),
.A2(n_592),
.B1(n_595),
.B2(n_603),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_382),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_391),
.Y(n_382)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_383),
.Y(n_391)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_544),
.B(n_548),
.Y(n_394)
);

OAI21x1_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_529),
.B(n_543),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_460),
.B(n_528),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_428),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_398),
.B(n_428),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_414),
.C(n_426),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_399),
.A2(n_400),
.B1(n_426),
.B2(n_427),
.Y(n_493)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_403),
.Y(n_406)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_414),
.B(n_493),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_416),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_446),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_429),
.B(n_447),
.C(n_454),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_439),
.B1(n_444),
.B2(n_445),
.Y(n_429)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_430),
.B(n_445),
.Y(n_538)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_439),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_453),
.B2(n_454),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

OAI21x1_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_494),
.B(n_527),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_492),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_462),
.B(n_492),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_487),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_463),
.A2(n_487),
.B1(n_488),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_463),
.Y(n_509)
);

OAI32xp33_ASAP7_75t_L g463 ( 
.A1(n_464),
.A2(n_465),
.A3(n_470),
.B1(n_473),
.B2(n_478),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_483),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx8_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_510),
.B(n_526),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_508),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_496),
.B(n_508),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_511),
.A2(n_522),
.B(n_525),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_515),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_514),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_524),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_524),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_531),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_532),
.A2(n_533),
.B1(n_536),
.B2(n_537),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_539),
.C(n_541),
.Y(n_547)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_538),
.A2(n_539),
.B1(n_541),
.B2(n_542),
.Y(n_537)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_538),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_539),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_545),
.B(n_547),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_545),
.B(n_547),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_604),
.C(n_615),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_597),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_557),
.A2(n_621),
.B(n_622),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_SL g557 ( 
.A(n_558),
.B(n_590),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_558),
.B(n_590),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_575),
.Y(n_558)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_559),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_568),
.C(n_574),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_560),
.B(n_574),
.Y(n_593)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_568),
.A2(n_569),
.B1(n_576),
.B2(n_589),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_568),
.A2(n_569),
.B1(n_593),
.B2(n_594),
.Y(n_592)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_569),
.B(n_613),
.C(n_614),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_570),
.Y(n_578)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_574),
.A2(n_582),
.B1(n_587),
.B2(n_588),
.Y(n_581)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_574),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_574),
.B(n_577),
.C(n_588),
.Y(n_611)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_576),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_577),
.B(n_581),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_579),
.Y(n_610)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_582),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx6_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_595),
.C(n_596),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_592),
.Y(n_603)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_593),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_596),
.B(n_602),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_598),
.B(n_601),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_598),
.B(n_601),
.Y(n_621)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

A2O1A1O1Ixp25_ASAP7_75t_L g619 ( 
.A1(n_605),
.A2(n_616),
.B(n_620),
.C(n_623),
.D(n_624),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_606),
.B(n_612),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_612),
.Y(n_623)
);

BUFx24_ASAP7_75t_SL g628 ( 
.A(n_606),
.Y(n_628)
);

FAx1_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_609),
.CI(n_611),
.CON(n_606),
.SN(n_606)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_607),
.B(n_609),
.C(n_611),
.Y(n_617)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);


endmodule