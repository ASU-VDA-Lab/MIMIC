module fake_jpeg_11334_n_604 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_604);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_604;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_535;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_63),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_65),
.Y(n_193)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_68),
.Y(n_181)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_83),
.Y(n_128)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_74),
.Y(n_140)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_81),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_22),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_82),
.A2(n_56),
.B1(n_32),
.B2(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_16),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_92),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_16),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_98),
.B(n_118),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_102),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_23),
.B(n_15),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_23),
.B(n_14),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_107),
.Y(n_134)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_24),
.B(n_14),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_108),
.Y(n_194)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_40),
.Y(n_112)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_20),
.Y(n_114)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_30),
.Y(n_117)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_120),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

NAND2x1_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_46),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_31),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_74),
.A2(n_45),
.B1(n_51),
.B2(n_37),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_123),
.A2(n_50),
.B1(n_2),
.B2(n_4),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_129),
.B(n_136),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_122),
.A2(n_36),
.B1(n_49),
.B2(n_40),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_130),
.A2(n_138),
.B1(n_157),
.B2(n_169),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_37),
.C(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_94),
.A2(n_49),
.B1(n_35),
.B2(n_51),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_144),
.A2(n_177),
.B1(n_34),
.B2(n_46),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_49),
.B1(n_35),
.B2(n_26),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_55),
.C(n_47),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_165),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_72),
.B(n_44),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_164),
.B(n_191),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_63),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_104),
.A2(n_35),
.B1(n_55),
.B2(n_47),
.Y(n_169)
);

INVx6_ASAP7_75t_SL g170 ( 
.A(n_65),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

BUFx12f_ASAP7_75t_SL g174 ( 
.A(n_92),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_174),
.B(n_62),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_56),
.B1(n_32),
.B2(n_25),
.Y(n_177)
);

INVx6_ASAP7_75t_SL g183 ( 
.A(n_108),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_183),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_76),
.A2(n_38),
.B1(n_26),
.B2(n_42),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_186),
.A2(n_42),
.B1(n_38),
.B2(n_34),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_89),
.B(n_29),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_116),
.A2(n_24),
.B1(n_29),
.B2(n_44),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_68),
.B1(n_67),
.B2(n_64),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_201),
.Y(n_282)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_128),
.A2(n_118),
.A3(n_106),
.B1(n_95),
.B2(n_96),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_211),
.Y(n_278)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_212),
.A2(n_235),
.B1(n_239),
.B2(n_168),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_213),
.A2(n_215),
.B1(n_238),
.B2(n_241),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_171),
.A2(n_133),
.B1(n_134),
.B2(n_150),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_217),
.Y(n_311)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_218),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_222),
.Y(n_305)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_223),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_135),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_224),
.B(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_225),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_226),
.A2(n_228),
.B1(n_243),
.B2(n_268),
.Y(n_317)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_227),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_187),
.A2(n_147),
.B1(n_180),
.B2(n_140),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_229),
.Y(n_324)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_141),
.Y(n_230)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_230),
.Y(n_309)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_152),
.B(n_14),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_124),
.B(n_131),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_234),
.B(n_246),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_158),
.A2(n_81),
.B1(n_91),
.B2(n_85),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_130),
.A2(n_97),
.B1(n_88),
.B2(n_79),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_240),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_186),
.A2(n_60),
.B1(n_59),
.B2(n_50),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_137),
.Y(n_243)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_178),
.Y(n_244)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_245),
.B(n_250),
.Y(n_297)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

AO22x2_ASAP7_75t_L g247 ( 
.A1(n_167),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_258),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_248),
.A2(n_264),
.B1(n_269),
.B2(n_193),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_13),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_249),
.B(n_259),
.Y(n_275)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_257),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_169),
.A2(n_13),
.B(n_12),
.C(n_11),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_253),
.B(n_5),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_13),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_254),
.B(n_260),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_167),
.Y(n_257)
);

AO22x2_ASAP7_75t_L g258 ( 
.A1(n_178),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_145),
.B(n_185),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_126),
.B(n_13),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_125),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_261),
.Y(n_308)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_262),
.B(n_263),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_147),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_138),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_149),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_266),
.Y(n_326)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_143),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_267),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_162),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_157),
.A2(n_146),
.B1(n_168),
.B2(n_184),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_272),
.A2(n_281),
.B1(n_293),
.B2(n_325),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_146),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_279),
.B(n_280),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_214),
.B(n_184),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_224),
.A2(n_198),
.B1(n_166),
.B2(n_176),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_299),
.C(n_302),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_206),
.B(n_198),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_285),
.B(n_287),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_206),
.B(n_166),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_189),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_288),
.B(n_296),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_212),
.A2(n_176),
.B1(n_181),
.B2(n_189),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_209),
.A2(n_148),
.B1(n_181),
.B2(n_163),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_304),
.B1(n_316),
.B2(n_228),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_148),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_258),
.B(n_5),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_209),
.A2(n_163),
.B1(n_193),
.B2(n_142),
.Y(n_316)
);

BUFx12_ASAP7_75t_L g320 ( 
.A(n_210),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_320),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_211),
.B(n_187),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_202),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_200),
.A2(n_142),
.B1(n_194),
.B2(n_8),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_234),
.C(n_232),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_328),
.B(n_336),
.C(n_337),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_291),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_329),
.B(n_342),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_332),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_200),
.B1(n_263),
.B2(n_217),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_226),
.C(n_222),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_246),
.C(n_229),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_274),
.A2(n_235),
.B1(n_247),
.B2(n_264),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.Y(n_376)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_341),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_291),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_274),
.A2(n_300),
.B1(n_299),
.B2(n_302),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_300),
.A2(n_247),
.B1(n_258),
.B2(n_244),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_278),
.A2(n_247),
.B1(n_253),
.B2(n_218),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_281),
.A2(n_243),
.B1(n_216),
.B2(n_207),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_347),
.A2(n_352),
.B1(n_311),
.B2(n_292),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_356),
.Y(n_398)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_296),
.A2(n_219),
.B1(n_255),
.B2(n_261),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_288),
.B(n_307),
.C(n_270),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_353),
.A2(n_354),
.B(n_359),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_283),
.A2(n_204),
.B(n_230),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_205),
.B(n_223),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_355),
.A2(n_365),
.B(n_311),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_291),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

AOI32xp33_ASAP7_75t_L g359 ( 
.A1(n_287),
.A2(n_242),
.A3(n_257),
.B1(n_8),
.B2(n_6),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_304),
.A2(n_7),
.B(n_8),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_360),
.A2(n_361),
.B(n_363),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_297),
.B(n_7),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_313),
.B(n_7),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_312),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_315),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_7),
.B(n_8),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_286),
.B(n_310),
.C(n_303),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_309),
.Y(n_374)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_367),
.B(n_324),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_275),
.A2(n_303),
.B1(n_308),
.B2(n_312),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_320),
.B1(n_340),
.B2(n_327),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_326),
.A2(n_284),
.B(n_308),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_276),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_284),
.B(n_319),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_370),
.A2(n_289),
.B1(n_277),
.B2(n_298),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_330),
.A2(n_271),
.B1(n_290),
.B2(n_273),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_371),
.A2(n_378),
.B1(n_382),
.B2(n_401),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_328),
.C(n_329),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_271),
.B1(n_290),
.B2(n_295),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_381),
.A2(n_347),
.B1(n_359),
.B2(n_364),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_330),
.A2(n_273),
.B1(n_315),
.B2(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_354),
.A2(n_309),
.B(n_292),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_388),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_324),
.B(n_305),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_390),
.B(n_407),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_323),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_395),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_305),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_399),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_276),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_345),
.A2(n_314),
.B1(n_318),
.B2(n_289),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_349),
.B(n_314),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_405),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_336),
.A2(n_277),
.B1(n_298),
.B2(n_318),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_404),
.A2(n_355),
.B1(n_370),
.B2(n_339),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_348),
.B(n_289),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_406),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_351),
.B(n_289),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_408),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_418),
.C(n_419),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_384),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_411),
.B(n_412),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_396),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_395),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_417),
.B(n_423),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_348),
.C(n_356),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_366),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_343),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_429),
.C(n_442),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_369),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_422),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_393),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_425),
.A2(n_443),
.B1(n_401),
.B2(n_404),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_368),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_427),
.B(n_437),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_374),
.B(n_353),
.C(n_342),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_392),
.A2(n_360),
.B1(n_337),
.B2(n_331),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_432),
.A2(n_438),
.B1(n_385),
.B2(n_394),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_390),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_433),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_390),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_434),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_380),
.A2(n_363),
.B1(n_361),
.B2(n_370),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_436),
.A2(n_385),
.B(n_375),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_357),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_401),
.A2(n_363),
.B1(n_361),
.B2(n_341),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_379),
.Y(n_439)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_399),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_412),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_344),
.C(n_338),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_376),
.A2(n_335),
.B1(n_365),
.B2(n_367),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_444),
.A2(n_457),
.B1(n_425),
.B2(n_428),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_429),
.B(n_398),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_465),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_447),
.A2(n_408),
.B1(n_426),
.B2(n_432),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_398),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_466),
.C(n_421),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_435),
.A2(n_371),
.B1(n_382),
.B2(n_376),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_450),
.A2(n_426),
.B1(n_428),
.B2(n_431),
.Y(n_491)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_454),
.Y(n_479)
);

AOI22x1_ASAP7_75t_L g455 ( 
.A1(n_416),
.A2(n_382),
.B1(n_371),
.B2(n_378),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_SL g503 ( 
.A1(n_455),
.A2(n_413),
.B(n_388),
.C(n_438),
.Y(n_503)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_414),
.Y(n_456)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_456),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_435),
.A2(n_376),
.B1(n_408),
.B2(n_381),
.Y(n_457)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_459),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_422),
.B(n_373),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_473),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_462),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_463),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_418),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_464),
.B(n_468),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_420),
.B(n_410),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_415),
.B(n_394),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_409),
.B(n_387),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_409),
.B(n_387),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_439),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_475),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_476),
.B(n_460),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_423),
.Y(n_480)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_440),
.Y(n_483)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

BUFx12_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_474),
.Y(n_485)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_486),
.A2(n_491),
.B1(n_375),
.B2(n_388),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_449),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_487),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_489),
.A2(n_503),
.B1(n_447),
.B2(n_450),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_458),
.A2(n_416),
.B(n_434),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_494),
.B(n_469),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_453),
.B(n_465),
.C(n_460),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_497),
.C(n_478),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_458),
.A2(n_433),
.B(n_427),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_453),
.B(n_413),
.C(n_411),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_459),
.Y(n_498)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_498),
.Y(n_516)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_501),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_417),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_469),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_448),
.B(n_415),
.Y(n_501)
);

AOI21x1_ASAP7_75t_SL g539 ( 
.A1(n_505),
.A2(n_507),
.B(n_518),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_510),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_471),
.Y(n_509)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_509),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_445),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_524),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_444),
.C(n_466),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_519),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_514),
.A2(n_388),
.B1(n_472),
.B2(n_467),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_502),
.A2(n_471),
.B(n_463),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_457),
.C(n_455),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_520),
.A2(n_507),
.B1(n_506),
.B2(n_522),
.Y(n_536)
);

FAx1_ASAP7_75t_SL g521 ( 
.A(n_490),
.B(n_424),
.CI(n_441),
.CON(n_521),
.SN(n_521)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_503),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_478),
.B(n_424),
.C(n_441),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_495),
.C(n_477),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_436),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_489),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_525),
.B(n_480),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_481),
.A2(n_479),
.B1(n_499),
.B2(n_496),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_526),
.A2(n_495),
.B1(n_491),
.B2(n_482),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_483),
.B(n_475),
.Y(n_527)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_529),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_530),
.B(n_531),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_503),
.C(n_493),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_533),
.B(n_542),
.Y(n_547)
);

AO21x1_ASAP7_75t_L g534 ( 
.A1(n_505),
.A2(n_500),
.B(n_503),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_534),
.A2(n_545),
.B1(n_520),
.B2(n_509),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_536),
.A2(n_521),
.B1(n_524),
.B2(n_512),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_537),
.A2(n_397),
.B1(n_484),
.B2(n_386),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_503),
.C(n_493),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_540),
.B(n_543),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_488),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_508),
.B(n_482),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_518),
.A2(n_488),
.B(n_482),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_544),
.A2(n_504),
.B1(n_527),
.B2(n_515),
.Y(n_549)
);

OA22x2_ASAP7_75t_L g546 ( 
.A1(n_504),
.A2(n_498),
.B1(n_472),
.B2(n_467),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_521),
.Y(n_553)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_519),
.C(n_525),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_552),
.C(n_540),
.Y(n_568)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_551),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_511),
.C(n_514),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_556),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_555),
.A2(n_561),
.B1(n_531),
.B2(n_533),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_539),
.A2(n_516),
.B(n_446),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_538),
.A2(n_517),
.B1(n_516),
.B2(n_446),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_557),
.A2(n_558),
.B1(n_534),
.B2(n_545),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_528),
.A2(n_388),
.B1(n_391),
.B2(n_386),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_539),
.A2(n_484),
.B(n_406),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_562),
.Y(n_567)
);

BUFx24_ASAP7_75t_SL g562 ( 
.A(n_532),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_566),
.A2(n_569),
.B1(n_573),
.B2(n_547),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_568),
.B(n_572),
.C(n_574),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_530),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_570),
.B(n_571),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_560),
.B(n_542),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_543),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_555),
.A2(n_553),
.B1(n_548),
.B2(n_556),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_541),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_541),
.C(n_546),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_SL g585 ( 
.A(n_575),
.B(n_372),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_563),
.A2(n_559),
.B(n_551),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_576),
.B(n_584),
.Y(n_592)
);

AO21x1_ASAP7_75t_L g577 ( 
.A1(n_563),
.A2(n_557),
.B(n_558),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_577),
.B(n_578),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_567),
.A2(n_546),
.B(n_389),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_579),
.B(n_582),
.Y(n_586)
);

AOI321xp33_ASAP7_75t_L g582 ( 
.A1(n_564),
.A2(n_383),
.A3(n_391),
.B1(n_379),
.B2(n_389),
.C(n_400),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_574),
.B(n_406),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_583),
.B(n_585),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_568),
.A2(n_383),
.B(n_400),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_581),
.A2(n_564),
.B(n_575),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_589),
.B(n_590),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_580),
.B(n_573),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_580),
.B(n_572),
.C(n_569),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_591),
.B(n_577),
.Y(n_596)
);

NOR2x1_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_565),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_593),
.A2(n_587),
.B(n_588),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_587),
.B(n_586),
.C(n_565),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_594),
.B(n_596),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_598),
.B(n_595),
.C(n_593),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_599),
.A2(n_597),
.B1(n_372),
.B2(n_358),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_600),
.Y(n_601)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_601),
.A2(n_397),
.B(n_334),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_602),
.B(n_350),
.C(n_320),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_603),
.B(n_320),
.Y(n_604)
);


endmodule