module fake_jpeg_16818_n_358 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_45),
.Y(n_71)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_21),
.B(n_20),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx2_ASAP7_75t_SL g116 ( 
.A(n_56),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_38),
.C(n_17),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_47),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_69),
.Y(n_78)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_28),
.Y(n_120)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_37),
.B1(n_41),
.B2(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_96),
.B1(n_106),
.B2(n_114),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_37),
.B1(n_41),
.B2(n_51),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_97),
.B1(n_102),
.B2(n_109),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_29),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_117),
.Y(n_129)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_48),
.B(n_49),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_98),
.B(n_40),
.Y(n_137)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_29),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_50),
.B(n_47),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_103),
.B(n_109),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_53),
.B1(n_52),
.B2(n_51),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_27),
.C(n_36),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_27),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_45),
.B1(n_48),
.B2(n_18),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_35),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_56),
.B(n_50),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_77),
.Y(n_111)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_24),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_115),
.B1(n_26),
.B2(n_34),
.Y(n_135)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_35),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_36),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_18),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_34),
.B1(n_33),
.B2(n_26),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_120),
.B1(n_38),
.B2(n_17),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_46),
.B(n_44),
.C(n_28),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_121),
.Y(n_175)
);

AOI22x1_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_53),
.B1(n_52),
.B2(n_51),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_136),
.B1(n_140),
.B2(n_149),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_44),
.A3(n_52),
.B1(n_53),
.B2(n_40),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_135),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_86),
.B1(n_97),
.B2(n_87),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_114),
.B(n_80),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_40),
.B1(n_39),
.B2(n_33),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_86),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_148),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_84),
.A2(n_34),
.B1(n_33),
.B2(n_26),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_86),
.A2(n_38),
.B1(n_17),
.B2(n_25),
.Y(n_150)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_88),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_156),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_123),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_154),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_109),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_116),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_164),
.B1(n_126),
.B2(n_147),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_161),
.A2(n_178),
.B(n_138),
.Y(n_201)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

BUFx24_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_107),
.B1(n_91),
.B2(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_82),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_173),
.Y(n_192)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_89),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_78),
.C(n_83),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_99),
.C(n_111),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_100),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_142),
.B1(n_131),
.B2(n_145),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_182),
.A2(n_188),
.B1(n_196),
.B2(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_153),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_156),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_143),
.B1(n_150),
.B2(n_121),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_140),
.B1(n_105),
.B2(n_97),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_197),
.A2(n_208),
.B1(n_111),
.B2(n_99),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_148),
.B1(n_134),
.B2(n_147),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_163),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_201),
.A2(n_203),
.B(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

HAxp5_ASAP7_75t_SL g203 ( 
.A(n_175),
.B(n_172),
.CON(n_203),
.SN(n_203)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_134),
.B1(n_92),
.B2(n_132),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_160),
.B1(n_162),
.B2(n_132),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_170),
.A2(n_138),
.B(n_143),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_149),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_97),
.B1(n_101),
.B2(n_112),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_201),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_194),
.C(n_199),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_180),
.B(n_189),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_219),
.B(n_236),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_171),
.B(n_173),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_220),
.B(n_221),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_127),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_222),
.B(n_224),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_180),
.A2(n_174),
.A3(n_169),
.B1(n_179),
.B2(n_165),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_209),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_146),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_159),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_228),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_192),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_25),
.C(n_32),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_237),
.Y(n_254)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_10),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_208),
.B(n_197),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_32),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_195),
.A2(n_0),
.B(n_1),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_0),
.Y(n_239)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_9),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_10),
.B(n_16),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_244),
.B1(n_251),
.B2(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_199),
.B1(n_207),
.B2(n_198),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_248),
.B(n_239),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_218),
.C(n_211),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_199),
.B1(n_193),
.B2(n_200),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_183),
.B1(n_190),
.B2(n_2),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_258),
.A2(n_4),
.B1(n_6),
.B2(n_12),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_183),
.B(n_190),
.C(n_9),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_229),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_32),
.B(n_25),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_0),
.Y(n_261)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_284),
.B1(n_287),
.B2(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_272),
.C(n_275),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_218),
.C(n_215),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_233),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_277),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_238),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_237),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_221),
.C(n_220),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_231),
.C(n_240),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_241),
.B(n_230),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_283),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_227),
.C(n_224),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_7),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_7),
.B(n_13),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_1),
.C(n_2),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_257),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_9),
.Y(n_286)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_290),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_245),
.B1(n_242),
.B2(n_243),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_302),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_246),
.B1(n_247),
.B2(n_243),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_292),
.A2(n_305),
.B1(n_280),
.B2(n_264),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_261),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_269),
.C(n_277),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_255),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_260),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_244),
.B(n_250),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_254),
.B(n_251),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_3),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_272),
.A2(n_264),
.B1(n_254),
.B2(n_262),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_279),
.B(n_260),
.CI(n_264),
.CON(n_306),
.SN(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_6),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_309),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_294),
.C(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_256),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_311),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_314),
.B1(n_319),
.B2(n_300),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_289),
.A2(n_304),
.B1(n_302),
.B2(n_295),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_2),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_317),
.B(n_318),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_291),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_2),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_303),
.B1(n_293),
.B2(n_299),
.Y(n_322)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_327),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_326),
.C(n_320),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_294),
.C(n_305),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_306),
.B1(n_292),
.B2(n_297),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_306),
.B(n_297),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_328),
.B(n_318),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_295),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_309),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_339),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_329),
.A2(n_308),
.B1(n_313),
.B2(n_315),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_336),
.A2(n_325),
.B1(n_330),
.B2(n_13),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_314),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_SL g343 ( 
.A(n_337),
.B(n_330),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_340),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_321),
.C(n_316),
.Y(n_339)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_341),
.Y(n_346)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_343),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_347),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_335),
.A2(n_12),
.B(n_13),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_339),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_344),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_351),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_342),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_352),
.B(n_346),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_338),
.B(n_350),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_333),
.C(n_14),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_14),
.Y(n_357)
);

NAND2x1_ASAP7_75t_SL g358 ( 
.A(n_357),
.B(n_14),
.Y(n_358)
);


endmodule