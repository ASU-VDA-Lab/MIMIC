module fake_netlist_6_1206_n_590 (n_52, n_16, n_1, n_46, n_18, n_21, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_42, n_8, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_80, n_41, n_86, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_590);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_42;
input n_8;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_80;
input n_41;
input n_86;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_590;

wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_125;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_300;
wire n_222;
wire n_248;
wire n_179;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_119;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_581;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_96;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_112;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_93;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_89;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_98;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_92;
wire n_513;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_548;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_175;
wire n_117;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_583;
wire n_123;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_90;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_14),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_49),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_42),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_20),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_25),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_0),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_38),
.Y(n_116)
);

BUFx8_ASAP7_75t_SL g117 ( 
.A(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_16),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_76),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_58),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_56),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_31),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_15),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_3),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_21),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_40),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_0),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_57),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_35),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_9),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_75),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_26),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_55),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_44),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_17),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_13),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_34),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_50),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_68),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_4),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_81),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_11),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_7),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_28),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_32),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_9),
.Y(n_158)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_16),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_14),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_47),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_46),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

BUFx2_ASAP7_75t_SL g165 ( 
.A(n_71),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_1),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_65),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_80),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_45),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_29),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_2),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_94),
.B(n_30),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_2),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_37),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_5),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_179)
);

AND2x4_ASAP7_75t_L g180 ( 
.A(n_102),
.B(n_61),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_102),
.B(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_108),
.A2(n_8),
.B(n_10),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_91),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

BUFx8_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_113),
.B(n_11),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

OAI21x1_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_101),
.B(n_103),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_130),
.B(n_13),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_60),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_90),
.B(n_66),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_91),
.Y(n_213)
);

CKINVDCx11_ASAP7_75t_R g214 ( 
.A(n_95),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_92),
.B(n_73),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_105),
.B(n_106),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_109),
.B(n_87),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_146),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_152),
.A2(n_74),
.B(n_82),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

CKINVDCx6p67_ASAP7_75t_R g222 ( 
.A(n_104),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_91),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_93),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_112),
.B(n_169),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_99),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_97),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_119),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_129),
.B(n_144),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_142),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_127),
.A2(n_143),
.B1(n_137),
.B2(n_134),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_118),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_124),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_128),
.Y(n_235)
);

AND2x6_ASAP7_75t_L g236 ( 
.A(n_131),
.B(n_170),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_136),
.B(n_153),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

CKINVDCx6p67_ASAP7_75t_R g239 ( 
.A(n_116),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_158),
.B(n_160),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_141),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_121),
.A2(n_138),
.B1(n_168),
.B2(n_122),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_147),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_148),
.B(n_164),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_157),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_184),
.B(n_96),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_201),
.Y(n_248)
);

BUFx6f_ASAP7_75t_SL g249 ( 
.A(n_173),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g250 ( 
.A(n_173),
.B(n_161),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_185),
.A2(n_169),
.B1(n_112),
.B2(n_123),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_184),
.B(n_98),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_172),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_100),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_173),
.B(n_167),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_228),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_185),
.B(n_111),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_115),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_175),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_172),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_201),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_240),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_174),
.B(n_140),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_193),
.A2(n_125),
.B1(n_126),
.B2(n_133),
.Y(n_280)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_228),
.B(n_149),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_171),
.B(n_151),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_204),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_192),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_192),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_200),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_178),
.A2(n_156),
.B(n_117),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_177),
.B(n_226),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_200),
.Y(n_291)
);

AND3x2_ASAP7_75t_L g292 ( 
.A(n_171),
.B(n_209),
.C(n_180),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_200),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_176),
.B(n_199),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_185),
.B(n_216),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_226),
.B(n_240),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_226),
.B(n_215),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_226),
.B(n_215),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_231),
.A2(n_216),
.B1(n_237),
.B2(n_245),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_181),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_183),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_178),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_186),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_211),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_236),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_221),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_221),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_259),
.B(n_180),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_181),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_217),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g316 ( 
.A(n_251),
.B(n_217),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_259),
.B(n_217),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_236),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_257),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_247),
.B(n_263),
.Y(n_322)
);

OAI221xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_208),
.B1(n_202),
.B2(n_246),
.C(n_209),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_263),
.B(n_232),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_264),
.B(n_231),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_259),
.B(n_212),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_236),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_257),
.B(n_236),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_300),
.B(n_242),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_269),
.B(n_236),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_239),
.B1(n_222),
.B2(n_238),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_248),
.A2(n_215),
.B1(n_212),
.B2(n_238),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_269),
.B(n_236),
.Y(n_334)
);

NAND2x1_ASAP7_75t_L g335 ( 
.A(n_250),
.B(n_220),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_252),
.B(n_230),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_254),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_269),
.B(n_212),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_250),
.B(n_188),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_250),
.B(n_188),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_252),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_278),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_273),
.A2(n_246),
.B1(n_229),
.B2(n_227),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_250),
.B(n_244),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_276),
.B(n_222),
.Y(n_346)
);

NOR2xp67_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_244),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_253),
.B(n_239),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_255),
.B(n_244),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_249),
.A2(n_227),
.B1(n_229),
.B2(n_235),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_285),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_322),
.B(n_289),
.Y(n_352)
);

NOR2x1p5_ASAP7_75t_SL g353 ( 
.A(n_311),
.B(n_271),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_310),
.A2(n_262),
.B(n_304),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_310),
.A2(n_262),
.B(n_304),
.Y(n_355)
);

BUFx8_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_324),
.A2(n_194),
.B(n_187),
.C(n_191),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_214),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_271),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_307),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_312),
.C(n_325),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_339),
.A2(n_317),
.B(n_326),
.Y(n_366)
);

BUFx4f_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

O2A1O1Ixp33_ASAP7_75t_L g368 ( 
.A1(n_305),
.A2(n_241),
.B(n_233),
.C(n_234),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_317),
.A2(n_282),
.B(n_258),
.Y(n_369)
);

NOR2x1_ASAP7_75t_R g370 ( 
.A(n_326),
.B(n_179),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_316),
.B(n_272),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_314),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_316),
.A2(n_249),
.B1(n_281),
.B2(n_289),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_305),
.A2(n_194),
.B1(n_220),
.B2(n_211),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_272),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_224),
.Y(n_376)
);

CKINVDCx8_ASAP7_75t_R g377 ( 
.A(n_330),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_268),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_306),
.A2(n_274),
.B(n_265),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_333),
.B(n_233),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_267),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_323),
.A2(n_220),
.B1(n_235),
.B2(n_243),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_338),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_277),
.B(n_267),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_243),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_268),
.B(n_260),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_332),
.B(n_234),
.Y(n_387)
);

NOR3xp33_ASAP7_75t_L g388 ( 
.A(n_344),
.B(n_224),
.C(n_241),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_328),
.A2(n_256),
.B(n_291),
.Y(n_390)
);

O2A1O1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_319),
.A2(n_266),
.B(n_279),
.C(n_253),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_343),
.B(n_270),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_331),
.A2(n_256),
.B(n_288),
.Y(n_394)
);

O2A1O1Ixp33_ASAP7_75t_L g395 ( 
.A1(n_350),
.A2(n_279),
.B(n_266),
.C(n_183),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_218),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_345),
.A2(n_191),
.B1(n_189),
.B2(n_223),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_327),
.A2(n_189),
.B(n_213),
.C(n_210),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_334),
.A2(n_256),
.B(n_288),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_213),
.B(n_197),
.C(n_205),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_315),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_308),
.B(n_219),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_313),
.A2(n_287),
.B(n_293),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_372),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_287),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_379),
.A2(n_270),
.B(n_205),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

AO21x2_ASAP7_75t_L g408 ( 
.A1(n_352),
.A2(n_206),
.B(n_197),
.Y(n_408)
);

AOI21x1_ASAP7_75t_L g409 ( 
.A1(n_354),
.A2(n_207),
.B(n_219),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_361),
.B(n_207),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_351),
.A2(n_270),
.B(n_182),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_392),
.Y(n_414)
);

OAI22x1_ASAP7_75t_L g415 ( 
.A1(n_364),
.A2(n_172),
.B1(n_182),
.B2(n_190),
.Y(n_415)
);

BUFx8_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_383),
.Y(n_417)
);

AOI21xp33_ASAP7_75t_L g418 ( 
.A1(n_371),
.A2(n_182),
.B(n_190),
.Y(n_418)
);

AOI221xp5_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_190),
.B1(n_376),
.B2(n_388),
.C(n_368),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_366),
.A2(n_355),
.B(n_359),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_190),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_396),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_385),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_358),
.B(n_367),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_374),
.A2(n_398),
.B(n_403),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_372),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_386),
.B(n_390),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_394),
.A2(n_399),
.B(n_369),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_372),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_400),
.A2(n_393),
.B(n_378),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_391),
.A2(n_380),
.B(n_353),
.C(n_395),
.Y(n_433)
);

OAI21x1_ASAP7_75t_SL g434 ( 
.A1(n_401),
.A2(n_381),
.B(n_397),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_356),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_370),
.A2(n_324),
.B(n_364),
.C(n_308),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_370),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_351),
.A2(n_269),
.B(n_339),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_SL g439 ( 
.A(n_377),
.B(n_323),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_374),
.A2(n_357),
.B(n_398),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_361),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_R g443 ( 
.A(n_383),
.B(n_214),
.Y(n_443)
);

AO32x2_ASAP7_75t_L g444 ( 
.A1(n_382),
.A2(n_373),
.A3(n_333),
.B1(n_401),
.B2(n_193),
.Y(n_444)
);

AO31x2_ASAP7_75t_L g445 ( 
.A1(n_357),
.A2(n_382),
.A3(n_398),
.B(n_366),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_357),
.A2(n_351),
.B(n_285),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_402),
.B(n_305),
.Y(n_447)
);

O2A1O1Ixp5_ASAP7_75t_L g448 ( 
.A1(n_352),
.A2(n_380),
.B(n_335),
.C(n_366),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_365),
.Y(n_449)
);

AOI21xp33_ASAP7_75t_L g450 ( 
.A1(n_364),
.A2(n_324),
.B(n_316),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_402),
.B(n_305),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_305),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_364),
.B(n_361),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_364),
.B(n_361),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_351),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_357),
.A2(n_351),
.B(n_285),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_451),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_451),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_414),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_407),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

AO21x2_ASAP7_75t_L g464 ( 
.A1(n_446),
.A2(n_458),
.B(n_426),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_450),
.B(n_446),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_450),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_449),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_424),
.B(n_452),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_413),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_442),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_426),
.B(n_420),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_439),
.A2(n_453),
.B1(n_456),
.B2(n_429),
.Y(n_472)
);

AO21x2_ASAP7_75t_L g473 ( 
.A1(n_433),
.A2(n_438),
.B(n_434),
.Y(n_473)
);

OA21x2_ASAP7_75t_L g474 ( 
.A1(n_418),
.A2(n_406),
.B(n_448),
.Y(n_474)
);

NOR2x1_ASAP7_75t_R g475 ( 
.A(n_435),
.B(n_425),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_457),
.A2(n_431),
.B1(n_427),
.B2(n_405),
.Y(n_476)
);

NAND2x1p5_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_404),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_437),
.A2(n_423),
.B1(n_416),
.B2(n_422),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_404),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_444),
.B(n_421),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_417),
.B(n_441),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_441),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_441),
.A2(n_419),
.B1(n_416),
.B2(n_415),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_430),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_419),
.A2(n_412),
.B(n_444),
.C(n_428),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_440),
.B(n_408),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

BUFx2_ASAP7_75t_SL g493 ( 
.A(n_479),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_492),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_486),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_490),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_463),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_459),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_461),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_467),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_462),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_466),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_464),
.A2(n_471),
.B(n_488),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_459),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_469),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_472),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_487),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_469),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_481),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_483),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_508),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_495),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_500),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

OR2x2_ASAP7_75t_SL g520 ( 
.A(n_510),
.B(n_491),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_482),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_494),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_497),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_499),
.A2(n_476),
.B1(n_478),
.B2(n_482),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_502),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_502),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_479),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_503),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_473),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_496),
.B(n_471),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_485),
.Y(n_532)
);

OAI221xp5_ASAP7_75t_L g533 ( 
.A1(n_509),
.A2(n_489),
.B1(n_477),
.B2(n_484),
.C(n_474),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_524),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_515),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_496),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_531),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_496),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_515),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_516),
.B(n_496),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_496),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_523),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_531),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_544),
.B(n_514),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_535),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_538),
.B(n_543),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_517),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_540),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_516),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_534),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_530),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_534),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_546),
.B(n_526),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_547),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_548),
.B(n_537),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_548),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_552),
.B(n_537),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_536),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_550),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_545),
.B(n_536),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_554),
.Y(n_563)
);

AOI321xp33_ASAP7_75t_L g564 ( 
.A1(n_555),
.A2(n_525),
.A3(n_549),
.B1(n_532),
.B2(n_533),
.C(n_505),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_560),
.A2(n_526),
.B1(n_525),
.B2(n_541),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_553),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_556),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_561),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_567),
.Y(n_569)
);

AOI322xp5_ASAP7_75t_L g570 ( 
.A1(n_564),
.A2(n_558),
.A3(n_562),
.B1(n_559),
.B2(n_563),
.C1(n_529),
.C2(n_527),
.Y(n_570)
);

OAI211xp5_ASAP7_75t_SL g571 ( 
.A1(n_568),
.A2(n_559),
.B(n_529),
.C(n_528),
.Y(n_571)
);

OAI221xp5_ASAP7_75t_L g572 ( 
.A1(n_570),
.A2(n_565),
.B1(n_560),
.B2(n_567),
.C(n_489),
.Y(n_572)
);

AOI21xp33_ASAP7_75t_L g573 ( 
.A1(n_571),
.A2(n_560),
.B(n_553),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_572),
.B(n_569),
.C(n_532),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_573),
.B(n_475),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_574),
.B(n_566),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_575),
.B(n_566),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_577),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_576),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_577),
.B(n_519),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_578),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_578),
.B(n_498),
.Y(n_582)
);

XNOR2x1_ASAP7_75t_L g583 ( 
.A(n_579),
.B(n_518),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_581),
.B(n_580),
.Y(n_584)
);

OAI22x1_ASAP7_75t_L g585 ( 
.A1(n_584),
.A2(n_580),
.B1(n_583),
.B2(n_582),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_585),
.A2(n_526),
.B1(n_518),
.B2(n_519),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_586),
.A2(n_526),
.B1(n_519),
.B2(n_518),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_587),
.Y(n_588)
);

AO21x2_ASAP7_75t_L g589 ( 
.A1(n_588),
.A2(n_498),
.B(n_513),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_589),
.A2(n_493),
.B1(n_506),
.B2(n_501),
.Y(n_590)
);


endmodule