module fake_jpeg_30081_n_50 (n_3, n_2, n_1, n_0, n_4, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx4f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.C(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_7),
.B(n_10),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_26),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_9),
.B(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_28),
.B1(n_26),
.B2(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_25),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_34),
.C(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_1),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_34),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_43),
.B(n_38),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_36),
.B1(n_37),
.B2(n_6),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_46),
.B(n_4),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

AOI221xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_0),
.B1(n_4),
.B2(n_46),
.C(n_44),
.Y(n_50)
);


endmodule