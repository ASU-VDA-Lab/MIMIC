module real_jpeg_9677_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_213;
wire n_179;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_3),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_59),
.B(n_71),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_69),
.B1(n_75),
.B2(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_135),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_36),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_36),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_26),
.B1(n_31),
.B2(n_188),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_3),
.A2(n_58),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_3),
.B(n_58),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_10),
.A2(n_69),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_10),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_76),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_69),
.B1(n_75),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_11),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_78),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_78),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_12),
.A2(n_69),
.B1(n_75),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_12),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_109),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_109),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_109),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_14),
.A2(n_36),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_16),
.A2(n_69),
.B1(n_75),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_16),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_92),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_92),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_92),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_17),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_17),
.A2(n_36),
.B1(n_37),
.B2(n_64),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_64),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_96),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_21),
.B(n_96),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_47),
.B1(n_80),
.B2(n_81),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_23),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_46),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_26),
.A2(n_31),
.B1(n_50),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_26),
.A2(n_31),
.B1(n_85),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_26),
.A2(n_31),
.B1(n_171),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_26),
.A2(n_31),
.B1(n_173),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_26),
.A2(n_31),
.B1(n_204),
.B2(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_27),
.A2(n_28),
.B1(n_117),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_27),
.A2(n_28),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_30),
.B1(n_38),
.B2(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_29),
.B(n_41),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_29),
.B(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_30),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_31),
.B(n_113),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_40),
.B1(n_42),
.B2(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_35),
.A2(n_40),
.B1(n_52),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_35),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_35),
.A2(n_40),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_35),
.A2(n_40),
.B1(n_179),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_35),
.A2(n_40),
.B1(n_202),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_35),
.A2(n_40),
.B1(n_138),
.B2(n_210),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_38),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_37),
.B1(n_57),
.B2(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_36),
.B(n_62),
.Y(n_217)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_37),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_39),
.Y(n_183)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_40),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_40),
.B(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_51),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_66),
.B1(n_67),
.B2(n_79),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_61),
.B1(n_63),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_56),
.A2(n_61),
.B1(n_95),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_56),
.A2(n_61),
.B1(n_104),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_56),
.A2(n_61),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_56),
.A2(n_61),
.B1(n_157),
.B2(n_212),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_59),
.B1(n_70),
.B2(n_71),
.Y(n_73)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_60),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_61),
.B(n_113),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_73),
.B1(n_74),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_73),
.B1(n_91),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_72),
.C(n_73),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_70),
.B(n_113),
.C(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_73),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.C(n_93),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_86),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_88),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.C(n_100),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_99),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_100),
.A2(n_101),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_105),
.C(n_110),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_162),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_144),
.B(n_161),
.Y(n_122)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_123),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_141),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_141),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_128),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_128),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_136),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_130),
.B1(n_136),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_145),
.B(n_147),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_153),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_148),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_151),
.Y(n_240)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_159),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_155),
.A2(n_156),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_158),
.B(n_159),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_160),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_242),
.C(n_243),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_236),
.B(n_241),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_222),
.B(n_235),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_206),
.B(n_221),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_196),
.B(n_205),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_185),
.B(n_195),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_174),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_180),
.B2(n_184),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_184),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_194),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.C(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_208),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.CI(n_214),
.CON(n_208),
.SN(n_208)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_219),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_224),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_232),
.C(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_231),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);


endmodule