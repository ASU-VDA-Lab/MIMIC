module fake_jpeg_7204_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx8_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_1),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_19),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_48),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_29),
.B1(n_30),
.B2(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_61),
.B1(n_43),
.B2(n_25),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_59),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_19),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_39),
.B(n_17),
.Y(n_76)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_31),
.B1(n_21),
.B2(n_24),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_28),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_29),
.B1(n_30),
.B2(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_68),
.Y(n_86)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_77),
.B1(n_81),
.B2(n_62),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_59),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_82),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_30),
.B1(n_33),
.B2(n_25),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_96),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_97),
.B1(n_71),
.B2(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_44),
.B1(n_58),
.B2(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_89),
.B1(n_93),
.B2(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_101),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_21),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_32),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_44),
.B1(n_58),
.B2(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_56),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_60),
.B1(n_57),
.B2(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_79),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_103),
.C(n_21),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_46),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_2),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_111),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_31),
.B(n_5),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_31),
.A3(n_75),
.B1(n_32),
.B2(n_16),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_100),
.B1(n_102),
.B2(n_66),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_118),
.B1(n_89),
.B2(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_119),
.Y(n_134)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_3),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_85),
.A3(n_103),
.B1(n_83),
.B2(n_96),
.C1(n_116),
.C2(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_66),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_60),
.C(n_64),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_84),
.C(n_94),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_115),
.B(n_138),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_132),
.C(n_139),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_94),
.B(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_137),
.B1(n_140),
.B2(n_113),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_95),
.C(n_103),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_103),
.B1(n_32),
.B2(n_16),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_118),
.B1(n_121),
.B2(n_107),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_31),
.B1(n_15),
.B2(n_14),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_144),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_140),
.B1(n_136),
.B2(n_6),
.Y(n_165)
);

OAI321xp33_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_108),
.A3(n_104),
.B1(n_117),
.B2(n_119),
.C(n_110),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_104),
.C(n_106),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_154),
.C(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_105),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

AO221x1_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.C(n_135),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_12),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_123),
.B(n_129),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_157),
.B(n_142),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_123),
.B(n_129),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_7),
.B(n_8),
.Y(n_177)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_143),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_153),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_154),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_176),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_143),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_10),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_172),
.B(n_158),
.C(n_165),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_163),
.CI(n_9),
.CON(n_191),
.SN(n_191)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_157),
.B(n_170),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_160),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_160),
.C(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_162),
.B1(n_163),
.B2(n_169),
.Y(n_189)
);

OAI21x1_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_182),
.B(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_174),
.C(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_191),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_7),
.B(n_9),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_195),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_179),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_191),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_10),
.B(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_10),
.Y(n_203)
);


endmodule