module fake_jpeg_11295_n_103 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_4),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_37),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_14),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_3),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_86),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_21),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_22),
.C(n_23),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_24),
.B(n_28),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_96),
.Y(n_98)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_93),
.B1(n_92),
.B2(n_83),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_90),
.B(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);


endmodule