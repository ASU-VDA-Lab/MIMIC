module fake_jpeg_27046_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_10),
.B1(n_12),
.B2(n_19),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

CKINVDCx12_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_24),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_20),
.C(n_16),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_24),
.C(n_22),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_35),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_23),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_39),
.B1(n_26),
.B2(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_15),
.B1(n_19),
.B2(n_11),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_27),
.B1(n_26),
.B2(n_11),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_52),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_34),
.C(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_3),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_62),
.C(n_65),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_34),
.C(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_55),
.C(n_47),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_4),
.B(n_5),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_4),
.B(n_5),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_74),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_54),
.B1(n_50),
.B2(n_45),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_78),
.B1(n_67),
.B2(n_59),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_42),
.C(n_34),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_65),
.C(n_57),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_63),
.B(n_6),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_78),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.C(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_70),
.C(n_76),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_57),
.B(n_64),
.C(n_7),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_77),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_88),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_70),
.C(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_82),
.B(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_71),
.C(n_8),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_97),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_71),
.B(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_91),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_101),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.Y(n_105)
);


endmodule