module fake_jpeg_1443_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_43),
.B1(n_36),
.B2(n_46),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_40),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_54),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_63),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_41),
.B1(n_47),
.B2(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_71),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_70),
.B1(n_15),
.B2(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_72),
.Y(n_79)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_49),
.B1(n_52),
.B2(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_4),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_75),
.Y(n_83)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_77),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_19),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_54),
.B(n_20),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_26),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_16),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_5),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_6),
.C(n_7),
.Y(n_95)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_77),
.B(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_95),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_6),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_10),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_22),
.B(n_32),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_27),
.B(n_31),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_7),
.B(n_8),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_103),
.B(n_85),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_13),
.B1(n_14),
.B2(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_9),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_87),
.C(n_84),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_11),
.C(n_12),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_89),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_90),
.A3(n_85),
.B1(n_12),
.B2(n_13),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.C(n_115),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_28),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_91),
.C(n_98),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_113),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_125),
.B(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_108),
.B(n_105),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_111),
.B1(n_93),
.B2(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_112),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_114),
.B(n_127),
.C(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

NAND2x1p5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_30),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_34),
.Y(n_133)
);


endmodule