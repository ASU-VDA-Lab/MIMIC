module fake_jpeg_16157_n_24 (n_3, n_2, n_1, n_0, n_4, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx6_ASAP7_75t_SL g7 ( 
.A(n_1),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_4),
.B(n_0),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g9 ( 
.A1(n_1),
.A2(n_2),
.B1(n_0),
.B2(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_15),
.B(n_6),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_10),
.C(n_9),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_14),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_19),
.C(n_2),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_SL g19 ( 
.A1(n_14),
.A2(n_9),
.B(n_6),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_7),
.B1(n_3),
.B2(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_22),
.B(n_5),
.Y(n_24)
);


endmodule