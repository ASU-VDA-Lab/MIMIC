module fake_jpeg_16018_n_91 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_23),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_8),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_17),
.B1(n_5),
.B2(n_6),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_63),
.B1(n_8),
.B2(n_11),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_29),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_60),
.B(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

AO21x1_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_62),
.B(n_64),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_28),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_68),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_48),
.B1(n_39),
.B2(n_31),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_57),
.B1(n_53),
.B2(n_63),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_57),
.B1(n_58),
.B2(n_35),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_40),
.B1(n_50),
.B2(n_64),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_42),
.B1(n_33),
.B2(n_35),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_74),
.B(n_67),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_30),
.C(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_80),
.B(n_72),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_83),
.C(n_80),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_85),
.C(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_70),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_33),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_77),
.B1(n_76),
.B2(n_65),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_67),
.B(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_89),
.B1(n_66),
.B2(n_42),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_90),
.A2(n_45),
.B(n_36),
.Y(n_91)
);


endmodule