module fake_aes_3313_n_30 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_SL g12 ( .A(n_9), .B(n_7), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_6), .B(n_11), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_16), .B(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_16), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
NAND3xp33_ASAP7_75t_L g22 ( .A(n_21), .B(n_20), .C(n_17), .Y(n_22) );
AOI221xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .B1(n_14), .B2(n_15), .C(n_13), .Y(n_23) );
OAI21xp5_ASAP7_75t_SL g24 ( .A1(n_23), .A2(n_14), .B(n_12), .Y(n_24) );
AOI221xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_1), .B1(n_2), .B2(n_3), .C(n_4), .Y(n_25) );
NOR3xp33_ASAP7_75t_L g26 ( .A(n_24), .B(n_25), .C(n_3), .Y(n_26) );
AND2x4_ASAP7_75t_L g27 ( .A(n_24), .B(n_2), .Y(n_27) );
O2A1O1Ixp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_8), .B(n_10), .C(n_5), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
AOI21xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_26), .B(n_5), .Y(n_30) );
endmodule