module real_aes_2645_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_602;
wire n_139;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g577 ( .A(n_0), .B(n_185), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_1), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g143 ( .A(n_2), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_3), .B(n_539), .Y(n_538) );
NAND2xp33_ASAP7_75t_SL g620 ( .A(n_4), .B(n_172), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_5), .B(n_152), .Y(n_176) );
INVx1_ASAP7_75t_L g613 ( .A(n_6), .Y(n_613) );
INVx1_ASAP7_75t_L g198 ( .A(n_7), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_8), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_9), .Y(n_214) );
AND2x2_ASAP7_75t_L g536 ( .A(n_10), .B(n_229), .Y(n_536) );
INVx2_ASAP7_75t_L g151 ( .A(n_11), .Y(n_151) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_12), .B(n_110), .C(n_112), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_12), .Y(n_507) );
INVx1_ASAP7_75t_L g186 ( .A(n_13), .Y(n_186) );
AOI221x1_ASAP7_75t_L g616 ( .A1(n_14), .A2(n_203), .B1(n_541), .B2(n_617), .C(n_619), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_15), .B(n_539), .Y(n_600) );
INVx1_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
INVx1_ASAP7_75t_L g183 ( .A(n_17), .Y(n_183) );
INVx1_ASAP7_75t_SL g258 ( .A(n_18), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_19), .B(n_163), .Y(n_162) );
AOI33xp33_ASAP7_75t_L g235 ( .A1(n_20), .A2(n_50), .A3(n_140), .B1(n_158), .B2(n_236), .B3(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_21), .A2(n_541), .B(n_542), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_22), .B(n_185), .Y(n_543) );
AOI221xp5_ASAP7_75t_SL g587 ( .A1(n_23), .A2(n_40), .B1(n_539), .B2(n_541), .C(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g207 ( .A(n_24), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_25), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_26), .A2(n_119), .B1(n_120), .B2(n_500), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_26), .Y(n_119) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_27), .A2(n_92), .B(n_151), .Y(n_150) );
OR2x2_ASAP7_75t_L g153 ( .A(n_27), .B(n_92), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_28), .B(n_188), .Y(n_604) );
INVxp67_ASAP7_75t_L g615 ( .A(n_29), .Y(n_615) );
AND2x2_ASAP7_75t_L g562 ( .A(n_30), .B(n_228), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_31), .B(n_196), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_32), .A2(n_541), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_33), .B(n_188), .Y(n_589) );
AND2x2_ASAP7_75t_L g146 ( .A(n_34), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g157 ( .A(n_34), .Y(n_157) );
AND2x2_ASAP7_75t_L g172 ( .A(n_34), .B(n_143), .Y(n_172) );
INVxp67_ASAP7_75t_L g112 ( .A(n_35), .Y(n_112) );
OR2x6_ASAP7_75t_L g509 ( .A(n_35), .B(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_36), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_37), .B(n_196), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_38), .A2(n_137), .B1(n_149), .B2(n_152), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_39), .B(n_169), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_41), .A2(n_82), .B1(n_155), .B2(n_541), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_42), .B(n_163), .Y(n_259) );
AOI22xp5_ASAP7_75t_SL g814 ( .A1(n_43), .A2(n_73), .B1(n_815), .B2(n_816), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_43), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_44), .B(n_185), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_45), .B(n_174), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_46), .B(n_163), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_47), .Y(n_148) );
AND2x2_ASAP7_75t_L g580 ( .A(n_48), .B(n_228), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_49), .B(n_228), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_51), .B(n_163), .Y(n_226) );
INVx1_ASAP7_75t_L g141 ( .A(n_52), .Y(n_141) );
INVx1_ASAP7_75t_L g165 ( .A(n_52), .Y(n_165) );
XOR2x2_ASAP7_75t_L g813 ( .A(n_53), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g227 ( .A(n_54), .B(n_228), .Y(n_227) );
AOI221xp5_ASAP7_75t_L g195 ( .A1(n_55), .A2(n_75), .B1(n_155), .B2(n_196), .C(n_197), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_56), .B(n_196), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_57), .B(n_539), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_58), .B(n_149), .Y(n_216) );
AOI21xp5_ASAP7_75t_SL g246 ( .A1(n_59), .A2(n_155), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g553 ( .A(n_60), .B(n_228), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_61), .B(n_188), .Y(n_578) );
INVx1_ASAP7_75t_L g179 ( .A(n_62), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_63), .B(n_185), .Y(n_551) );
AND2x2_ASAP7_75t_SL g605 ( .A(n_64), .B(n_229), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_65), .A2(n_541), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g225 ( .A(n_66), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_67), .B(n_188), .Y(n_544) );
AND2x2_ASAP7_75t_SL g569 ( .A(n_68), .B(n_174), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_69), .Y(n_822) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_70), .A2(n_155), .B(n_224), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_71), .A2(n_90), .B1(n_125), .B2(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_71), .Y(n_126) );
INVx1_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
INVx1_ASAP7_75t_L g167 ( .A(n_72), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_73), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_74), .B(n_196), .Y(n_238) );
AND2x2_ASAP7_75t_L g260 ( .A(n_76), .B(n_203), .Y(n_260) );
INVx1_ASAP7_75t_L g180 ( .A(n_77), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_78), .A2(n_155), .B(n_257), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_79), .A2(n_155), .B(n_161), .C(n_173), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_80), .B(n_539), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_81), .A2(n_85), .B1(n_196), .B2(n_539), .Y(n_567) );
INVx1_ASAP7_75t_L g114 ( .A(n_83), .Y(n_114) );
AND2x2_ASAP7_75t_SL g244 ( .A(n_84), .B(n_203), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_86), .A2(n_155), .B1(n_233), .B2(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_87), .B(n_185), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_88), .B(n_185), .Y(n_590) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_89), .A2(n_123), .B1(n_124), .B2(n_127), .Y(n_122) );
INVx1_ASAP7_75t_L g127 ( .A(n_89), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_90), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_90), .B(n_130), .C(n_471), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_91), .A2(n_541), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g248 ( .A(n_93), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_94), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_95), .B(n_188), .Y(n_550) );
AND2x2_ASAP7_75t_L g239 ( .A(n_96), .B(n_203), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_97), .A2(n_205), .B(n_206), .C(n_208), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_98), .B(n_539), .Y(n_579) );
INVxp67_ASAP7_75t_L g618 ( .A(n_99), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_100), .B(n_188), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_101), .A2(n_541), .B(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g502 ( .A(n_102), .Y(n_502) );
BUFx2_ASAP7_75t_SL g828 ( .A(n_102), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_103), .B(n_163), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_116), .B(n_829), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_107), .B(n_830), .Y(n_829) );
INVx3_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_109), .B(n_113), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_114), .B(n_115), .Y(n_510) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_513), .Y(n_116) );
AOI22xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_501), .B1(n_511), .B2(n_512), .Y(n_117) );
INVx2_ASAP7_75t_L g500 ( .A(n_120), .Y(n_500) );
XNOR2x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_128), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_125), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_SL g522 ( .A1(n_125), .A2(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_434), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_357), .Y(n_129) );
INVxp67_ASAP7_75t_L g521 ( .A(n_130), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_304), .C(n_337), .Y(n_130) );
AOI211xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_261), .B(n_270), .C(n_294), .Y(n_131) );
OAI21xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_190), .B(n_240), .Y(n_132) );
OR2x2_ASAP7_75t_L g314 ( .A(n_133), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g469 ( .A(n_133), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_134), .A2(n_360), .B1(n_364), .B2(n_366), .Y(n_359) );
AND2x2_ASAP7_75t_L g396 ( .A(n_134), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_175), .Y(n_134) );
INVx1_ASAP7_75t_L g293 ( .A(n_135), .Y(n_293) );
AND2x4_ASAP7_75t_L g310 ( .A(n_135), .B(n_291), .Y(n_310) );
INVx2_ASAP7_75t_L g332 ( .A(n_135), .Y(n_332) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_135), .Y(n_415) );
AND2x2_ASAP7_75t_L g486 ( .A(n_135), .B(n_243), .Y(n_486) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_154), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_144), .C(n_148), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g196 ( .A(n_139), .B(n_145), .Y(n_196) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
OR2x6_ASAP7_75t_L g170 ( .A(n_140), .B(n_159), .Y(n_170) );
INVxp33_ASAP7_75t_L g236 ( .A(n_140), .Y(n_236) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g160 ( .A(n_141), .B(n_143), .Y(n_160) );
AND2x4_ASAP7_75t_L g188 ( .A(n_141), .B(n_166), .Y(n_188) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g541 ( .A(n_146), .B(n_160), .Y(n_541) );
INVx2_ASAP7_75t_L g159 ( .A(n_147), .Y(n_159) );
AND2x6_ASAP7_75t_L g185 ( .A(n_147), .B(n_164), .Y(n_185) );
INVx4_ASAP7_75t_L g203 ( .A(n_149), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_149), .B(n_213), .Y(n_212) );
AOI21x1_ASAP7_75t_L g573 ( .A1(n_149), .A2(n_574), .B(n_580), .Y(n_573) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
AND2x4_ASAP7_75t_L g152 ( .A(n_151), .B(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_SL g229 ( .A(n_151), .B(n_153), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_152), .B(n_171), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_152), .A2(n_246), .B(n_250), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_152), .A2(n_538), .B(n_540), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_152), .B(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_152), .B(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_152), .B(n_618), .Y(n_617) );
NOR3xp33_ASAP7_75t_L g619 ( .A(n_152), .B(n_181), .C(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_155), .A2(n_196), .B1(n_612), .B2(n_614), .Y(n_611) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_160), .Y(n_155) );
NOR2x1p5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
INVx1_ASAP7_75t_L g237 ( .A(n_158), .Y(n_237) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_168), .B(n_171), .Y(n_161) );
INVx1_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
AND2x4_ASAP7_75t_L g539 ( .A(n_163), .B(n_172), .Y(n_539) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_166), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_170), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_SL g197 ( .A1(n_170), .A2(n_171), .B(n_198), .C(n_199), .Y(n_197) );
INVxp67_ASAP7_75t_L g205 ( .A(n_170), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_170), .A2(n_171), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_170), .A2(n_171), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_170), .A2(n_171), .B(n_258), .C(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g233 ( .A(n_171), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_171), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_171), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_171), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_171), .A2(n_577), .B(n_578), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_171), .A2(n_589), .B(n_590), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_171), .A2(n_603), .B(n_604), .Y(n_602) );
INVx5_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_173), .A2(n_231), .B(n_239), .Y(n_230) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_173), .A2(n_231), .B(n_239), .Y(n_275) );
AOI21x1_ASAP7_75t_L g565 ( .A1(n_173), .A2(n_566), .B(n_569), .Y(n_565) );
INVx2_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_174), .A2(n_195), .B(n_200), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_174), .A2(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g251 ( .A(n_175), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g280 ( .A(n_175), .Y(n_280) );
INVx3_ASAP7_75t_L g291 ( .A(n_175), .Y(n_291) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_182), .B(n_189), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_181), .B(n_207), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B1(n_186), .B2(n_187), .Y(n_182) );
INVxp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVxp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_190), .A2(n_481), .B1(n_483), .B2(n_485), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_190), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_218), .Y(n_191) );
INVx3_ASAP7_75t_L g264 ( .A(n_192), .Y(n_264) );
AND2x2_ASAP7_75t_L g272 ( .A(n_192), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_192), .Y(n_302) );
NAND2x1_ASAP7_75t_SL g496 ( .A(n_192), .B(n_263), .Y(n_496) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g269 ( .A(n_194), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_194), .B(n_275), .Y(n_287) );
AND2x2_ASAP7_75t_L g300 ( .A(n_194), .B(n_201), .Y(n_300) );
AND2x4_ASAP7_75t_L g307 ( .A(n_194), .B(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_194), .Y(n_356) );
INVxp67_ASAP7_75t_L g363 ( .A(n_194), .Y(n_363) );
INVx1_ASAP7_75t_L g368 ( .A(n_194), .Y(n_368) );
INVx1_ASAP7_75t_L g217 ( .A(n_196), .Y(n_217) );
INVx1_ASAP7_75t_L g267 ( .A(n_201), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_201), .B(n_277), .Y(n_286) );
INVx2_ASAP7_75t_L g354 ( .A(n_201), .Y(n_354) );
INVx1_ASAP7_75t_L g393 ( .A(n_201), .Y(n_393) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_211), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B1(n_209), .B2(n_210), .Y(n_202) );
INVx3_ASAP7_75t_L g210 ( .A(n_203), .Y(n_210) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_210), .A2(n_221), .B(n_227), .Y(n_220) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_210), .A2(n_221), .B(n_227), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_215), .B1(n_216), .B2(n_217), .Y(n_211) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g323 ( .A(n_218), .B(n_300), .Y(n_323) );
AND2x2_ASAP7_75t_L g391 ( .A(n_218), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g405 ( .A(n_218), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_218), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_230), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2x1_ASAP7_75t_L g268 ( .A(n_220), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g361 ( .A(n_220), .B(n_354), .Y(n_361) );
AND2x2_ASAP7_75t_L g452 ( .A(n_220), .B(n_274), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_228), .Y(n_253) );
OA21x2_ASAP7_75t_L g586 ( .A1(n_228), .A2(n_587), .B(n_591), .Y(n_586) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g263 ( .A(n_230), .Y(n_263) );
INVx2_ASAP7_75t_L g308 ( .A(n_230), .Y(n_308) );
AND2x2_ASAP7_75t_L g353 ( .A(n_230), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_232), .B(n_238), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_251), .Y(n_241) );
AND2x2_ASAP7_75t_L g395 ( .A(n_242), .B(n_396), .Y(n_395) );
OR2x6_ASAP7_75t_L g454 ( .A(n_242), .B(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx4_ASAP7_75t_L g284 ( .A(n_243), .Y(n_284) );
AND2x4_ASAP7_75t_L g292 ( .A(n_243), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g327 ( .A(n_243), .B(n_252), .Y(n_327) );
INVx2_ASAP7_75t_L g376 ( .A(n_243), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_243), .B(n_350), .Y(n_425) );
AND2x2_ASAP7_75t_L g462 ( .A(n_243), .B(n_280), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_243), .B(n_345), .Y(n_470) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g303 ( .A(n_251), .B(n_292), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_251), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_251), .B(n_330), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_251), .B(n_343), .Y(n_464) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_252), .Y(n_282) );
AND2x2_ASAP7_75t_L g290 ( .A(n_252), .B(n_291), .Y(n_290) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
INVx2_ASAP7_75t_L g316 ( .A(n_252), .Y(n_316) );
INVx1_ASAP7_75t_L g349 ( .A(n_252), .Y(n_349) );
INVx1_ASAP7_75t_L g397 ( .A(n_252), .Y(n_397) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_260), .Y(n_252) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_253), .A2(n_547), .B(n_553), .Y(n_546) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_253), .A2(n_556), .B(n_562), .Y(n_555) );
AO21x2_ASAP7_75t_L g594 ( .A1(n_253), .A2(n_556), .B(n_562), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_263), .B(n_266), .Y(n_339) );
OR2x2_ASAP7_75t_L g411 ( .A(n_263), .B(n_412), .Y(n_411) );
AND4x1_ASAP7_75t_SL g457 ( .A(n_263), .B(n_439), .C(n_458), .D(n_459), .Y(n_457) );
OR2x2_ASAP7_75t_L g481 ( .A(n_264), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g318 ( .A(n_267), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_267), .B(n_276), .Y(n_468) );
AND2x2_ASAP7_75t_L g493 ( .A(n_268), .B(n_353), .Y(n_493) );
OAI32xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_278), .A3(n_283), .B1(n_285), .B2(n_288), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g366 ( .A(n_273), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g466 ( .A(n_273), .B(n_420), .Y(n_466) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
AND2x2_ASAP7_75t_L g362 ( .A(n_274), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g448 ( .A(n_274), .Y(n_448) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_275), .B(n_277), .Y(n_482) );
INVx3_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_276), .B(n_404), .Y(n_477) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_277), .Y(n_336) );
AND2x2_ASAP7_75t_L g355 ( .A(n_277), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g489 ( .A(n_279), .Y(n_489) );
NAND2x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g329 ( .A(n_280), .Y(n_329) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_280), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_283), .B(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g321 ( .A(n_284), .B(n_289), .Y(n_321) );
AND2x4_ASAP7_75t_L g343 ( .A(n_284), .B(n_293), .Y(n_343) );
AND2x4_ASAP7_75t_SL g414 ( .A(n_284), .B(n_415), .Y(n_414) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_284), .B(n_365), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_285), .A2(n_408), .B1(n_411), .B2(n_413), .Y(n_407) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_SL g427 ( .A(n_286), .Y(n_427) );
INVx2_ASAP7_75t_L g319 ( .A(n_287), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_290), .B(n_296), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_290), .A2(n_426), .B1(n_429), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g350 ( .A(n_291), .Y(n_350) );
AND2x2_ASAP7_75t_L g373 ( .A(n_291), .B(n_332), .Y(n_373) );
INVx2_ASAP7_75t_L g296 ( .A(n_292), .Y(n_296) );
OAI21xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_297), .B(n_301), .Y(n_294) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_298), .A2(n_370), .B1(n_374), .B2(n_375), .Y(n_369) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_299), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_299), .B(n_367), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_299), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
NOR3xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_320), .C(n_324), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_309), .B1(n_314), .B2(n_317), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g334 ( .A(n_307), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g374 ( .A(n_307), .B(n_361), .Y(n_374) );
AND2x2_ASAP7_75t_L g426 ( .A(n_307), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g443 ( .A(n_307), .B(n_393), .Y(n_443) );
AND2x2_ASAP7_75t_L g498 ( .A(n_307), .B(n_392), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx4_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
AND2x2_ASAP7_75t_L g375 ( .A(n_310), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_L g380 ( .A(n_313), .Y(n_380) );
AND2x2_ASAP7_75t_L g389 ( .A(n_313), .B(n_373), .Y(n_389) );
INVx1_ASAP7_75t_L g424 ( .A(n_315), .Y(n_424) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_318), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_319), .B(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B(n_333), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_326), .B(n_365), .Y(n_474) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AOI21xp33_ASAP7_75t_SL g337 ( .A1(n_329), .A2(n_338), .B(n_340), .Y(n_337) );
AND2x2_ASAP7_75t_L g484 ( .A(n_329), .B(n_343), .Y(n_484) );
AND2x4_ASAP7_75t_L g347 ( .A(n_330), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g381 ( .A(n_330), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_330), .B(n_397), .Y(n_463) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI21xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_346), .B(n_351), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_343), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_343), .B(n_348), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_344), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g406 ( .A(n_344), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_344), .Y(n_410) );
AND2x2_ASAP7_75t_L g494 ( .A(n_344), .B(n_462), .Y(n_494) );
AND2x2_ASAP7_75t_L g497 ( .A(n_344), .B(n_414), .Y(n_497) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_349), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g476 ( .A(n_353), .Y(n_476) );
AND2x2_ASAP7_75t_L g367 ( .A(n_354), .B(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_357), .B(n_435), .Y(n_518) );
INVxp67_ASAP7_75t_L g520 ( .A(n_357), .Y(n_520) );
NAND4xp75_ASAP7_75t_L g357 ( .A(n_358), .B(n_377), .C(n_398), .D(n_416), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_369), .Y(n_358) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_361), .B(n_448), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_362), .B(n_427), .Y(n_433) );
NAND2xp5_ASAP7_75t_R g449 ( .A(n_365), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g499 ( .A(n_365), .Y(n_499) );
INVx2_ASAP7_75t_L g412 ( .A(n_367), .Y(n_412) );
BUFx3_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g455 ( .A(n_373), .Y(n_455) );
AND2x2_ASAP7_75t_L g409 ( .A(n_375), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g431 ( .A(n_376), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B(n_384), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_380), .B(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_381), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_383), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B1(n_390), .B2(n_394), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
OA21x2_ASAP7_75t_L g399 ( .A1(n_392), .A2(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g420 ( .A(n_392), .Y(n_420) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g451 ( .A(n_393), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g459 ( .A(n_393), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_394), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g429 ( .A(n_397), .B(n_430), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_405), .B(n_407), .Y(n_398) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g446 ( .A(n_403), .B(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
INVx2_ASAP7_75t_SL g450 ( .A(n_414), .Y(n_450) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_428), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B1(n_423), .B2(n_426), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g479 ( .A(n_423), .Y(n_479) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_471), .Y(n_434) );
INVxp67_ASAP7_75t_L g524 ( .A(n_435), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_444), .C(n_456), .Y(n_435) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_449), .B1(n_451), .B2(n_453), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_460), .C(n_467), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVxp67_ASAP7_75t_L g523 ( .A(n_471), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_490), .Y(n_471) );
NOR3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_480), .C(n_487), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B1(n_478), .B2(n_479), .Y(n_473) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g487 ( .A(n_481), .B(n_486), .C(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI222xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B1(n_495), .B2(n_497), .C1(n_498), .C2(n_499), .Y(n_490) );
INVx1_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
NOR2x1_ASAP7_75t_R g511 ( .A(n_502), .B(n_506), .Y(n_511) );
CKINVDCx14_ASAP7_75t_R g512 ( .A(n_503), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g820 ( .A(n_503), .B(n_821), .C(n_825), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
BUFx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x6_ASAP7_75t_SL g528 ( .A(n_507), .B(n_509), .Y(n_528) );
OR2x6_ASAP7_75t_SL g812 ( .A(n_507), .B(n_508), .Y(n_812) );
OR2x2_ASAP7_75t_L g824 ( .A(n_507), .B(n_509), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_509), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_817), .C(n_820), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_813), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_525), .B1(n_529), .B2(n_810), .Y(n_515) );
AO22x2_ASAP7_75t_L g819 ( .A1(n_516), .A2(n_526), .B1(n_529), .B2(n_811), .Y(n_819) );
AOI211x1_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .C(n_522), .Y(n_516) );
INVx4_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_740), .Y(n_530) );
NOR4xp25_ASAP7_75t_SL g531 ( .A(n_532), .B(n_633), .C(n_677), .D(n_704), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_596), .B1(n_606), .B2(n_621), .C(n_623), .Y(n_532) );
AOI32xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_563), .A3(n_570), .B1(n_581), .B2(n_592), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_534), .B(n_776), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_534), .A2(n_746), .B1(n_804), .B2(n_807), .Y(n_803) );
AND2x4_ASAP7_75t_SL g534 ( .A(n_535), .B(n_545), .Y(n_534) );
INVx5_ASAP7_75t_L g595 ( .A(n_535), .Y(n_595) );
OR2x2_ASAP7_75t_L g622 ( .A(n_535), .B(n_594), .Y(n_622) );
AND2x4_ASAP7_75t_L g624 ( .A(n_535), .B(n_555), .Y(n_624) );
INVx2_ASAP7_75t_L g639 ( .A(n_535), .Y(n_639) );
OR2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_564), .Y(n_651) );
AND2x2_ASAP7_75t_L g658 ( .A(n_535), .B(n_554), .Y(n_658) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_535), .B(n_583), .Y(n_700) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_535), .Y(n_757) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx3_ASAP7_75t_SL g652 ( .A(n_545), .Y(n_652) );
AND2x2_ASAP7_75t_L g671 ( .A(n_545), .B(n_595), .Y(n_671) );
AOI32xp33_ASAP7_75t_L g786 ( .A1(n_545), .A2(n_657), .A3(n_687), .B1(n_717), .B2(n_752), .Y(n_786) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_554), .Y(n_545) );
AND2x2_ASAP7_75t_L g626 ( .A(n_546), .B(n_564), .Y(n_626) );
OR2x2_ASAP7_75t_L g642 ( .A(n_546), .B(n_555), .Y(n_642) );
INVx1_ASAP7_75t_L g665 ( .A(n_546), .Y(n_665) );
INVx2_ASAP7_75t_L g681 ( .A(n_546), .Y(n_681) );
AND2x2_ASAP7_75t_L g718 ( .A(n_546), .B(n_583), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_546), .B(n_555), .Y(n_737) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_546), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g773 ( .A(n_555), .B(n_564), .Y(n_773) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_555), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .Y(n_556) );
OR2x2_ASAP7_75t_L g621 ( .A(n_563), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g627 ( .A(n_563), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g640 ( .A(n_563), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g802 ( .A(n_563), .B(n_671), .Y(n_802) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g731 ( .A(n_564), .B(n_681), .Y(n_731) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_565), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_570), .B(n_698), .Y(n_800) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_571), .B(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
AND2x2_ASAP7_75t_L g631 ( .A(n_572), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_572), .B(n_609), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_572), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g689 ( .A(n_572), .Y(n_689) );
OR2x2_ASAP7_75t_L g708 ( .A(n_572), .B(n_635), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_572), .Y(n_715) );
NOR2xp33_ASAP7_75t_R g767 ( .A(n_572), .B(n_598), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_572), .B(n_610), .Y(n_771) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_579), .Y(n_574) );
AOI32xp33_ASAP7_75t_L g794 ( .A1(n_581), .A2(n_630), .A3(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx2_ASAP7_75t_L g661 ( .A(n_583), .Y(n_661) );
AND2x4_ASAP7_75t_L g680 ( .A(n_583), .B(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_583), .B(n_652), .Y(n_709) );
OR2x2_ASAP7_75t_L g763 ( .A(n_583), .B(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g721 ( .A(n_584), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g779 ( .A(n_584), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_585), .B(n_598), .Y(n_745) );
AND2x2_ASAP7_75t_L g782 ( .A(n_585), .B(n_748), .Y(n_782) );
INVx2_ASAP7_75t_L g632 ( .A(n_586), .Y(n_632) );
INVx2_ASAP7_75t_L g635 ( .A(n_586), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_586), .B(n_598), .Y(n_655) );
INVx1_ASAP7_75t_L g686 ( .A(n_586), .Y(n_686) );
OR2x2_ASAP7_75t_L g712 ( .A(n_586), .B(n_598), .Y(n_712) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_586), .Y(n_764) );
BUFx3_ASAP7_75t_L g793 ( .A(n_586), .Y(n_793) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g662 ( .A(n_593), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_593), .B(n_680), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_593), .B(n_751), .Y(n_750) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_594), .B(n_665), .Y(n_664) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_594), .A2(n_661), .B(n_679), .Y(n_694) );
OAI32xp33_ASAP7_75t_L g716 ( .A1(n_595), .A2(n_717), .A3(n_719), .B1(n_721), .B2(n_723), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_595), .B(n_680), .Y(n_789) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g722 ( .A(n_597), .Y(n_722) );
NOR2x1p5_ASAP7_75t_L g792 ( .A(n_597), .B(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g608 ( .A(n_598), .B(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_SL g630 ( .A(n_598), .B(n_610), .Y(n_630) );
OR2x2_ASAP7_75t_L g634 ( .A(n_598), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g669 ( .A(n_598), .Y(n_669) );
AND2x2_ASAP7_75t_L g687 ( .A(n_598), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g698 ( .A(n_598), .B(n_610), .Y(n_698) );
OR2x2_ASAP7_75t_L g760 ( .A(n_598), .B(n_761), .Y(n_760) );
OR2x2_ASAP7_75t_L g777 ( .A(n_598), .B(n_708), .Y(n_777) );
INVx1_ASAP7_75t_L g809 ( .A(n_598), .Y(n_809) );
OR2x6_ASAP7_75t_L g598 ( .A(n_599), .B(n_605), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_607), .B(n_686), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_608), .B(n_720), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g724 ( .A1(n_608), .A2(n_725), .B1(n_730), .B2(n_732), .C1(n_735), .C2(n_738), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_608), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g752 ( .A(n_608), .B(n_631), .Y(n_752) );
AND2x2_ASAP7_75t_L g714 ( .A(n_609), .B(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g729 ( .A(n_609), .B(n_634), .Y(n_729) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_610), .B(n_635), .Y(n_667) );
AND2x4_ASAP7_75t_L g688 ( .A(n_610), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g748 ( .A(n_610), .B(n_669), .Y(n_748) );
AND2x4_ASAP7_75t_L g610 ( .A(n_611), .B(n_616), .Y(n_610) );
INVx1_ASAP7_75t_SL g628 ( .A(n_622), .Y(n_628) );
NAND2xp33_ASAP7_75t_SL g797 ( .A(n_622), .B(n_652), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B(n_627), .C(n_629), .Y(n_623) );
INVx2_ASAP7_75t_SL g674 ( .A(n_624), .Y(n_674) );
AND2x2_ASAP7_75t_L g678 ( .A(n_625), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_626), .B(n_674), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_626), .A2(n_664), .B(n_700), .C(n_701), .Y(n_699) );
AND2x2_ASAP7_75t_L g776 ( .A(n_626), .B(n_757), .Y(n_776) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x4_ASAP7_75t_L g675 ( .A(n_630), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g780 ( .A(n_630), .Y(n_780) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_643), .C(n_670), .Y(n_633) );
INVx2_ASAP7_75t_L g645 ( .A(n_634), .Y(n_645) );
OR2x2_ASAP7_75t_L g692 ( .A(n_634), .B(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_635), .Y(n_676) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_638), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g730 ( .A(n_638), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_638), .B(n_718), .Y(n_784) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g742 ( .A1(n_640), .A2(n_743), .B1(n_744), .B2(n_746), .C1(n_749), .C2(n_752), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_641), .A2(n_706), .B1(n_709), .B2(n_710), .C(n_716), .Y(n_705) );
AND2x2_ASAP7_75t_L g743 ( .A(n_641), .B(n_700), .Y(n_743) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp33_ASAP7_75t_SL g656 ( .A(n_642), .B(n_657), .Y(n_656) );
AOI221x1_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B1(n_653), .B2(n_656), .C(n_659), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g796 ( .A(n_646), .B(n_734), .Y(n_796) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g654 ( .A(n_647), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
OAI32xp33_ASAP7_75t_L g762 ( .A1(n_652), .A2(n_693), .A3(n_763), .B1(n_765), .B2(n_769), .Y(n_762) );
OAI21xp33_ASAP7_75t_SL g781 ( .A1(n_653), .A2(n_782), .B(n_783), .Y(n_781) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_666), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
OR2x2_ASAP7_75t_L g663 ( .A(n_661), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g736 ( .A(n_661), .B(n_737), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_665), .A2(n_691), .B1(n_694), .B2(n_695), .C(n_699), .Y(n_690) );
INVx1_ASAP7_75t_L g766 ( .A(n_665), .Y(n_766) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_665), .Y(n_772) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_674), .B(n_739), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_682), .B(n_690), .Y(n_677) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_681), .Y(n_751) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_687), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_684), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g703 ( .A(n_686), .Y(n_703) );
INVx1_ASAP7_75t_L g693 ( .A(n_688), .Y(n_693) );
AND2x2_ASAP7_75t_SL g702 ( .A(n_688), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_688), .B(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_688), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g707 ( .A(n_698), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_703), .Y(n_768) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_724), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g720 ( .A(n_708), .Y(n_720) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_SL g734 ( .A(n_712), .Y(n_734) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_714), .B(n_792), .Y(n_791) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_715), .Y(n_728) );
BUFx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_726), .B(n_729), .Y(n_725) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g739 ( .A(n_731), .Y(n_739) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g758 ( .A(n_737), .Y(n_758) );
NOR4xp25_ASAP7_75t_L g740 ( .A(n_741), .B(n_774), .C(n_785), .D(n_798), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_753), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_743), .A2(n_754), .B(n_759), .C(n_762), .Y(n_753) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_756), .B(n_758), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g765 ( .A1(n_756), .A2(n_766), .B(n_767), .C(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
OAI21xp33_ASAP7_75t_SL g769 ( .A1(n_770), .A2(n_772), .B(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_SL g804 ( .A(n_773), .B(n_805), .Y(n_804) );
OAI221xp5_ASAP7_75t_SL g774 ( .A1(n_775), .A2(n_777), .B1(n_778), .B2(n_779), .C(n_781), .Y(n_774) );
INVx1_ASAP7_75t_SL g778 ( .A(n_776), .Y(n_778) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND3xp33_ASAP7_75t_SL g785 ( .A(n_786), .B(n_787), .C(n_794), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
OAI21xp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_801), .B(n_803), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVxp33_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
CKINVDCx11_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_813), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
BUFx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
CKINVDCx11_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
CKINVDCx8_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
endmodule