module real_jpeg_16962_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_1),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_2),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_6),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_3),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_3),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_3),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_3),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_5),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_6),
.B(n_58),
.Y(n_57)
);

AOI31xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_109),
.A3(n_113),
.B(n_116),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_6),
.B(n_55),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_6),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_6),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_7),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_7),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_7),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_7),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_7),
.B(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_7),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_8),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_8),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_8),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_73),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_12),
.B(n_149),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_13),
.Y(n_153)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_14),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_161),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_159),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_103),
.Y(n_17)
);

NOR2xp67_ASAP7_75t_SL g160 ( 
.A(n_18),
.B(n_103),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_62),
.C(n_88),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_19),
.A2(n_20),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_48),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_31),
.Y(n_21)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_22),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_23),
.B(n_27),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_29),
.Y(n_225)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_31),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.C(n_42),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_32),
.A2(n_42),
.B1(n_43),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_32),
.Y(n_191)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

XOR2x2_ASAP7_75t_L g189 ( 
.A(n_37),
.B(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_48),
.B(n_133),
.C(n_134),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_49),
.B(n_54),
.C(n_57),
.Y(n_157)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_51),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_54),
.B(n_198),
.C(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_54),
.A2(n_61),
.B1(n_200),
.B2(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_62),
.A2(n_88),
.B1(n_89),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_62),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_72),
.C(n_76),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_63),
.B(n_72),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_67),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_68),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_68),
.A2(n_209),
.B1(n_210),
.B2(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_76),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_84),
.Y(n_76)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_77),
.A2(n_78),
.B1(n_84),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_84),
.Y(n_182)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_85),
.Y(n_212)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_101),
.C(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_131),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_121),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_156),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_148),
.B1(n_154),
.B2(n_155),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_144),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_230),
.B(n_236),
.Y(n_162)
);

OAI21x1_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_192),
.B(n_229),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_183),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.C(n_181),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_172),
.C(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_174),
.B1(n_181),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_175),
.B(n_178),
.Y(n_199)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_203),
.B(n_228),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_199),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_213),
.B(n_227),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_208),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_223),
.B(n_226),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

NOR2x1p5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_235),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);


endmodule