module real_aes_14359_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_892;
wire n_372;
wire n_528;
wire n_202;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
OA21x2_ASAP7_75t_L g151 ( .A1(n_0), .A2(n_50), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g212 ( .A(n_0), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_1), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g141 ( .A(n_2), .B(n_142), .Y(n_141) );
NAND2xp33_ASAP7_75t_L g570 ( .A(n_3), .B(n_224), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g201 ( .A1(n_4), .A2(n_97), .B1(n_181), .B2(n_202), .C(n_204), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_5), .B(n_150), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_6), .B(n_560), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_7), .B(n_248), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_8), .B(n_268), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_9), .Y(n_553) );
INVx1_ASAP7_75t_L g140 ( .A(n_10), .Y(n_140) );
BUFx3_ASAP7_75t_L g144 ( .A(n_10), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_11), .B(n_156), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g669 ( .A1(n_12), .A2(n_278), .B(n_623), .C(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_13), .A2(n_18), .B1(n_522), .B2(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_13), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_14), .Y(n_304) );
BUFx10_ASAP7_75t_L g869 ( .A(n_15), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_16), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_17), .B(n_191), .Y(n_600) );
NAND2xp33_ASAP7_75t_SL g128 ( .A(n_18), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g522 ( .A(n_18), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_19), .B(n_230), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_20), .B(n_233), .Y(n_301) );
OAI21xp33_ASAP7_75t_L g402 ( .A1(n_20), .A2(n_66), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_21), .B(n_189), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_22), .B(n_588), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_23), .A2(n_571), .B(n_662), .C(n_663), .Y(n_661) );
O2A1O1Ixp5_ASAP7_75t_L g205 ( .A1(n_24), .A2(n_206), .B(n_207), .C(n_209), .Y(n_205) );
AND2x2_ASAP7_75t_L g580 ( .A(n_25), .B(n_150), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g893 ( .A(n_26), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_27), .B(n_233), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_28), .A2(n_76), .B1(n_184), .B2(n_248), .Y(n_562) );
INVx1_ASAP7_75t_L g163 ( .A(n_29), .Y(n_163) );
INVx1_ASAP7_75t_L g546 ( .A(n_30), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_31), .B(n_185), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_32), .B(n_184), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_33), .B(n_233), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_34), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g110 ( .A(n_35), .Y(n_110) );
AND3x2_ASAP7_75t_L g891 ( .A(n_35), .B(n_112), .C(n_114), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_36), .Y(n_888) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_37), .B(n_204), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_38), .B(n_233), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_39), .B(n_206), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_40), .B(n_156), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_41), .Y(n_671) );
AND2x4_ASAP7_75t_L g162 ( .A(n_42), .B(n_163), .Y(n_162) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_43), .B(n_142), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_44), .Y(n_310) );
INVx1_ASAP7_75t_L g273 ( .A(n_45), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_46), .Y(n_179) );
AND2x2_ASAP7_75t_L g137 ( .A(n_47), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_48), .B(n_184), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_49), .A2(n_91), .B1(n_184), .B2(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g211 ( .A(n_50), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_51), .B(n_150), .Y(n_197) );
INVx1_ASAP7_75t_L g152 ( .A(n_52), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_53), .B(n_138), .Y(n_154) );
AND2x4_ASAP7_75t_L g107 ( .A(n_54), .B(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_55), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_56), .B(n_224), .Y(n_276) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_57), .B(n_78), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_58), .B(n_184), .Y(n_249) );
AND2x2_ASAP7_75t_L g612 ( .A(n_59), .B(n_234), .Y(n_612) );
INVx1_ASAP7_75t_L g108 ( .A(n_60), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_61), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_62), .B(n_588), .Y(n_587) );
NAND2x1_ASAP7_75t_L g622 ( .A(n_63), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g149 ( .A(n_64), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_65), .B(n_156), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_66), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_67), .B(n_206), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_68), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_69), .B(n_184), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_70), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_71), .B(n_175), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_72), .B(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_74), .B(n_286), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_75), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_77), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_79), .B(n_233), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_80), .B(n_204), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_81), .B(n_234), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_82), .B(n_138), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_83), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_84), .B(n_191), .Y(n_619) );
NAND2xp33_ASAP7_75t_SL g541 ( .A(n_85), .B(n_192), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_86), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_87), .B(n_138), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_88), .A2(n_126), .B1(n_863), .B2(n_864), .Y(n_125) );
INVx1_ASAP7_75t_L g863 ( .A(n_88), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_89), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_90), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
INVx1_ASAP7_75t_L g182 ( .A(n_92), .Y(n_182) );
BUFx3_ASAP7_75t_L g254 ( .A(n_92), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_93), .B(n_311), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_94), .Y(n_664) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_95), .Y(n_118) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_96), .B(n_274), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_98), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_99), .B(n_138), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_116), .B(n_892), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_102), .B(n_893), .Y(n_892) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_111), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_109), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g525 ( .A(n_109), .Y(n_525) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_110), .B(n_113), .Y(n_123) );
OR2x6_ASAP7_75t_L g867 ( .A(n_111), .B(n_868), .Y(n_867) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g122 ( .A(n_115), .Y(n_122) );
OR2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_124), .Y(n_116) );
INVxp67_ASAP7_75t_L g884 ( .A(n_117), .Y(n_884) );
NOR2x1_ASAP7_75t_SL g117 ( .A(n_118), .B(n_119), .Y(n_117) );
BUFx12f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g877 ( .A(n_121), .Y(n_877) );
NOR2x1p5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_865), .B(n_870), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_526), .Y(n_126) );
OR2x2_ASAP7_75t_L g864 ( .A(n_127), .B(n_526), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_521), .B(n_524), .Y(n_127) );
INVx2_ASAP7_75t_L g523 ( .A(n_129), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_129), .B(n_881), .Y(n_883) );
NOR2x1p5_ASAP7_75t_L g129 ( .A(n_130), .B(n_462), .Y(n_129) );
NAND4xp75_ASAP7_75t_L g130 ( .A(n_131), .B(n_364), .C(n_409), .D(n_440), .Y(n_130) );
NOR2xp67_ASAP7_75t_L g131 ( .A(n_132), .B(n_336), .Y(n_131) );
OAI321xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_164), .A3(n_236), .B1(n_257), .B2(n_293), .C(n_319), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_133), .A2(n_341), .B1(n_343), .B2(n_344), .Y(n_340) );
AND2x2_ASAP7_75t_L g457 ( .A(n_133), .B(n_258), .Y(n_457) );
AOI211xp5_ASAP7_75t_L g520 ( .A1(n_133), .A2(n_425), .B(n_453), .C(n_486), .Y(n_520) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g280 ( .A(n_134), .B(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_SL g502 ( .A(n_134), .B(n_261), .Y(n_502) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g335 ( .A(n_135), .B(n_281), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_135), .B(n_261), .Y(n_351) );
INVx1_ASAP7_75t_L g363 ( .A(n_135), .Y(n_363) );
AND2x2_ASAP7_75t_L g374 ( .A(n_135), .B(n_327), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_135), .B(n_416), .Y(n_415) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_148), .B(n_158), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B(n_145), .Y(n_136) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
INVx2_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
INVx1_ASAP7_75t_L g274 ( .A(n_139), .Y(n_274) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g203 ( .A(n_140), .Y(n_203) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
INVx3_ASAP7_75t_L g270 ( .A(n_143), .Y(n_270) );
INVx2_ASAP7_75t_L g543 ( .A(n_143), .Y(n_543) );
INVx2_ASAP7_75t_L g560 ( .A(n_143), .Y(n_560) );
INVx2_ASAP7_75t_L g588 ( .A(n_143), .Y(n_588) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx2_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
NAND3xp33_ASAP7_75t_L g561 ( .A(n_146), .B(n_406), .C(n_556), .Y(n_561) );
O2A1O1Ixp5_ASAP7_75t_L g620 ( .A1(n_146), .A2(n_174), .B(n_621), .C(n_622), .Y(n_620) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
NOR2xp67_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
AOI21xp33_ASAP7_75t_L g158 ( .A1(n_149), .A2(n_159), .B(n_160), .Y(n_158) );
INVxp33_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
INVx1_ASAP7_75t_L g216 ( .A(n_150), .Y(n_216) );
INVx1_ASAP7_75t_L g264 ( .A(n_150), .Y(n_264) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_150), .Y(n_579) );
NOR2xp67_ASAP7_75t_SL g604 ( .A(n_150), .B(n_315), .Y(n_604) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g235 ( .A(n_151), .Y(n_235) );
BUFx2_ASAP7_75t_L g244 ( .A(n_151), .Y(n_244) );
INVxp33_ASAP7_75t_L g547 ( .A(n_151), .Y(n_547) );
INVx1_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_157), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_157), .A2(n_606), .B(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR3xp33_ASAP7_75t_L g200 ( .A(n_161), .B(n_201), .C(n_205), .Y(n_200) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g196 ( .A(n_162), .Y(n_196) );
BUFx6f_ASAP7_75t_SL g255 ( .A(n_162), .Y(n_255) );
INVx1_ASAP7_75t_L g315 ( .A(n_162), .Y(n_315) );
INVx1_ASAP7_75t_L g557 ( .A(n_162), .Y(n_557) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_165), .A2(n_381), .B1(n_419), .B2(n_428), .C1(n_430), .C2(n_432), .Y(n_418) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_198), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g443 ( .A(n_167), .Y(n_443) );
AND2x4_ASAP7_75t_L g499 ( .A(n_167), .B(n_461), .Y(n_499) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g322 ( .A(n_168), .B(n_300), .Y(n_322) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx3_ASAP7_75t_L g329 ( .A(n_169), .Y(n_329) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_197), .Y(n_169) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_170), .A2(n_219), .B(n_232), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_170), .A2(n_219), .B(n_232), .Y(n_297) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_170), .A2(n_172), .B(n_197), .Y(n_318) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_170), .A2(n_593), .B(n_601), .Y(n_592) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_170), .A2(n_616), .B(n_624), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_170), .A2(n_593), .B(n_601), .Y(n_630) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_186), .B(n_195), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .B1(n_181), .B2(n_183), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g189 ( .A(n_176), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_176), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g248 ( .A(n_176), .Y(n_248) );
INVx2_ASAP7_75t_L g311 ( .A(n_176), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_180), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g313 ( .A(n_181), .Y(n_313) );
BUFx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g194 ( .A(n_182), .Y(n_194) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g224 ( .A(n_185), .Y(n_224) );
INVx1_ASAP7_75t_L g286 ( .A(n_185), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_185), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .B(n_193), .Y(n_186) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OAI221xp5_ASAP7_75t_L g309 ( .A1(n_192), .A2(n_310), .B1(n_311), .B2(n_312), .C(n_313), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_193), .A2(n_227), .B(n_229), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_193), .A2(n_247), .B(n_249), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_193), .A2(n_285), .B(n_287), .Y(n_284) );
AO21x1_ASAP7_75t_L g537 ( .A1(n_193), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_193), .A2(n_586), .B(n_587), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_193), .A2(n_598), .B(n_600), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_193), .A2(n_618), .B(n_619), .Y(n_617) );
BUFx10_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_195), .B(n_210), .Y(n_665) );
INVx2_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g231 ( .A(n_196), .Y(n_231) );
AND2x2_ASAP7_75t_L g383 ( .A(n_198), .B(n_354), .Y(n_383) );
INVx1_ASAP7_75t_L g392 ( .A(n_198), .Y(n_392) );
AND2x2_ASAP7_75t_L g444 ( .A(n_198), .B(n_424), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_198), .B(n_322), .Y(n_447) );
AND2x2_ASAP7_75t_L g483 ( .A(n_198), .B(n_298), .Y(n_483) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_217), .Y(n_198) );
AND2x2_ASAP7_75t_L g321 ( .A(n_199), .B(n_297), .Y(n_321) );
INVx2_ASAP7_75t_L g332 ( .A(n_199), .Y(n_332) );
AO21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_210), .B(n_214), .Y(n_199) );
NAND2xp33_ASAP7_75t_L g404 ( .A(n_200), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g228 ( .A(n_202), .Y(n_228) );
INVx2_ASAP7_75t_L g599 ( .A(n_202), .Y(n_599) );
INVx2_ASAP7_75t_L g623 ( .A(n_202), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_202), .B(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_203), .Y(n_204) );
INVx2_ASAP7_75t_L g230 ( .A(n_204), .Y(n_230) );
INVx1_ASAP7_75t_L g662 ( .A(n_204), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_204), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g225 ( .A(n_209), .Y(n_225) );
INVx2_ASAP7_75t_L g278 ( .A(n_209), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_210), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g667 ( .A(n_210), .Y(n_667) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
AOI21x1_ASAP7_75t_L g316 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_316) );
NOR2xp33_ASAP7_75t_R g214 ( .A(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g331 ( .A(n_217), .Y(n_331) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_L g399 ( .A(n_218), .Y(n_399) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_226), .B(n_231), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_225), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g558 ( .A(n_225), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_228), .A2(n_583), .B(n_584), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_231), .A2(n_617), .B(n_620), .Y(n_616) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_234), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AOI31xp33_ASAP7_75t_L g491 ( .A1(n_236), .A2(n_331), .A3(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g361 ( .A(n_238), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_238), .B(n_382), .Y(n_488) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g377 ( .A(n_239), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g388 ( .A(n_239), .Y(n_388) );
INVx1_ASAP7_75t_L g482 ( .A(n_239), .Y(n_482) );
AND2x2_ASAP7_75t_L g486 ( .A(n_239), .B(n_281), .Y(n_486) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g334 ( .A(n_240), .B(n_261), .Y(n_334) );
AND2x2_ASAP7_75t_L g408 ( .A(n_240), .B(n_363), .Y(n_408) );
AND2x2_ASAP7_75t_L g453 ( .A(n_240), .B(n_260), .Y(n_453) );
BUFx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g259 ( .A(n_241), .Y(n_259) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_245), .B(n_256), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_243), .A2(n_255), .B(n_545), .Y(n_548) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx3_ASAP7_75t_L g403 ( .A(n_244), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_250), .B(n_255), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .Y(n_250) );
AO21x1_ASAP7_75t_L g540 ( .A1(n_253), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_253), .A2(n_595), .B(n_596), .Y(n_594) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g268 ( .A(n_254), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_254), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
AOI211x1_ASAP7_75t_L g581 ( .A1(n_254), .A2(n_580), .B(n_582), .C(n_585), .Y(n_581) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_255), .A2(n_266), .B(n_275), .Y(n_265) );
INVx1_ASAP7_75t_L g292 ( .A(n_255), .Y(n_292) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_255), .A2(n_565), .B(n_568), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_255), .A2(n_579), .B(n_580), .Y(n_578) );
OAI21x1_ASAP7_75t_L g593 ( .A1(n_255), .A2(n_594), .B(n_597), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_280), .Y(n_257) );
AND2x2_ASAP7_75t_L g432 ( .A(n_258), .B(n_368), .Y(n_432) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g324 ( .A(n_259), .B(n_261), .Y(n_324) );
INVx2_ASAP7_75t_L g339 ( .A(n_259), .Y(n_339) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_L g379 ( .A(n_261), .Y(n_379) );
INVx1_ASAP7_75t_L g396 ( .A(n_261), .Y(n_396) );
INVx1_ASAP7_75t_L g416 ( .A(n_261), .Y(n_416) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_261), .Y(n_470) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_265), .B(n_279), .Y(n_262) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_269), .B(n_271), .Y(n_266) );
INVx1_ASAP7_75t_L g571 ( .A(n_268), .Y(n_571) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
AOI21x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_277), .B(n_278), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_278), .A2(n_289), .B(n_290), .Y(n_288) );
BUFx3_ASAP7_75t_L g344 ( .A(n_280), .Y(n_344) );
AND2x2_ASAP7_75t_L g458 ( .A(n_280), .B(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
INVx1_ASAP7_75t_L g349 ( .A(n_281), .Y(n_349) );
INVx1_ASAP7_75t_L g368 ( .A(n_281), .Y(n_368) );
AND2x2_ASAP7_75t_L g378 ( .A(n_281), .B(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_281), .Y(n_517) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B(n_291), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_298), .Y(n_293) );
INVxp67_ASAP7_75t_L g343 ( .A(n_294), .Y(n_343) );
AND2x2_ASAP7_75t_L g513 ( .A(n_294), .B(n_376), .Y(n_513) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_295), .B(n_298), .Y(n_478) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g461 ( .A(n_296), .B(n_332), .Y(n_461) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g338 ( .A(n_298), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g417 ( .A(n_298), .B(n_321), .Y(n_417) );
AND2x2_ASAP7_75t_L g434 ( .A(n_298), .B(n_330), .Y(n_434) );
AND2x2_ASAP7_75t_L g472 ( .A(n_298), .B(n_461), .Y(n_472) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_317), .Y(n_298) );
INVx1_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g355 ( .A(n_300), .Y(n_355) );
AND2x2_ASAP7_75t_L g376 ( .A(n_300), .B(n_318), .Y(n_376) );
INVx1_ASAP7_75t_L g422 ( .A(n_300), .Y(n_422) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_302), .B(n_402), .C(n_404), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_309), .C(n_314), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_307), .C(n_308), .Y(n_303) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_308), .A2(n_566), .B(n_567), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_308), .A2(n_610), .B(n_611), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g406 ( .A(n_316), .Y(n_406) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g354 ( .A(n_318), .B(n_355), .Y(n_354) );
AOI32xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .A3(n_325), .B1(n_328), .B2(n_333), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g359 ( .A(n_321), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g372 ( .A(n_321), .B(n_354), .Y(n_372) );
AND2x2_ASAP7_75t_L g375 ( .A(n_321), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g455 ( .A(n_321), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_321), .B(n_390), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_322), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI32xp33_ASAP7_75t_L g371 ( .A1(n_324), .A2(n_372), .A3(n_373), .B1(n_375), .B2(n_377), .Y(n_371) );
AND2x2_ASAP7_75t_L g411 ( .A(n_324), .B(n_368), .Y(n_411) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g480 ( .A(n_326), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g362 ( .A(n_327), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g345 ( .A(n_328), .Y(n_345) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g429 ( .A(n_329), .Y(n_429) );
INVx2_ASAP7_75t_L g439 ( .A(n_329), .Y(n_439) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_329), .Y(n_509) );
OR2x2_ASAP7_75t_L g519 ( .A(n_329), .B(n_401), .Y(n_519) );
INVx1_ASAP7_75t_L g342 ( .A(n_330), .Y(n_342) );
AND2x4_ASAP7_75t_SL g353 ( .A(n_330), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx2_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
AND2x2_ASAP7_75t_L g421 ( .A(n_332), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
AND2x2_ASAP7_75t_L g367 ( .A(n_334), .B(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_334), .Y(n_436) );
INVx1_ASAP7_75t_L g358 ( .A(n_335), .Y(n_358) );
INVx2_ASAP7_75t_L g454 ( .A(n_335), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B1(n_345), .B2(n_346), .C(n_352), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g449 ( .A(n_339), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g459 ( .A(n_339), .Y(n_459) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_344), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_347), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AND3x1_ASAP7_75t_L g428 ( .A(n_348), .B(n_408), .C(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g381 ( .A(n_350), .Y(n_381) );
AND2x2_ASAP7_75t_L g475 ( .A(n_350), .B(n_368), .Y(n_475) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g450 ( .A(n_351), .Y(n_450) );
AOI32xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .A3(n_358), .B1(n_359), .B2(n_361), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g476 ( .A1(n_353), .A2(n_477), .B1(n_479), .B2(n_483), .C1(n_484), .C2(n_487), .Y(n_476) );
AND2x2_ASAP7_75t_L g460 ( .A(n_354), .B(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
INVx3_ASAP7_75t_L g382 ( .A(n_362), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g364 ( .A(n_365), .B(n_384), .Y(n_364) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_369), .B(n_371), .C(n_380), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_367), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g512 ( .A(n_368), .B(n_453), .Y(n_512) );
INVx1_ASAP7_75t_L g493 ( .A(n_369), .Y(n_493) );
NOR2x1p5_ASAP7_75t_SL g437 ( .A(n_370), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g393 ( .A(n_372), .Y(n_393) );
INVx1_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g468 ( .A(n_374), .B(n_469), .Y(n_468) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_383), .Y(n_380) );
NOR2xp67_ASAP7_75t_SL g484 ( .A(n_381), .B(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .B1(n_393), .B2(n_394), .C(n_397), .Y(n_384) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_386), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g474 ( .A(n_390), .B(n_461), .Y(n_474) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_395), .A2(n_420), .B(n_423), .Y(n_419) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g407 ( .A(n_396), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g497 ( .A(n_396), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_407), .Y(n_397) );
AND2x2_ASAP7_75t_L g503 ( .A(n_398), .B(n_443), .Y(n_503) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx2_ASAP7_75t_L g427 ( .A(n_399), .Y(n_427) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g431 ( .A(n_401), .Y(n_431) );
OR2x2_ASAP7_75t_L g438 ( .A(n_401), .B(n_439), .Y(n_438) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_403), .A2(n_564), .B(n_572), .Y(n_563) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_406), .B(n_556), .C(n_558), .Y(n_555) );
AND4x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_418), .C(n_433), .D(n_435), .Y(n_409) );
OAI31xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .A3(n_413), .B(n_417), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_411), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g445 ( .A(n_414), .Y(n_445) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g481 ( .A(n_415), .B(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g505 ( .A(n_415), .B(n_459), .Y(n_505) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_416), .Y(n_425) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g424 ( .A(n_422), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .C(n_426), .Y(n_423) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_424), .Y(n_492) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g430 ( .A(n_427), .B(n_431), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_427), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_429), .Y(n_466) );
OAI21xp33_ASAP7_75t_L g435 ( .A1(n_432), .A2(n_436), .B(n_437), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_438), .A2(n_448), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_445), .B(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_451), .B2(n_455), .C(n_456), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_460), .Y(n_456) );
AND2x2_ASAP7_75t_L g501 ( .A(n_459), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_461), .B(n_509), .Y(n_508) );
NAND4xp75_ASAP7_75t_L g462 ( .A(n_463), .B(n_476), .C(n_489), .D(n_506), .Y(n_462) );
OA211x2_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_467), .B(n_471), .C(n_473), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
AO22x1_ASAP7_75t_L g500 ( .A1(n_474), .A2(n_501), .B1(n_503), .B2(n_504), .Y(n_500) );
INVxp67_ASAP7_75t_L g495 ( .A(n_475), .Y(n_495) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_480), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AOI221x1_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_494), .B1(n_496), .B2(n_498), .C(n_500), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g498 ( .A(n_492), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g516 ( .A(n_502), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_511), .B1(n_513), .B2(n_514), .C(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g880 ( .A(n_523), .Y(n_880) );
BUFx8_ASAP7_75t_L g528 ( .A(n_524), .Y(n_528) );
BUFx6f_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_746), .Y(n_529) );
NOR4xp25_ASAP7_75t_L g530 ( .A(n_531), .B(n_648), .C(n_692), .D(n_732), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_573), .B(n_625), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_549), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_533), .B(n_723), .Y(n_766) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g826 ( .A(n_534), .B(n_723), .Y(n_826) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_535), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_535), .B(n_641), .Y(n_837) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g635 ( .A(n_536), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g639 ( .A(n_536), .Y(n_639) );
AND2x2_ASAP7_75t_L g708 ( .A(n_536), .B(n_563), .Y(n_708) );
AND2x2_ASAP7_75t_L g736 ( .A(n_536), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g760 ( .A(n_536), .B(n_675), .Y(n_760) );
AND2x2_ASAP7_75t_L g790 ( .A(n_536), .B(n_675), .Y(n_790) );
AO31x2_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_540), .A3(n_544), .B(n_548), .Y(n_536) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_549), .B(n_736), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_549), .B(n_681), .Y(n_763) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_563), .Y(n_549) );
AND2x2_ASAP7_75t_L g638 ( .A(n_550), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g634 ( .A(n_551), .Y(n_634) );
AND2x2_ASAP7_75t_L g674 ( .A(n_551), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g682 ( .A(n_551), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g703 ( .A(n_551), .Y(n_703) );
AND2x2_ASAP7_75t_L g723 ( .A(n_551), .B(n_563), .Y(n_723) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_551), .Y(n_759) );
INVxp67_ASAP7_75t_L g789 ( .A(n_551), .Y(n_789) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_559), .B1(n_561), .B2(n_562), .Y(n_554) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g636 ( .A(n_563), .Y(n_636) );
INVx1_ASAP7_75t_L g641 ( .A(n_563), .Y(n_641) );
INVx1_ASAP7_75t_L g683 ( .A(n_563), .Y(n_683) );
AND2x2_ASAP7_75t_L g861 ( .A(n_563), .B(n_770), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_571), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_589), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g704 ( .A(n_575), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g710 ( .A(n_575), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_575), .B(n_696), .Y(n_731) );
AND2x2_ASAP7_75t_L g755 ( .A(n_575), .B(n_643), .Y(n_755) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g678 ( .A(n_576), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g832 ( .A(n_576), .B(n_776), .Y(n_832) );
AND2x2_ASAP7_75t_L g838 ( .A(n_576), .B(n_659), .Y(n_838) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g632 ( .A(n_577), .Y(n_632) );
AND2x2_ASAP7_75t_L g652 ( .A(n_577), .B(n_630), .Y(n_652) );
INVx2_ASAP7_75t_L g687 ( .A(n_577), .Y(n_687) );
INVx1_ASAP7_75t_L g719 ( .A(n_577), .Y(n_719) );
AND2x2_ASAP7_75t_L g726 ( .A(n_577), .B(n_679), .Y(n_726) );
AND2x2_ASAP7_75t_L g762 ( .A(n_577), .B(n_718), .Y(n_762) );
BUFx2_ASAP7_75t_L g801 ( .A(n_577), .Y(n_801) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_577), .Y(n_824) );
OR2x6_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_589), .A2(n_680), .B1(n_721), .B2(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_613), .Y(n_590) );
INVx4_ASAP7_75t_L g643 ( .A(n_591), .Y(n_643) );
NAND2xp33_ASAP7_75t_SL g694 ( .A(n_591), .B(n_695), .Y(n_694) );
OAI32xp33_ASAP7_75t_L g839 ( .A1(n_591), .A2(n_724), .A3(n_840), .B1(n_841), .B2(n_843), .Y(n_839) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_602), .Y(n_591) );
INVx2_ASAP7_75t_L g691 ( .A(n_592), .Y(n_691) );
AND2x4_ASAP7_75t_L g631 ( .A(n_602), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g651 ( .A(n_602), .Y(n_651) );
INVx2_ASAP7_75t_L g679 ( .A(n_602), .Y(n_679) );
AND2x2_ASAP7_75t_L g705 ( .A(n_602), .B(n_691), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_602), .B(n_614), .Y(n_711) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_608), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_604), .A2(n_609), .B(n_612), .Y(n_608) );
AND2x2_ASAP7_75t_L g793 ( .A(n_613), .B(n_726), .Y(n_793) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_613), .Y(n_842) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_614), .Y(n_655) );
AND2x2_ASAP7_75t_L g696 ( .A(n_614), .B(n_691), .Y(n_696) );
AND2x2_ASAP7_75t_L g775 ( .A(n_614), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g647 ( .A(n_615), .Y(n_647) );
INVx1_ASAP7_75t_L g690 ( .A(n_615), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_633), .B1(n_637), .B2(n_642), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_628), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g821 ( .A(n_628), .Y(n_821) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g728 ( .A(n_629), .B(n_646), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g847 ( .A1(n_629), .A2(n_734), .B1(n_814), .B2(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g786 ( .A(n_630), .B(n_679), .Y(n_786) );
AND2x2_ASAP7_75t_L g749 ( .A(n_631), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g771 ( .A(n_631), .B(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_631), .Y(n_830) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_632), .Y(n_817) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_634), .Y(n_713) );
AND2x2_ASAP7_75t_L g768 ( .A(n_634), .B(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g778 ( .A(n_634), .B(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g818 ( .A(n_634), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_634), .B(n_819), .Y(n_834) );
AND2x2_ASAP7_75t_L g673 ( .A(n_635), .B(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g797 ( .A(n_635), .Y(n_797) );
AOI33xp33_ASAP7_75t_L g831 ( .A1(n_635), .A2(n_643), .A3(n_714), .B1(n_832), .B2(n_833), .B3(n_838), .Y(n_831) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_637), .B(n_657), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_637), .A2(n_694), .B1(n_697), .B2(n_704), .Y(n_693) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
AND2x2_ASAP7_75t_L g792 ( .A(n_638), .B(n_769), .Y(n_792) );
AND2x4_ASAP7_75t_L g860 ( .A(n_638), .B(n_861), .Y(n_860) );
AND2x2_ASAP7_75t_L g722 ( .A(n_639), .B(n_659), .Y(n_722) );
INVx1_ASAP7_75t_L g819 ( .A(n_639), .Y(n_819) );
BUFx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_641), .Y(n_700) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_642), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g815 ( .A(n_642), .Y(n_815) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
OAI21xp33_ASAP7_75t_L g858 ( .A1(n_643), .A2(n_822), .B(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g677 ( .A(n_645), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g740 ( .A(n_645), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_645), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g718 ( .A(n_647), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_653), .B(n_656), .C(n_672), .Y(n_648) );
NAND2x1_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_650), .A2(n_856), .B1(n_858), .B2(n_862), .Y(n_855) );
INVx4_ASAP7_75t_R g650 ( .A(n_651), .Y(n_650) );
OAI32xp33_ASAP7_75t_L g820 ( .A1(n_651), .A2(n_821), .A3(n_822), .B1(n_823), .B2(n_825), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_651), .B(n_836), .Y(n_835) );
AND2x2_ASAP7_75t_L g654 ( .A(n_652), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g822 ( .A(n_657), .B(n_797), .Y(n_822) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_659), .Y(n_681) );
BUFx2_ASAP7_75t_L g715 ( .A(n_659), .Y(n_715) );
INVx1_ASAP7_75t_L g737 ( .A(n_659), .Y(n_737) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_660), .B(n_668), .Y(n_659) );
NAND2x1p5_ASAP7_75t_L g675 ( .A(n_660), .B(n_668), .Y(n_675) );
OA21x2_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_665), .B(n_666), .Y(n_660) );
OR2x2_ASAP7_75t_L g668 ( .A(n_665), .B(n_669), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B1(n_680), .B2(n_684), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g764 ( .A1(n_673), .A2(n_765), .B1(n_771), .B2(n_773), .C1(n_778), .C2(n_780), .Y(n_764) );
AND2x2_ASAP7_75t_L g707 ( .A(n_674), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g702 ( .A(n_675), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g770 ( .A(n_675), .Y(n_770) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g756 ( .A1(n_677), .A2(n_757), .B1(n_761), .B2(n_763), .Y(n_756) );
INVx2_ASAP7_75t_L g777 ( .A(n_678), .Y(n_777) );
AND2x4_ASAP7_75t_SL g686 ( .A(n_679), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
AND2x4_ASAP7_75t_SL g729 ( .A(n_682), .B(n_722), .Y(n_729) );
INVx1_ASAP7_75t_L g814 ( .A(n_682), .Y(n_814) );
AND2x2_ASAP7_75t_L g769 ( .A(n_683), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g741 ( .A(n_686), .Y(n_741) );
INVx1_ASAP7_75t_L g781 ( .A(n_686), .Y(n_781) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_SL g750 ( .A(n_689), .Y(n_750) );
INVx1_ASAP7_75t_L g806 ( .A(n_689), .Y(n_806) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
BUFx2_ASAP7_75t_L g836 ( .A(n_690), .Y(n_836) );
INVx1_ASAP7_75t_L g776 ( .A(n_691), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_706), .C(n_720), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_696), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
OR2x2_ASAP7_75t_L g796 ( .A(n_701), .B(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g809 ( .A(n_702), .B(n_708), .Y(n_809) );
INVx1_ASAP7_75t_L g735 ( .A(n_703), .Y(n_735) );
AND2x2_ASAP7_75t_L g716 ( .A(n_705), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_705), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g807 ( .A(n_705), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B1(n_712), .B2(n_716), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g745 ( .A(n_711), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_711), .A2(n_834), .B1(n_835), .B2(n_837), .Y(n_833) );
AND2x4_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_718), .Y(n_772) );
OR2x2_ASAP7_75t_L g857 ( .A(n_718), .B(n_719), .Y(n_857) );
AOI32xp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_724), .A3(n_727), .B1(n_729), .B2(n_730), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx2_ASAP7_75t_L g752 ( .A(n_723), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_723), .B(n_736), .Y(n_840) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND3xp33_ASAP7_75t_SL g851 ( .A(n_727), .B(n_807), .C(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g804 ( .A(n_729), .Y(n_804) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_738), .B(n_742), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_740), .A2(n_813), .B1(n_815), .B2(n_816), .Y(n_812) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_810), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_764), .C(n_782), .D(n_794), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .B1(n_753), .B2(n_755), .C(n_756), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g854 ( .A(n_752), .B(n_760), .Y(n_854) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
OR2x2_ASAP7_75t_L g843 ( .A(n_758), .B(n_797), .Y(n_843) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g779 ( .A(n_760), .Y(n_779) );
OR2x2_ASAP7_75t_L g813 ( .A(n_760), .B(n_814), .Y(n_813) );
OR2x2_ASAP7_75t_L g850 ( .A(n_760), .B(n_824), .Y(n_850) );
INVx1_ASAP7_75t_L g783 ( .A(n_761), .Y(n_783) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_763), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g862 ( .A(n_768), .B(n_819), .Y(n_862) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g848 ( .A(n_775), .Y(n_848) );
OAI32xp33_ASAP7_75t_L g803 ( .A1(n_780), .A2(n_804), .A3(n_805), .B1(n_807), .B2(n_808), .Y(n_803) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
O2A1O1Ixp33_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B(n_787), .C(n_791), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g802 ( .A(n_786), .Y(n_802) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
INVx1_ASAP7_75t_L g852 ( .A(n_793), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_798), .B(n_803), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NAND4xp25_ASAP7_75t_L g810 ( .A(n_811), .B(n_827), .C(n_844), .D(n_855), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_820), .Y(n_811) );
NAND3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .C(n_819), .Y(n_816) );
AOI322xp5_ASAP7_75t_L g844 ( .A1(n_821), .A2(n_845), .A3(n_846), .B1(n_847), .B2(n_849), .C1(n_851), .C2(n_853), .Y(n_844) );
OAI21xp33_ASAP7_75t_L g828 ( .A1(n_822), .A2(n_829), .B(n_831), .Y(n_828) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_824), .Y(n_846) );
INVx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_SL g827 ( .A(n_828), .B(n_839), .Y(n_827) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_SL g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx6_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx3_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_869), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_869), .B(n_891), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_885), .B(n_887), .Y(n_870) );
OAI21xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_878), .B(n_884), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx2_ASAP7_75t_SL g874 ( .A(n_875), .Y(n_874) );
BUFx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
BUFx3_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B(n_883), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_886), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
endmodule