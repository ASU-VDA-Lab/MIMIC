module fake_jpeg_12808_n_148 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NAND2x1_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_57),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_29),
.A3(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_42),
.B(n_39),
.C(n_38),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_23),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_60),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_69),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_66),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_37),
.B1(n_30),
.B2(n_18),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_51),
.B1(n_55),
.B2(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_24),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_30),
.B(n_22),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_74),
.B(n_1),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_22),
.B1(n_19),
.B2(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_10),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_7),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_12),
.B(n_5),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_56),
.B1(n_59),
.B2(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_85),
.B1(n_87),
.B2(n_68),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_55),
.C(n_45),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_94),
.C(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_48),
.B1(n_39),
.B2(n_3),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_66),
.B1(n_62),
.B2(n_61),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_78),
.B(n_68),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_1),
.C(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NAND2x1p5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_73),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_102),
.C(n_108),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_84),
.C(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_104),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_85),
.B1(n_93),
.B2(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_107),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_67),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_83),
.C(n_101),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_106),
.B(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_86),
.B1(n_100),
.B2(n_107),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.C(n_98),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_91),
.C(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_99),
.C(n_98),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_110),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

XOR2x2_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_115),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_111),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_94),
.B(n_125),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_133),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_137),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_127),
.B1(n_67),
.B2(n_92),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_132),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_143),
.C(n_135),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_5),
.A3(n_6),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_2),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_86),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.C(n_141),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_140),
.Y(n_147)
);


endmodule