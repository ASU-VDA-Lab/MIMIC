module fake_ariane_1004_n_2405 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_2405);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2405;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_1196;
wire n_462;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_2370;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2203;
wire n_2133;
wire n_2076;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2394;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_2395;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2324;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_1251;
wire n_412;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_37),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_6),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_173),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_130),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_197),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_168),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_144),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_24),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_5),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_3),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_124),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_156),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_3),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_201),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_94),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_202),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_101),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_147),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_63),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_171),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_31),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_233),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_71),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_22),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_71),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_125),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_181),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_186),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_8),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_142),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_198),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_31),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_29),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_143),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_217),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_182),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_216),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_167),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_228),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_47),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_47),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_19),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_161),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_28),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_52),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_120),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_110),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_85),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_94),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_121),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_61),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_209),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_44),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_21),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_85),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_175),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_24),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_70),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_191),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_60),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_5),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_154),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_150),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_109),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_123),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_0),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_63),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_15),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_126),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_37),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_164),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_70),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_100),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_118),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_1),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_162),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_215),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_65),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_136),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_97),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_23),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_157),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_174),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_148),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_188),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_36),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_60),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_46),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_72),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_10),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_214),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_138),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_232),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_58),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_221),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_48),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_13),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_86),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_133),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_140),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_18),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_158),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_106),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_42),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_240),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_61),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_34),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_14),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_236),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_93),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_30),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_141),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_199),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_50),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_96),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_235),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_205),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_75),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_72),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_80),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_163),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_16),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_208),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_239),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_93),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_177),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_33),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_58),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_76),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_113),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_213),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_99),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_25),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_92),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_45),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_46),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_103),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_127),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_159),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_39),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_137),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_49),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_179),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_7),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_51),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_234),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_51),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_36),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_49),
.Y(n_397)
);

BUFx8_ASAP7_75t_SL g398 ( 
.A(n_29),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_87),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_67),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_32),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_59),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_165),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_206),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_95),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_33),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_62),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_116),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_135),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_77),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_77),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_145),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_241),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_176),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_218),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_102),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_117),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_102),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_100),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_129),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_170),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_223),
.Y(n_422)
);

INVx4_ASAP7_75t_R g423 ( 
.A(n_52),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_30),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_66),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_86),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_88),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_64),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_43),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_1),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_9),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_53),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_178),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_196),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_128),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_4),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_106),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_212),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_34),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_43),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_14),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_0),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_119),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_180),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_237),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_66),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_55),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_22),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_203),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_78),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_183),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_229),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_101),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_146),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_195),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_55),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_230),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_166),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_231),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_75),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_87),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_225),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_131),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_38),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_222),
.Y(n_465)
);

BUFx2_ASAP7_75t_SL g466 ( 
.A(n_112),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_6),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_108),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_132),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_103),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_185),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_114),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_105),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_263),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_263),
.B(n_2),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_383),
.B(n_2),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_263),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_261),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_263),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_263),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_398),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_263),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_263),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_464),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_366),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_390),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_331),
.Y(n_487)
);

INVxp33_ASAP7_75t_SL g488 ( 
.A(n_269),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_333),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_263),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_306),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_383),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_431),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_439),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_306),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_365),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_286),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_242),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_374),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_306),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_306),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_306),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_306),
.Y(n_503)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_383),
.B(n_4),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_414),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_306),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_R g507 ( 
.A(n_298),
.B(n_304),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_286),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_305),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_306),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_7),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_302),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_290),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_253),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_290),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_308),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_268),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_290),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_313),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_290),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_290),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_377),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_377),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_302),
.B(n_368),
.Y(n_524)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_250),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_309),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_314),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_316),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_318),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_342),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_359),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_377),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_329),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_377),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_377),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_242),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_437),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_437),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_337),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_344),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_323),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_323),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_399),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_345),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_243),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_368),
.B(n_8),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_326),
.B(n_9),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_326),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_328),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_328),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_352),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_472),
.B(n_10),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_354),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_355),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_356),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_338),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_243),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_411),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_338),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_382),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_258),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_362),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_382),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_363),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_416),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_370),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_373),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_416),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_376),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_448),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_442),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_381),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_313),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_442),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_453),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_453),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_472),
.B(n_11),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_380),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_388),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_393),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_294),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_294),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_413),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_386),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_386),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_460),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_471),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_381),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_395),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_413),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_471),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_256),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_252),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_251),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_251),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_396),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_259),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_277),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_251),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_397),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_288),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_496),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_522),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_514),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_466),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_519),
.B(n_339),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_499),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_505),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_480),
.A2(n_283),
.B(n_255),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_522),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_522),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_485),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_519),
.B(n_509),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_522),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_487),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_492),
.B(n_262),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_480),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_474),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_586),
.B(n_262),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_586),
.B(n_407),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_474),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_477),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_486),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_477),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_517),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_479),
.Y(n_629)
);

OA21x2_ASAP7_75t_L g630 ( 
.A1(n_475),
.A2(n_296),
.B(n_292),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_530),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_479),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_497),
.B(n_407),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_482),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_549),
.B(n_265),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_478),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_489),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_482),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_531),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_483),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_493),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_483),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_516),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_507),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_513),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_591),
.B(n_456),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_SL g648 ( 
.A(n_593),
.B(n_456),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_490),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_498),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_481),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_491),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_497),
.B(n_265),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_491),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_495),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_575),
.B(n_300),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_495),
.Y(n_657)
);

CKINVDCx8_ASAP7_75t_R g658 ( 
.A(n_484),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_576),
.B(n_319),
.Y(n_659)
);

CKINVDCx8_ASAP7_75t_R g660 ( 
.A(n_526),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_576),
.B(n_325),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_500),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_527),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_513),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_591),
.B(n_327),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_500),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_R g667 ( 
.A(n_528),
.B(n_258),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_529),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_515),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_533),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_L g671 ( 
.A(n_542),
.B(n_405),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_543),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_547),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_501),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_554),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_SL g676 ( 
.A1(n_546),
.A2(n_270),
.B1(n_274),
.B2(n_266),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_501),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_591),
.B(n_330),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_561),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_502),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_556),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_502),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_591),
.B(n_343),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_596),
.B(n_353),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_557),
.B(n_341),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_503),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_573),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_R g688 ( 
.A(n_558),
.B(n_266),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_503),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_506),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_565),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_506),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_510),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_596),
.B(n_360),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_584),
.B(n_341),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_510),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_515),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_589),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_518),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_518),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_567),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_569),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_570),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_632),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_693),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_632),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_632),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_653),
.B(n_537),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_693),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_605),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_623),
.B(n_647),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

AND2x2_ASAP7_75t_SL g713 ( 
.A(n_635),
.B(n_511),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_640),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_640),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_629),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_635),
.A2(n_488),
.B1(n_494),
.B2(n_550),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_640),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_609),
.A2(n_550),
.B1(n_349),
.B2(n_555),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_642),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_685),
.B(n_572),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_642),
.Y(n_722)
);

INVx8_ASAP7_75t_L g723 ( 
.A(n_644),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_619),
.B(n_581),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_622),
.B(n_582),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_642),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_620),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_629),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_693),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_650),
.B(n_583),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_653),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_663),
.B(n_592),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_633),
.B(n_508),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_623),
.B(n_599),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_620),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_649),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_607),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_621),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_676),
.B(n_524),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_649),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_615),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_629),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_649),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_620),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_655),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_660),
.A2(n_580),
.B1(n_274),
.B2(n_278),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_655),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_655),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_623),
.B(n_524),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_645),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_657),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_623),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_657),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_621),
.B(n_603),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_647),
.B(n_508),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_633),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_645),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_645),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_645),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_608),
.B(n_604),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_624),
.B(n_584),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_647),
.B(n_595),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_657),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_608),
.B(n_248),
.Y(n_764)
);

INVx4_ASAP7_75t_SL g765 ( 
.A(n_620),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_680),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_647),
.B(n_595),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_624),
.B(n_585),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_630),
.A2(n_525),
.B1(n_560),
.B2(n_548),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_616),
.B(n_564),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_662),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_684),
.B(n_600),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_668),
.B(n_244),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_625),
.B(n_627),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_620),
.Y(n_775)
);

NOR3xp33_ASAP7_75t_L g776 ( 
.A(n_676),
.B(n_461),
.C(n_278),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_658),
.B(n_597),
.Y(n_777)
);

INVx4_ASAP7_75t_SL g778 ( 
.A(n_620),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_656),
.B(n_512),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_625),
.B(n_585),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_671),
.B(n_587),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_680),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_651),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_646),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_680),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_662),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_670),
.B(n_244),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_662),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_627),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_615),
.B(n_604),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_680),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_630),
.A2(n_504),
.B1(n_476),
.B2(n_297),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_634),
.B(n_587),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_606),
.Y(n_795)
);

NOR2x1p5_ASAP7_75t_L g796 ( 
.A(n_672),
.B(n_270),
.Y(n_796)
);

AO22x2_ASAP7_75t_L g797 ( 
.A1(n_684),
.A2(n_590),
.B1(n_594),
.B2(n_588),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_646),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_690),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_673),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_690),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_681),
.B(n_246),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_695),
.B(n_600),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_606),
.Y(n_804)
);

AND2x6_ASAP7_75t_L g805 ( 
.A(n_634),
.B(n_248),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_613),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_695),
.B(n_601),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_690),
.Y(n_808)
);

INVx1_ASAP7_75t_SL g809 ( 
.A(n_628),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_638),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_694),
.B(n_601),
.Y(n_811)
);

AND2x6_ASAP7_75t_L g812 ( 
.A(n_638),
.B(n_248),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_636),
.B(n_282),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_697),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_643),
.B(n_588),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_652),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_613),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_659),
.B(n_544),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_697),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_667),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_630),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_691),
.B(n_246),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_614),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_630),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_610),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_614),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_617),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_646),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_SL g829 ( 
.A(n_658),
.B(n_598),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_675),
.B(n_590),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_697),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_652),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_700),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_617),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_659),
.B(n_544),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_699),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_701),
.B(n_247),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_L g838 ( 
.A(n_654),
.B(n_245),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_654),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_702),
.B(n_247),
.Y(n_840)
);

INVx5_ASAP7_75t_L g841 ( 
.A(n_646),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_646),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_694),
.B(n_545),
.Y(n_843)
);

OAI21xp33_ASAP7_75t_L g844 ( 
.A1(n_666),
.A2(n_301),
.B(n_299),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_661),
.B(n_545),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_666),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_674),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_674),
.B(n_245),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_677),
.B(n_594),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_703),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_677),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_682),
.B(n_520),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_688),
.A2(n_282),
.B1(n_291),
.B2(n_287),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_682),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_686),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_686),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_665),
.B(n_551),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_689),
.B(n_602),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_689),
.B(n_369),
.Y(n_859)
);

OAI22xp33_ASAP7_75t_L g860 ( 
.A1(n_660),
.A2(n_291),
.B1(n_295),
.B2(n_287),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_665),
.B(n_678),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_611),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_646),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_692),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_692),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_696),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_795),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_861),
.B(n_696),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_704),
.Y(n_869)
);

AND2x6_ASAP7_75t_SL g870 ( 
.A(n_739),
.B(n_315),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_713),
.A2(n_410),
.B1(n_427),
.B2(n_295),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_713),
.A2(n_641),
.B1(n_626),
.B2(n_648),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_790),
.Y(n_873)
);

AND3x1_ASAP7_75t_L g874 ( 
.A(n_776),
.B(n_334),
.C(n_320),
.Y(n_874)
);

AND2x4_ASAP7_75t_SL g875 ( 
.A(n_800),
.B(n_631),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_861),
.B(n_678),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_795),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_772),
.B(n_683),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_804),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_728),
.A2(n_683),
.B(n_612),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_713),
.A2(n_303),
.B1(n_321),
.B2(n_265),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_792),
.A2(n_303),
.B1(n_336),
.B2(n_321),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_723),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_738),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_804),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_741),
.B(n_733),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_712),
.B(n_612),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_723),
.B(n_551),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_790),
.B(n_636),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_711),
.B(n_293),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_741),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_772),
.B(n_811),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_733),
.B(n_618),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_708),
.B(n_637),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_811),
.B(n_249),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_704),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_781),
.A2(n_249),
.B1(n_257),
.B2(n_254),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_707),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_806),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_779),
.B(n_254),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_705),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_711),
.B(n_639),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_730),
.B(n_679),
.Y(n_903)
);

AND2x6_ASAP7_75t_SL g904 ( 
.A(n_739),
.B(n_335),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_806),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_731),
.A2(n_257),
.B1(n_267),
.B2(n_260),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_817),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_723),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_857),
.B(n_260),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_857),
.B(n_267),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_820),
.B(n_724),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_857),
.B(n_271),
.Y(n_912)
);

INVx8_ASAP7_75t_L g913 ( 
.A(n_723),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_817),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_708),
.B(n_687),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_823),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_853),
.A2(n_358),
.B(n_367),
.C(n_346),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_707),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_712),
.B(n_271),
.Y(n_919)
);

INVx8_ASAP7_75t_L g920 ( 
.A(n_764),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_712),
.B(n_272),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_721),
.B(n_272),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_760),
.B(n_273),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_760),
.B(n_273),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_760),
.B(n_275),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_716),
.B(n_275),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_838),
.B(n_372),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_808),
.A2(n_700),
.B(n_391),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_716),
.B(n_276),
.Y(n_929)
);

OAI22xp33_ASAP7_75t_L g930 ( 
.A1(n_853),
.A2(n_410),
.B1(n_432),
.B2(n_427),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_714),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_818),
.B(n_276),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_L g933 ( 
.A(n_860),
.B(n_384),
.C(n_375),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_731),
.A2(n_279),
.B1(n_281),
.B2(n_280),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_809),
.B(n_698),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_823),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_818),
.B(n_279),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_844),
.A2(n_762),
.B(n_767),
.C(n_858),
.Y(n_938)
);

INVx8_ASAP7_75t_L g939 ( 
.A(n_764),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_783),
.B(n_777),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_SL g941 ( 
.A1(n_866),
.A2(n_865),
.B(n_847),
.C(n_851),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_818),
.B(n_835),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_835),
.B(n_280),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_714),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_826),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_754),
.B(n_406),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_850),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_844),
.A2(n_392),
.B(n_401),
.C(n_385),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_718),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_737),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_718),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_726),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_835),
.B(n_281),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_850),
.B(n_303),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_726),
.Y(n_955)
);

INVx8_ASAP7_75t_L g956 ( 
.A(n_764),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_843),
.B(n_284),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_716),
.B(n_284),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_843),
.B(n_285),
.Y(n_959)
);

AND2x6_ASAP7_75t_SL g960 ( 
.A(n_739),
.B(n_402),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_705),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_725),
.B(n_285),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_826),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_750),
.B(n_289),
.Y(n_964)
);

NAND2x1p5_ASAP7_75t_L g965 ( 
.A(n_711),
.B(n_389),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_SL g966 ( 
.A1(n_717),
.A2(n_432),
.B1(n_440),
.B2(n_441),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_827),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_845),
.B(n_289),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_800),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_738),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_845),
.B(n_408),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_827),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_750),
.B(n_408),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_783),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_750),
.B(n_757),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_734),
.B(n_473),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_774),
.A2(n_847),
.B(n_839),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_755),
.B(n_321),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_762),
.B(n_767),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_800),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_762),
.B(n_767),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_793),
.A2(n_404),
.B(n_394),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_862),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_762),
.B(n_415),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_815),
.B(n_415),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_736),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_862),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_830),
.B(n_417),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_711),
.B(n_417),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_755),
.B(n_336),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_834),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_719),
.A2(n_752),
.B1(n_770),
.B2(n_756),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_736),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_834),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_710),
.Y(n_995)
);

NAND2x1_ASAP7_75t_L g996 ( 
.A(n_757),
.B(n_700),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_740),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_821),
.A2(n_400),
.B1(n_336),
.B2(n_351),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_756),
.B(n_440),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_752),
.B(n_420),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_789),
.B(n_420),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_825),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_757),
.B(n_421),
.Y(n_1003)
);

INVxp33_ASAP7_75t_L g1004 ( 
.A(n_813),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_789),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_829),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_810),
.B(n_421),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_810),
.B(n_433),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_816),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_759),
.B(n_441),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_740),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_813),
.B(n_446),
.Y(n_1012)
);

CKINVDCx11_ASAP7_75t_R g1013 ( 
.A(n_862),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_749),
.A2(n_451),
.B1(n_465),
.B2(n_463),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_816),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_821),
.A2(n_351),
.B1(n_400),
.B2(n_418),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_832),
.B(n_433),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_832),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_749),
.A2(n_449),
.B1(n_451),
.B2(n_454),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_846),
.B(n_434),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_755),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_846),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_759),
.B(n_434),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_856),
.B(n_438),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_856),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_836),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_821),
.A2(n_400),
.B1(n_351),
.B2(n_450),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_836),
.Y(n_1028)
);

NAND2xp33_ASAP7_75t_L g1029 ( 
.A(n_791),
.B(n_793),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_769),
.B(n_438),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_839),
.A2(n_447),
.B(n_424),
.C(n_419),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_759),
.B(n_445),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_807),
.B(n_445),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_807),
.B(n_803),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_709),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_739),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_807),
.B(n_449),
.Y(n_1037)
);

NAND3xp33_ASAP7_75t_L g1038 ( 
.A(n_746),
.B(n_467),
.C(n_446),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_755),
.B(n_467),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_749),
.A2(n_469),
.B1(n_454),
.B2(n_455),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_911),
.B(n_807),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1026),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1028),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_892),
.B(n_782),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_911),
.B(n_803),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_869),
.Y(n_1046)
);

NOR2xp67_ASAP7_75t_L g1047 ( 
.A(n_947),
.B(n_732),
.Y(n_1047)
);

AOI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_1004),
.A2(n_787),
.B(n_773),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_920),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_938),
.A2(n_854),
.B(n_855),
.C(n_851),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_891),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_974),
.B(n_742),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_869),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_913),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_915),
.B(n_802),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_876),
.B(n_803),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_896),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_867),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_877),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_927),
.B(n_884),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_878),
.B(n_942),
.Y(n_1061)
);

NAND2x2_ASAP7_75t_L g1062 ( 
.A(n_983),
.B(n_796),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_896),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_920),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_898),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_920),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_879),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_898),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_885),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_899),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_913),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_905),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_907),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_914),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_894),
.B(n_822),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_883),
.B(n_729),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_927),
.B(n_782),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_SL g1078 ( 
.A(n_974),
.B(n_470),
.C(n_837),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_920),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1002),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1002),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_979),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_933),
.A2(n_797),
.B1(n_966),
.B2(n_881),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_SL g1084 ( 
.A(n_930),
.B(n_470),
.C(n_840),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_916),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_946),
.B(n_742),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1021),
.B(n_782),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_936),
.Y(n_1088)
);

BUFx12f_ASAP7_75t_L g1089 ( 
.A(n_1013),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_SL g1090 ( 
.A(n_940),
.B(n_426),
.C(n_425),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_945),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_946),
.A2(n_796),
.B1(n_729),
.B2(n_859),
.Y(n_1092)
);

BUFx12f_ASAP7_75t_L g1093 ( 
.A(n_1013),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_918),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_963),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_967),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_972),
.Y(n_1097)
);

BUFx4f_ASAP7_75t_L g1098 ( 
.A(n_913),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_900),
.B(n_742),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_889),
.B(n_761),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_991),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_939),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_R g1103 ( 
.A(n_913),
.B(n_758),
.Y(n_1103)
);

OR2x4_ASAP7_75t_L g1104 ( 
.A(n_1012),
.B(n_854),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_939),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_884),
.B(n_785),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_935),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_939),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_969),
.B(n_768),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_939),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_956),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_902),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_868),
.A2(n_797),
.B1(n_824),
.B2(n_855),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_883),
.B(n_758),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_884),
.B(n_785),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_895),
.B(n_758),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_957),
.B(n_766),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_956),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_918),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_950),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_959),
.B(n_922),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1034),
.A2(n_797),
.B1(n_824),
.B2(n_864),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_931),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_956),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_994),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_886),
.B(n_797),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_873),
.B(n_552),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1004),
.B(n_785),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_902),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_931),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_944),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1009),
.Y(n_1133)
);

AND3x1_ASAP7_75t_SL g1134 ( 
.A(n_870),
.B(n_429),
.C(n_428),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_SL g1135 ( 
.A(n_1038),
.B(n_436),
.C(n_430),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_893),
.B(n_552),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1010),
.B(n_766),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_902),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_908),
.B(n_766),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_SL g1140 ( 
.A(n_903),
.B(n_824),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1015),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1018),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_875),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1010),
.B(n_801),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_956),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_908),
.B(n_801),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_888),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1022),
.Y(n_1148)
);

OR2x6_ASAP7_75t_L g1149 ( 
.A(n_888),
.B(n_780),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1035),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_962),
.B(n_801),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_944),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1025),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_970),
.B(n_791),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_983),
.B(n_709),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_949),
.Y(n_1156)
);

INVx6_ASAP7_75t_L g1157 ( 
.A(n_888),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_875),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_954),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_981),
.B(n_709),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_871),
.A2(n_865),
.B1(n_866),
.B2(n_864),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_949),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_970),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1035),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_951),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_976),
.B(n_706),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_992),
.B(n_799),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_951),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_978),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_987),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_952),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_990),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_SL g1173 ( 
.A(n_999),
.B(n_1031),
.C(n_917),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_995),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_R g1175 ( 
.A(n_987),
.B(n_838),
.Y(n_1175)
);

BUFx5_ASAP7_75t_L g1176 ( 
.A(n_1029),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_888),
.B(n_765),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1036),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_976),
.B(n_706),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_952),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_897),
.B(n_848),
.C(n_794),
.Y(n_1181)
);

BUFx4f_ASAP7_75t_L g1182 ( 
.A(n_890),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1006),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1039),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_961),
.Y(n_1185)
);

CKINVDCx8_ASAP7_75t_R g1186 ( 
.A(n_904),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_955),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_890),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_965),
.B(n_849),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_980),
.B(n_765),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_955),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_961),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1035),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_986),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_986),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_985),
.B(n_715),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_872),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_960),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_988),
.B(n_715),
.Y(n_1199)
);

CKINVDCx11_ASAP7_75t_R g1200 ( 
.A(n_961),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_993),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_SL g1202 ( 
.A(n_999),
.B(n_459),
.C(n_455),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1031),
.B(n_463),
.C(n_459),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_993),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_970),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_997),
.Y(n_1206)
);

INVx3_ASAP7_75t_SL g1207 ( 
.A(n_919),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_938),
.A2(n_971),
.B1(n_968),
.B2(n_937),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_997),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_923),
.Y(n_1210)
);

BUFx4f_ASAP7_75t_L g1211 ( 
.A(n_965),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1029),
.B(n_848),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_975),
.B(n_799),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1011),
.Y(n_1214)
);

AND2x6_ASAP7_75t_L g1215 ( 
.A(n_1011),
.B(n_720),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_977),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_901),
.Y(n_1217)
);

INVx5_ASAP7_75t_L g1218 ( 
.A(n_901),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_882),
.A2(n_748),
.B1(n_788),
.B2(n_720),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_932),
.B(n_722),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_943),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_953),
.B(n_722),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_924),
.B(n_747),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_874),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_909),
.B(n_747),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_996),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_1014),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_887),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_975),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_989),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_941),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1001),
.Y(n_1232)
);

BUFx12f_ASAP7_75t_L g1233 ( 
.A(n_917),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1228),
.A2(n_880),
.B(n_887),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1111),
.B(n_765),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1137),
.A2(n_941),
.B(n_921),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1216),
.A2(n_852),
.B(n_753),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1061),
.B(n_910),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1041),
.A2(n_984),
.B1(n_912),
.B2(n_1007),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1228),
.A2(n_928),
.B(n_753),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1045),
.B(n_925),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1113),
.A2(n_763),
.B(n_748),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1056),
.B(n_1033),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1136),
.B(n_1184),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1144),
.A2(n_921),
.B(n_919),
.Y(n_1245)
);

NAND2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1103),
.B(n_1212),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1210),
.B(n_1037),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1113),
.A2(n_788),
.B(n_763),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1121),
.A2(n_929),
.B(n_926),
.Y(n_1249)
);

OAI22x1_ASAP7_75t_L g1250 ( 
.A1(n_1197),
.A2(n_1040),
.B1(n_1019),
.B2(n_934),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1054),
.Y(n_1251)
);

NOR3xp33_ASAP7_75t_L g1252 ( 
.A(n_1048),
.B(n_1017),
.C(n_1008),
.Y(n_1252)
);

NOR2xp67_ASAP7_75t_L g1253 ( 
.A(n_1143),
.B(n_1020),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1122),
.A2(n_982),
.B(n_745),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1208),
.A2(n_948),
.B(n_743),
.C(n_751),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1122),
.A2(n_745),
.B(n_743),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1166),
.A2(n_929),
.B(n_926),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1128),
.B(n_1024),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1159),
.B(n_906),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1160),
.A2(n_964),
.B(n_958),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1044),
.A2(n_771),
.B(n_751),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1160),
.A2(n_964),
.B(n_958),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1128),
.B(n_1082),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1179),
.A2(n_1003),
.B(n_973),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1086),
.A2(n_1077),
.B(n_1151),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1181),
.A2(n_1003),
.B(n_973),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1044),
.A2(n_786),
.B(n_771),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_SL g1268 ( 
.A1(n_1163),
.A2(n_1000),
.B(n_786),
.Y(n_1268)
);

AND2x2_ASAP7_75t_SL g1269 ( 
.A(n_1211),
.B(n_998),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1167),
.A2(n_1223),
.B(n_1117),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1221),
.B(n_1016),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_L g1272 ( 
.A1(n_1231),
.A2(n_1032),
.B(n_1023),
.C(n_1077),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_L g1273 ( 
.A(n_1143),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1158),
.Y(n_1274)
);

AO21x2_ASAP7_75t_L g1275 ( 
.A1(n_1050),
.A2(n_1032),
.B(n_1023),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_SL g1276 ( 
.A1(n_1049),
.A2(n_735),
.B(n_727),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1230),
.B(n_1027),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1051),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1060),
.A2(n_819),
.B(n_814),
.Y(n_1279)
);

AOI221x1_ASAP7_75t_L g1280 ( 
.A1(n_1231),
.A2(n_948),
.B1(n_1030),
.B2(n_520),
.C(n_521),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1100),
.B(n_791),
.Y(n_1281)
);

AOI211x1_ASAP7_75t_L g1282 ( 
.A1(n_1042),
.A2(n_574),
.B(n_579),
.C(n_578),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1176),
.B(n_727),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1060),
.A2(n_819),
.B(n_814),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1043),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1050),
.A2(n_831),
.A3(n_833),
.B(n_574),
.Y(n_1286)
);

CKINVDCx8_ASAP7_75t_R g1287 ( 
.A(n_1158),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1174),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1126),
.B(n_791),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1058),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1099),
.A2(n_791),
.B(n_735),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1167),
.B(n_791),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1223),
.A2(n_828),
.B(n_842),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1196),
.A2(n_735),
.B(n_727),
.Y(n_1294)
);

OAI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1233),
.A2(n_563),
.B1(n_553),
.B2(n_559),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1232),
.A2(n_833),
.B(n_831),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1129),
.B(n_553),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1083),
.A2(n_422),
.B(n_409),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1232),
.A2(n_828),
.B(n_443),
.Y(n_1299)
);

OAI21xp33_ASAP7_75t_L g1300 ( 
.A1(n_1173),
.A2(n_469),
.B(n_465),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1169),
.B(n_764),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1084),
.B(n_444),
.C(n_435),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1176),
.B(n_727),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1199),
.A2(n_735),
.B(n_727),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1080),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1161),
.A2(n_828),
.B1(n_842),
.B2(n_744),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1232),
.A2(n_457),
.B(n_452),
.Y(n_1307)
);

AOI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_1055),
.A2(n_1107),
.B(n_1172),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1118),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1213),
.A2(n_744),
.B(n_735),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1220),
.A2(n_523),
.B(n_521),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1059),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1231),
.A2(n_562),
.A3(n_559),
.B(n_563),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1116),
.A2(n_842),
.B(n_764),
.Y(n_1314)
);

NOR2x1_ASAP7_75t_SL g1315 ( 
.A(n_1111),
.B(n_744),
.Y(n_1315)
);

NOR2xp67_ASAP7_75t_L g1316 ( 
.A(n_1075),
.B(n_841),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1127),
.B(n_1067),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1222),
.A2(n_764),
.B(n_841),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1225),
.A2(n_764),
.B(n_841),
.Y(n_1319)
);

AO22x1_ASAP7_75t_L g1320 ( 
.A1(n_1198),
.A2(n_562),
.B1(n_579),
.B2(n_578),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1089),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1089),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1046),
.A2(n_462),
.B(n_458),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1087),
.A2(n_841),
.B(n_812),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1213),
.A2(n_775),
.B(n_744),
.Y(n_1325)
);

OA22x2_ASAP7_75t_L g1326 ( 
.A1(n_1112),
.A2(n_577),
.B1(n_571),
.B2(n_568),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1087),
.A2(n_841),
.B(n_812),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1069),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1154),
.A2(n_532),
.B(n_523),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1070),
.B(n_1072),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1073),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_SL g1332 ( 
.A1(n_1163),
.A2(n_468),
.B(n_532),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1054),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1106),
.A2(n_841),
.B(n_812),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1053),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1111),
.B(n_765),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1053),
.A2(n_535),
.B(n_534),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1057),
.Y(n_1338)
);

OAI21xp33_ASAP7_75t_L g1339 ( 
.A1(n_1092),
.A2(n_310),
.B(n_307),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1161),
.A2(n_568),
.B(n_566),
.C(n_571),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1071),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1106),
.A2(n_744),
.B(n_775),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1057),
.A2(n_540),
.B(n_534),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1115),
.A2(n_775),
.B(n_863),
.Y(n_1344)
);

NOR2xp67_ASAP7_75t_L g1345 ( 
.A(n_1170),
.B(n_566),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1111),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1074),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1063),
.A2(n_577),
.A3(n_538),
.B(n_536),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1081),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1115),
.A2(n_805),
.B(n_812),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1085),
.B(n_775),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1154),
.A2(n_535),
.B(n_536),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1098),
.A2(n_775),
.B1(n_798),
.B2(n_784),
.Y(n_1353)
);

AOI221xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1083),
.A2(n_863),
.B1(n_798),
.B2(n_784),
.C(n_669),
.Y(n_1354)
);

OAI21xp33_ASAP7_75t_L g1355 ( 
.A1(n_1202),
.A2(n_371),
.B(n_311),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1176),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1088),
.A2(n_812),
.B(n_805),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1063),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1120),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1091),
.B(n_1095),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1098),
.A2(n_863),
.B(n_784),
.Y(n_1361)
);

AND2x6_ASAP7_75t_L g1362 ( 
.A(n_1118),
.B(n_784),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1226),
.A2(n_863),
.B(n_784),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1052),
.Y(n_1364)
);

AO32x2_ASAP7_75t_L g1365 ( 
.A1(n_1217),
.A2(n_812),
.A3(n_805),
.B1(n_778),
.B2(n_538),
.Y(n_1365)
);

NOR4xp25_ASAP7_75t_L g1366 ( 
.A(n_1090),
.B(n_539),
.C(n_540),
.D(n_541),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1096),
.B(n_778),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1049),
.A2(n_863),
.B(n_798),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1097),
.B(n_778),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1052),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1226),
.A2(n_798),
.B(n_312),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_SL g1372 ( 
.A1(n_1217),
.A2(n_541),
.B(n_539),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1176),
.B(n_798),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1176),
.B(n_778),
.Y(n_1374)
);

AO21x1_ASAP7_75t_L g1375 ( 
.A1(n_1140),
.A2(n_245),
.B(n_340),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1212),
.A2(n_805),
.B(n_812),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1065),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1101),
.B(n_11),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1170),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1125),
.B(n_12),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1149),
.A2(n_361),
.B(n_322),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1176),
.B(n_664),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1065),
.A2(n_1094),
.B(n_1068),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1211),
.B(n_12),
.Y(n_1384)
);

CKINVDCx6p67_ASAP7_75t_R g1385 ( 
.A(n_1093),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1093),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1068),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1094),
.A2(n_805),
.B(n_245),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1149),
.A2(n_364),
.B(n_324),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1131),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1071),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1119),
.A2(n_1130),
.B(n_1123),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1119),
.A2(n_805),
.B(n_245),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1118),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1176),
.B(n_664),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1149),
.A2(n_378),
.B(n_332),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1189),
.A2(n_379),
.B(n_347),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_SL g1398 ( 
.A1(n_1049),
.A2(n_15),
.B(n_16),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1182),
.B(n_17),
.Y(n_1399)
);

O2A1O1Ixp5_ASAP7_75t_L g1400 ( 
.A1(n_1205),
.A2(n_1164),
.B(n_1193),
.C(n_1150),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1265),
.A2(n_1102),
.B(n_1066),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1309),
.B(n_1155),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1235),
.Y(n_1403)
);

AND2x6_ASAP7_75t_L g1404 ( 
.A(n_1235),
.B(n_1177),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1234),
.A2(n_1130),
.B(n_1123),
.Y(n_1405)
);

BUFx12f_ASAP7_75t_L g1406 ( 
.A(n_1321),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1244),
.B(n_1183),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1288),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1270),
.B(n_1138),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1238),
.B(n_1233),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1285),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1359),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1234),
.A2(n_1237),
.B(n_1296),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1298),
.A2(n_1227),
.B1(n_1224),
.B2(n_1135),
.C(n_1078),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1296),
.A2(n_1152),
.B(n_1132),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1388),
.A2(n_1393),
.B(n_1284),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1278),
.Y(n_1417)
);

INVx6_ASAP7_75t_L g1418 ( 
.A(n_1309),
.Y(n_1418)
);

AO222x2_ASAP7_75t_L g1419 ( 
.A1(n_1259),
.A2(n_1186),
.B1(n_1134),
.B2(n_1227),
.C1(n_423),
.C2(n_1104),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1302),
.B(n_1252),
.C(n_1339),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1250),
.A2(n_1182),
.B1(n_1188),
.B2(n_1207),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_SL g1422 ( 
.A1(n_1258),
.A2(n_1205),
.B(n_1164),
.C(n_1150),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1383),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1309),
.B(n_1235),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1388),
.A2(n_1152),
.B(n_1132),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_SL g1426 ( 
.A(n_1287),
.B(n_1186),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1278),
.Y(n_1427)
);

AOI222xp33_ASAP7_75t_L g1428 ( 
.A1(n_1269),
.A2(n_1047),
.B1(n_1178),
.B2(n_1148),
.C1(n_1141),
.C2(n_1153),
.Y(n_1428)
);

NAND2x1p5_ASAP7_75t_L g1429 ( 
.A(n_1309),
.B(n_1177),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1317),
.B(n_1207),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1263),
.A2(n_1104),
.B1(n_1157),
.B2(n_1189),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1236),
.A2(n_1162),
.B(n_1156),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1349),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1305),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1356),
.A2(n_1189),
.B(n_1177),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1273),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1393),
.A2(n_1214),
.B(n_1187),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1279),
.A2(n_1214),
.B(n_1187),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1269),
.A2(n_1189),
.B1(n_1133),
.B2(n_1142),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1247),
.B(n_1109),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1336),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1246),
.A2(n_1218),
.B(n_1205),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1322),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1280),
.A2(n_1255),
.A3(n_1375),
.B(n_1245),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1295),
.A2(n_1157),
.B1(n_1171),
.B2(n_1194),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1336),
.B(n_1155),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1354),
.A2(n_1168),
.B(n_1165),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1323),
.A2(n_1191),
.B(n_1180),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1297),
.B(n_1241),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1345),
.A2(n_1157),
.B1(n_1147),
.B2(n_1200),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1290),
.B(n_1195),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1379),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1273),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1312),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1328),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1364),
.A2(n_1155),
.B1(n_1146),
.B2(n_1139),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1246),
.A2(n_1218),
.B(n_1164),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1276),
.B(n_1066),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1279),
.A2(n_1150),
.B(n_1193),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1370),
.B(n_1200),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1331),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_SL g1462 ( 
.A1(n_1277),
.A2(n_1175),
.B1(n_1062),
.B2(n_1203),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1271),
.A2(n_1175),
.B1(n_1062),
.B2(n_1114),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1300),
.A2(n_1219),
.B1(n_1193),
.B2(n_1229),
.C(n_1218),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1330),
.B(n_1139),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1336),
.Y(n_1466)
);

AOI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1382),
.A2(n_1209),
.B(n_1204),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1284),
.A2(n_1206),
.B(n_1201),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_SL g1469 ( 
.A(n_1274),
.B(n_1190),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1383),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1243),
.A2(n_1360),
.B1(n_1399),
.B2(n_1384),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1308),
.B(n_1139),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1392),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1385),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1281),
.A2(n_1146),
.B1(n_1076),
.B2(n_1229),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_SL g1476 ( 
.A(n_1346),
.B(n_1124),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1391),
.B(n_1076),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1239),
.A2(n_1146),
.B(n_1076),
.C(n_1190),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1295),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1392),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1274),
.B(n_1190),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1323),
.A2(n_1219),
.B(n_1215),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1346),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1249),
.A2(n_1064),
.B(n_1079),
.C(n_1105),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1391),
.B(n_1124),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1242),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_SL g1487 ( 
.A1(n_1268),
.A2(n_1266),
.B(n_1292),
.Y(n_1487)
);

NAND3xp33_ASAP7_75t_L g1488 ( 
.A(n_1355),
.B(n_1229),
.C(n_1218),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1347),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1251),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1260),
.A2(n_1229),
.B1(n_1066),
.B2(n_1102),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1261),
.A2(n_1110),
.B(n_1108),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1351),
.Y(n_1493)
);

INVx3_ASAP7_75t_SL g1494 ( 
.A(n_1321),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1390),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_SL g1496 ( 
.A1(n_1262),
.A2(n_1102),
.B(n_1079),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_SL g1497 ( 
.A1(n_1373),
.A2(n_1064),
.B(n_1105),
.C(n_1145),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1257),
.A2(n_1215),
.B(n_1110),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1255),
.A2(n_1114),
.B(n_1215),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1378),
.B(n_1185),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1322),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1368),
.B(n_1118),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1253),
.A2(n_1192),
.B1(n_1185),
.B2(n_1108),
.C(n_1145),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1261),
.A2(n_1108),
.B(n_1110),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1326),
.A2(n_1215),
.B1(n_1192),
.B2(n_1185),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1335),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1264),
.A2(n_1215),
.B(n_1103),
.Y(n_1507)
);

AO31x2_ASAP7_75t_L g1508 ( 
.A1(n_1340),
.A2(n_1192),
.A3(n_1185),
.B(n_664),
.Y(n_1508)
);

AO31x2_ASAP7_75t_L g1509 ( 
.A1(n_1340),
.A2(n_1192),
.A3(n_664),
.B(n_669),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1272),
.A2(n_1145),
.B(n_1124),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1335),
.Y(n_1511)
);

INVxp67_ASAP7_75t_L g1512 ( 
.A(n_1380),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1326),
.A2(n_1124),
.B1(n_805),
.B2(n_669),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1267),
.A2(n_317),
.B(n_403),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1338),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1316),
.A2(n_348),
.B1(n_387),
.B2(n_669),
.Y(n_1516)
);

CKINVDCx8_ASAP7_75t_R g1517 ( 
.A(n_1251),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1289),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1346),
.B(n_664),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1267),
.A2(n_245),
.B(n_340),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1358),
.Y(n_1521)
);

INVx3_ASAP7_75t_SL g1522 ( 
.A(n_1386),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1377),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1251),
.B(n_664),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1293),
.A2(n_669),
.B1(n_412),
.B2(n_357),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1240),
.A2(n_340),
.B(n_245),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1240),
.A2(n_340),
.B(n_245),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1299),
.A2(n_1343),
.B(n_1337),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1320),
.B(n_20),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1299),
.A2(n_340),
.B(n_669),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1251),
.B(n_20),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1387),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1337),
.A2(n_340),
.B(n_357),
.Y(n_1533)
);

AOI222xp33_ASAP7_75t_L g1534 ( 
.A1(n_1301),
.A2(n_412),
.B1(n_357),
.B2(n_350),
.C1(n_264),
.C2(n_248),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1242),
.B(n_21),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1387),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1343),
.A2(n_1303),
.B(n_1283),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1283),
.A2(n_340),
.B(n_357),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1248),
.B(n_23),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1307),
.A2(n_340),
.B(n_357),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1256),
.Y(n_1541)
);

AOI211xp5_ASAP7_75t_L g1542 ( 
.A1(n_1397),
.A2(n_412),
.B(n_350),
.C(n_264),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1348),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1303),
.A2(n_412),
.B(n_350),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1248),
.B(n_25),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1307),
.A2(n_412),
.B(n_350),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1348),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1256),
.Y(n_1548)
);

AOI22x1_ASAP7_75t_L g1549 ( 
.A1(n_1291),
.A2(n_350),
.B1(n_264),
.B2(n_248),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1373),
.A2(n_1395),
.B(n_1382),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_SL g1551 ( 
.A1(n_1332),
.A2(n_26),
.B(n_27),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1348),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1275),
.A2(n_1396),
.B1(n_1389),
.B2(n_1381),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1400),
.A2(n_27),
.B(n_28),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1286),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1348),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1286),
.B(n_32),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1318),
.A2(n_264),
.B(n_238),
.Y(n_1558)
);

AO21x2_ASAP7_75t_L g1559 ( 
.A1(n_1319),
.A2(n_264),
.B(n_226),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1395),
.A2(n_224),
.B(n_220),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1333),
.B(n_35),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1374),
.B(n_35),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1333),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1294),
.A2(n_219),
.B(n_211),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1286),
.B(n_38),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1304),
.A2(n_210),
.B(n_204),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1282),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1362),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1286),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1333),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1374),
.B(n_39),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1275),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_1572)
);

AOI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1310),
.A2(n_200),
.B(n_192),
.Y(n_1573)
);

AO21x2_ASAP7_75t_L g1574 ( 
.A1(n_1314),
.A2(n_190),
.B(n_189),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1325),
.A2(n_1254),
.B(n_1342),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1254),
.A2(n_187),
.B(n_184),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1362),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1313),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1333),
.B(n_40),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1311),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1479),
.A2(n_1311),
.B1(n_1398),
.B2(n_1386),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1471),
.A2(n_1366),
.B1(n_1371),
.B2(n_1372),
.C(n_1306),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1449),
.B(n_48),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1435),
.B(n_1341),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1495),
.Y(n_1585)
);

BUFx10_ASAP7_75t_L g1586 ( 
.A(n_1474),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1417),
.B(n_1313),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1449),
.B(n_50),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1511),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1408),
.Y(n_1590)
);

OAI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1529),
.A2(n_1571),
.B1(n_1562),
.B2(n_1469),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1412),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1517),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1410),
.B(n_1341),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1410),
.B(n_53),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1411),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1463),
.A2(n_1420),
.B1(n_1462),
.B2(n_1434),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_SL g1598 ( 
.A(n_1562),
.B(n_1341),
.Y(n_1598)
);

BUFx12f_ASAP7_75t_L g1599 ( 
.A(n_1501),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1511),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1414),
.A2(n_1369),
.B1(n_1367),
.B2(n_1341),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_SL g1602 ( 
.A1(n_1554),
.A2(n_1315),
.B(n_1344),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_1501),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1562),
.A2(n_1324),
.B1(n_1327),
.B2(n_1394),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1412),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1465),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1427),
.B(n_1394),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1454),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1428),
.A2(n_1419),
.B1(n_1409),
.B2(n_1512),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1403),
.B(n_1394),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1441),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1455),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1436),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1407),
.B(n_1394),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1517),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1409),
.B(n_1313),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1490),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1481),
.B(n_1579),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1443),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1555),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1555),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1403),
.B(n_1362),
.Y(n_1622)
);

INVx4_ASAP7_75t_L g1623 ( 
.A(n_1436),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1579),
.B(n_1430),
.Y(n_1624)
);

OAI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1572),
.A2(n_1439),
.B1(n_1518),
.B2(n_1421),
.C(n_1450),
.Y(n_1625)
);

AOI222xp33_ASAP7_75t_L g1626 ( 
.A1(n_1419),
.A2(n_1357),
.B1(n_1350),
.B2(n_1334),
.C1(n_1362),
.C2(n_62),
.Y(n_1626)
);

CKINVDCx11_ASAP7_75t_R g1627 ( 
.A(n_1443),
.Y(n_1627)
);

NOR2xp67_ASAP7_75t_L g1628 ( 
.A(n_1452),
.B(n_1361),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1494),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1461),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1489),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1526),
.A2(n_1363),
.B(n_1329),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1440),
.B(n_1362),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1441),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1451),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1441),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1451),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1494),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1413),
.A2(n_1352),
.B(n_1353),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1431),
.A2(n_1376),
.B1(n_1313),
.B2(n_1365),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1433),
.B(n_54),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1460),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1506),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1490),
.Y(n_1644)
);

OAI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1562),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1472),
.B(n_56),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1522),
.B(n_57),
.Y(n_1647)
);

BUFx4f_ASAP7_75t_SL g1648 ( 
.A(n_1406),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1406),
.Y(n_1649)
);

AOI222xp33_ASAP7_75t_L g1650 ( 
.A1(n_1464),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.C1(n_67),
.C2(n_68),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1413),
.A2(n_1365),
.B(n_1376),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1535),
.A2(n_1365),
.B1(n_69),
.B2(n_73),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_SL g1653 ( 
.A1(n_1457),
.A2(n_1442),
.B(n_1577),
.C(n_1568),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1477),
.B(n_68),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1402),
.Y(n_1655)
);

NAND4xp25_ASAP7_75t_L g1656 ( 
.A(n_1567),
.B(n_69),
.C(n_73),
.D(n_74),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1515),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1521),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1571),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1477),
.B(n_79),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1525),
.A2(n_1365),
.B(n_80),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1477),
.B(n_79),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1535),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_1663)
);

INVx3_ASAP7_75t_SL g1664 ( 
.A(n_1474),
.Y(n_1664)
);

CKINVDCx11_ASAP7_75t_R g1665 ( 
.A(n_1522),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1571),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_1666)
);

AOI21xp33_ASAP7_75t_L g1667 ( 
.A1(n_1534),
.A2(n_84),
.B(n_88),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1402),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1446),
.B(n_84),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1580),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.C(n_92),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1526),
.A2(n_115),
.B(n_169),
.Y(n_1671)
);

OAI21x1_ASAP7_75t_L g1672 ( 
.A1(n_1527),
.A2(n_111),
.B(n_160),
.Y(n_1672)
);

NAND2x1p5_ASAP7_75t_L g1673 ( 
.A(n_1424),
.B(n_172),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_R g1674 ( 
.A(n_1568),
.B(n_155),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1446),
.B(n_89),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1571),
.A2(n_90),
.B1(n_91),
.B2(n_95),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1403),
.B(n_122),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1557),
.B(n_96),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1523),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1532),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1446),
.B(n_97),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1539),
.A2(n_98),
.B1(n_99),
.B2(n_104),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1441),
.B(n_139),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1453),
.B(n_98),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1453),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1563),
.B(n_104),
.Y(n_1686)
);

OR2x6_ASAP7_75t_L g1687 ( 
.A(n_1478),
.B(n_134),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1539),
.A2(n_107),
.B1(n_153),
.B2(n_151),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1493),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1441),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1536),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1422),
.A2(n_107),
.B(n_149),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1424),
.Y(n_1693)
);

AOI221x1_ASAP7_75t_L g1694 ( 
.A1(n_1551),
.A2(n_1488),
.B1(n_1545),
.B2(n_1531),
.C(n_1561),
.Y(n_1694)
);

OAI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1545),
.A2(n_1553),
.B(n_1557),
.C(n_1565),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1486),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1551),
.A2(n_152),
.B1(n_1565),
.B2(n_1569),
.C(n_1500),
.Y(n_1697)
);

OAI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1505),
.A2(n_1426),
.B1(n_1456),
.B2(n_1568),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1491),
.B(n_1475),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1405),
.Y(n_1700)
);

NAND2xp33_ASAP7_75t_R g1701 ( 
.A(n_1577),
.B(n_1482),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1542),
.B(n_1445),
.C(n_1516),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1513),
.A2(n_1577),
.B1(n_1402),
.B2(n_1483),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1499),
.A2(n_1559),
.B1(n_1558),
.B2(n_1482),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1570),
.B(n_1466),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1424),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1466),
.B(n_1429),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1466),
.B(n_1483),
.Y(n_1708)
);

AOI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1558),
.A2(n_1559),
.B(n_1514),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1418),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1486),
.A2(n_1429),
.B1(n_1503),
.B2(n_1418),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1405),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1418),
.Y(n_1713)
);

AO21x2_ASAP7_75t_L g1714 ( 
.A1(n_1578),
.A2(n_1552),
.B(n_1556),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1404),
.A2(n_1499),
.B1(n_1418),
.B2(n_1485),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_R g1716 ( 
.A(n_1404),
.B(n_1483),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1543),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1547),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1423),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1404),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1404),
.A2(n_1499),
.B1(n_1485),
.B2(n_1559),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1404),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1485),
.B(n_1524),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1502),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1524),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1423),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1498),
.A2(n_1484),
.B(n_1510),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1482),
.A2(n_1558),
.B1(n_1574),
.B2(n_1578),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1574),
.A2(n_1447),
.B1(n_1448),
.B2(n_1514),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1447),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1519),
.B(n_1508),
.Y(n_1731)
);

AOI22x1_ASAP7_75t_L g1732 ( 
.A1(n_1487),
.A2(n_1401),
.B1(n_1496),
.B2(n_1519),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1733)
);

AO31x2_ASAP7_75t_L g1734 ( 
.A1(n_1541),
.A2(n_1548),
.A3(n_1473),
.B(n_1470),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1502),
.B(n_1458),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1502),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_SL g1737 ( 
.A1(n_1574),
.A2(n_1507),
.B1(n_1546),
.B2(n_1514),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1519),
.B(n_1447),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1422),
.B(n_1507),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1502),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1573),
.A2(n_1497),
.B(n_1549),
.C(n_1560),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1576),
.A2(n_1564),
.B(n_1566),
.C(n_1560),
.Y(n_1742)
);

OAI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1458),
.A2(n_1548),
.B1(n_1541),
.B2(n_1546),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1745)
);

NOR3xp33_ASAP7_75t_SL g1746 ( 
.A(n_1487),
.B(n_1497),
.C(n_1496),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1468),
.Y(n_1747)
);

BUFx12f_ASAP7_75t_L g1748 ( 
.A(n_1458),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1458),
.A2(n_1467),
.B1(n_1448),
.B2(n_1546),
.Y(n_1749)
);

NOR2x1_ASAP7_75t_L g1750 ( 
.A(n_1507),
.B(n_1432),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1432),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1448),
.A2(n_1432),
.B1(n_1540),
.B2(n_1576),
.Y(n_1753)
);

AOI21x1_ASAP7_75t_L g1754 ( 
.A1(n_1527),
.A2(n_1540),
.B(n_1544),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1470),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1468),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1540),
.A2(n_1480),
.B1(n_1473),
.B2(n_1438),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1509),
.B(n_1476),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1480),
.A2(n_1550),
.B1(n_1444),
.B2(n_1401),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1438),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1444),
.B(n_1550),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1444),
.B(n_1459),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1564),
.Y(n_1763)
);

BUFx3_ASAP7_75t_L g1764 ( 
.A(n_1459),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1415),
.Y(n_1765)
);

INVx6_ASAP7_75t_L g1766 ( 
.A(n_1566),
.Y(n_1766)
);

AO21x2_ASAP7_75t_L g1767 ( 
.A1(n_1520),
.A2(n_1416),
.B(n_1425),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1444),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1415),
.Y(n_1769)
);

OR2x6_ASAP7_75t_L g1770 ( 
.A(n_1425),
.B(n_1437),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1537),
.B(n_1504),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1444),
.A2(n_1537),
.B1(n_1575),
.B2(n_1544),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1437),
.B(n_1538),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1538),
.A2(n_1575),
.B1(n_1533),
.B2(n_1530),
.C(n_1528),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1530),
.A2(n_1492),
.B1(n_1504),
.B2(n_1528),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1533),
.A2(n_1416),
.B1(n_1492),
.B2(n_1520),
.Y(n_1776)
);

OAI21x1_ASAP7_75t_L g1777 ( 
.A1(n_1413),
.A2(n_1527),
.B(n_1526),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1449),
.B(n_1410),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_SL g1779 ( 
.A(n_1414),
.B(n_940),
.C(n_610),
.Y(n_1779)
);

BUFx4f_ASAP7_75t_SL g1780 ( 
.A(n_1599),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_SL g1781 ( 
.A1(n_1625),
.A2(n_1695),
.B1(n_1687),
.B2(n_1597),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1663),
.A2(n_1682),
.B1(n_1645),
.B2(n_1666),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1596),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1644),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1687),
.A2(n_1598),
.B1(n_1678),
.B2(n_1646),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1656),
.B2(n_1591),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1593),
.Y(n_1787)
);

INVx4_ASAP7_75t_L g1788 ( 
.A(n_1685),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1591),
.A2(n_1779),
.B1(n_1659),
.B2(n_1666),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1618),
.B(n_1624),
.Y(n_1790)
);

OA21x2_ASAP7_75t_L g1791 ( 
.A1(n_1709),
.A2(n_1729),
.B(n_1742),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1663),
.A2(n_1682),
.B1(n_1609),
.B2(n_1697),
.C(n_1650),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1608),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1645),
.A2(n_1676),
.B1(n_1659),
.B2(n_1702),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1676),
.A2(n_1687),
.B1(n_1667),
.B2(n_1670),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1612),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1630),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1631),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1585),
.Y(n_1799)
);

BUFx5_ASAP7_75t_L g1800 ( 
.A(n_1764),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1688),
.A2(n_1652),
.B1(n_1642),
.B2(n_1604),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1652),
.A2(n_1688),
.B1(n_1778),
.B2(n_1583),
.C(n_1588),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1696),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1698),
.A2(n_1606),
.B1(n_1595),
.B2(n_1604),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1643),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_SL g1806 ( 
.A1(n_1716),
.A2(n_1722),
.B1(n_1748),
.B2(n_1661),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1658),
.Y(n_1807)
);

AOI21xp33_ASAP7_75t_L g1808 ( 
.A1(n_1587),
.A2(n_1581),
.B(n_1633),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1592),
.B(n_1605),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_SL g1810 ( 
.A1(n_1716),
.A2(n_1722),
.B1(n_1748),
.B2(n_1727),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1627),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1698),
.A2(n_1704),
.B1(n_1616),
.B2(n_1699),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1644),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1641),
.A2(n_1581),
.B1(n_1768),
.B2(n_1582),
.C(n_1689),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1619),
.A2(n_1601),
.B1(n_1660),
.B2(n_1662),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1617),
.B(n_1681),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1742),
.A2(n_1653),
.B(n_1741),
.Y(n_1818)
);

OAI211xp5_ASAP7_75t_L g1819 ( 
.A1(n_1694),
.A2(n_1654),
.B(n_1675),
.C(n_1669),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1679),
.Y(n_1820)
);

OAI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1674),
.A2(n_1594),
.B1(n_1619),
.B2(n_1722),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1614),
.B(n_1590),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1699),
.A2(n_1601),
.B1(n_1647),
.B2(n_1627),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1599),
.A2(n_1722),
.B1(n_1728),
.B2(n_1684),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1674),
.A2(n_1715),
.B1(n_1673),
.B2(n_1721),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1607),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1705),
.B(n_1680),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1696),
.Y(n_1828)
);

OAI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1673),
.A2(n_1648),
.B1(n_1615),
.B2(n_1720),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1728),
.A2(n_1737),
.B1(n_1711),
.B2(n_1665),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1711),
.A2(n_1665),
.B1(n_1717),
.B2(n_1718),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_SL g1832 ( 
.A1(n_1744),
.A2(n_1766),
.B1(n_1735),
.B2(n_1731),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1729),
.A2(n_1745),
.B1(n_1739),
.B2(n_1692),
.C(n_1738),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1649),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1706),
.B(n_1693),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1739),
.A2(n_1686),
.B1(n_1752),
.B2(n_1761),
.C(n_1730),
.Y(n_1836)
);

BUFx8_ASAP7_75t_SL g1837 ( 
.A(n_1603),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_SL g1838 ( 
.A1(n_1766),
.A2(n_1735),
.B1(n_1720),
.B2(n_1740),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1638),
.A2(n_1735),
.B(n_1622),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1752),
.A2(n_1640),
.B1(n_1762),
.B2(n_1759),
.C(n_1751),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1747),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_SL g1842 ( 
.A1(n_1766),
.A2(n_1740),
.B1(n_1724),
.B2(n_1736),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_L g1843 ( 
.A(n_1628),
.B(n_1746),
.C(n_1750),
.Y(n_1843)
);

OAI31xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1732),
.A2(n_1703),
.A3(n_1677),
.B(n_1683),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1640),
.A2(n_1648),
.B1(n_1657),
.B2(n_1691),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1724),
.A2(n_1736),
.B1(n_1683),
.B2(n_1733),
.Y(n_1846)
);

BUFx3_ASAP7_75t_L g1847 ( 
.A(n_1685),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1691),
.A2(n_1603),
.B1(n_1736),
.B2(n_1724),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1693),
.B(n_1708),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1629),
.A2(n_1613),
.B1(n_1623),
.B2(n_1664),
.Y(n_1850)
);

OAI33xp33_ASAP7_75t_L g1851 ( 
.A1(n_1772),
.A2(n_1749),
.A3(n_1758),
.B1(n_1690),
.B2(n_1743),
.B3(n_1775),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_SL g1852 ( 
.A1(n_1736),
.A2(n_1683),
.B1(n_1677),
.B2(n_1763),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1584),
.A2(n_1677),
.B1(n_1589),
.B2(n_1600),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1723),
.B(n_1655),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1655),
.B(n_1668),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1756),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1664),
.A2(n_1668),
.B1(n_1622),
.B2(n_1713),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1622),
.A2(n_1610),
.B1(n_1710),
.B2(n_1725),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1714),
.A2(n_1707),
.B1(n_1719),
.B2(n_1726),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1763),
.A2(n_1602),
.B1(n_1701),
.B2(n_1671),
.Y(n_1860)
);

AOI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1743),
.A2(n_1753),
.B1(n_1757),
.B2(n_1726),
.C(n_1719),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1611),
.B(n_1636),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1714),
.A2(n_1755),
.B1(n_1610),
.B2(n_1621),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1755),
.A2(n_1610),
.B1(n_1620),
.B2(n_1621),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1611),
.A2(n_1636),
.B1(n_1634),
.B2(n_1586),
.Y(n_1865)
);

BUFx12f_ASAP7_75t_L g1866 ( 
.A(n_1586),
.Y(n_1866)
);

AOI222xp33_ASAP7_75t_L g1867 ( 
.A1(n_1765),
.A2(n_1760),
.B1(n_1634),
.B2(n_1636),
.C1(n_1757),
.C2(n_1774),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1776),
.A2(n_1764),
.B1(n_1773),
.B2(n_1771),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1653),
.A2(n_1672),
.B1(n_1770),
.B2(n_1771),
.Y(n_1869)
);

AOI222xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1700),
.A2(n_1712),
.B1(n_1769),
.B2(n_1771),
.C1(n_1776),
.C2(n_1777),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1651),
.B(n_1770),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1734),
.B(n_1770),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_SL g1873 ( 
.A1(n_1632),
.A2(n_1767),
.B1(n_1639),
.B2(n_1734),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1734),
.B(n_1767),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1632),
.A2(n_1626),
.B1(n_1609),
.B2(n_1233),
.Y(n_1875)
);

OAI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1632),
.A2(n_1656),
.B1(n_717),
.B2(n_940),
.C(n_635),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1635),
.B(n_1417),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1685),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1618),
.B(n_1624),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1596),
.Y(n_1881)
);

OAI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1656),
.A2(n_1298),
.B1(n_1479),
.B2(n_1645),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1596),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1592),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1596),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1635),
.B(n_1417),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1604),
.A2(n_1356),
.B(n_1270),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1635),
.B(n_1417),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1778),
.B(n_1585),
.Y(n_1891)
);

OAI221xp5_ASAP7_75t_L g1892 ( 
.A1(n_1656),
.A2(n_717),
.B1(n_940),
.B2(n_635),
.C(n_881),
.Y(n_1892)
);

OAI21x1_ASAP7_75t_L g1893 ( 
.A1(n_1754),
.A2(n_1413),
.B(n_1777),
.Y(n_1893)
);

OR2x6_ASAP7_75t_L g1894 ( 
.A(n_1748),
.B(n_1735),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1754),
.A2(n_1413),
.B(n_1777),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1635),
.B(n_1417),
.Y(n_1896)
);

OA21x2_ASAP7_75t_L g1897 ( 
.A1(n_1709),
.A2(n_1729),
.B(n_1742),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1592),
.Y(n_1898)
);

AO31x2_ASAP7_75t_L g1899 ( 
.A1(n_1749),
.A2(n_1742),
.A3(n_1578),
.B(n_1739),
.Y(n_1899)
);

OAI211xp5_ASAP7_75t_L g1900 ( 
.A1(n_1656),
.A2(n_1682),
.B(n_1663),
.C(n_853),
.Y(n_1900)
);

OAI221xp5_ASAP7_75t_L g1901 ( 
.A1(n_1656),
.A2(n_717),
.B1(n_940),
.B2(n_635),
.C(n_881),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1619),
.A2(n_1603),
.B1(n_1443),
.B2(n_1609),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_SL g1903 ( 
.A1(n_1625),
.A2(n_1695),
.B1(n_487),
.B2(n_489),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1618),
.B(n_1624),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1625),
.A2(n_1695),
.B1(n_487),
.B2(n_489),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1656),
.A2(n_1298),
.B1(n_1479),
.B2(n_1645),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1635),
.B(n_1417),
.Y(n_1907)
);

CKINVDCx20_ASAP7_75t_R g1908 ( 
.A(n_1603),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1909)
);

OAI322xp33_ASAP7_75t_L g1910 ( 
.A1(n_1645),
.A2(n_261),
.A3(n_1659),
.B1(n_1676),
.B2(n_1666),
.C1(n_930),
.C2(n_635),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1618),
.B(n_1624),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_SL g1912 ( 
.A1(n_1625),
.A2(n_1695),
.B1(n_487),
.B2(n_489),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1696),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1663),
.A2(n_1682),
.B1(n_1597),
.B2(n_1479),
.Y(n_1914)
);

OAI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1656),
.A2(n_713),
.B(n_1420),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1618),
.B(n_1624),
.Y(n_1916)
);

AOI222xp33_ASAP7_75t_L g1917 ( 
.A1(n_1609),
.A2(n_1298),
.B1(n_966),
.B2(n_881),
.C1(n_1233),
.C2(n_676),
.Y(n_1917)
);

OR2x6_ASAP7_75t_L g1918 ( 
.A(n_1748),
.B(n_1735),
.Y(n_1918)
);

OAI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1656),
.A2(n_1298),
.B1(n_1479),
.B2(n_1645),
.Y(n_1919)
);

AOI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1604),
.A2(n_1356),
.B(n_1270),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1663),
.A2(n_1682),
.B1(n_1597),
.B2(n_1479),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_L g1923 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1663),
.A2(n_1682),
.B1(n_1597),
.B2(n_1479),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1696),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1656),
.A2(n_717),
.B1(n_940),
.B2(n_635),
.C(n_881),
.Y(n_1928)
);

AOI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1645),
.A2(n_930),
.B1(n_719),
.B2(n_717),
.C(n_966),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1626),
.A2(n_1609),
.B1(n_1233),
.B2(n_1656),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1627),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1604),
.A2(n_1356),
.B(n_1270),
.Y(n_1932)
);

AOI21xp33_ASAP7_75t_L g1933 ( 
.A1(n_1626),
.A2(n_1471),
.B(n_1420),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1597),
.B(n_1656),
.Y(n_1934)
);

OAI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1656),
.A2(n_717),
.B1(n_940),
.B2(n_635),
.C(n_881),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1627),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1656),
.A2(n_713),
.B(n_1420),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1596),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1644),
.Y(n_1939)
);

OAI21xp33_ASAP7_75t_L g1940 ( 
.A1(n_1656),
.A2(n_1682),
.B(n_1663),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1618),
.B(n_1624),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1800),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1871),
.B(n_1899),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1809),
.B(n_1803),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1841),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1803),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1856),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1828),
.B(n_1913),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1828),
.B(n_1913),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1814),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1927),
.Y(n_1951)
);

BUFx2_ASAP7_75t_L g1952 ( 
.A(n_1927),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1799),
.B(n_1783),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1856),
.Y(n_1954)
);

INVxp67_ASAP7_75t_SL g1955 ( 
.A(n_1874),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1891),
.B(n_1827),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1793),
.B(n_1796),
.Y(n_1957)
);

NOR2x1_ASAP7_75t_L g1958 ( 
.A(n_1843),
.B(n_1814),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1899),
.B(n_1791),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1898),
.B(n_1872),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1788),
.B(n_1878),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1797),
.B(n_1798),
.Y(n_1962)
);

INVx4_ASAP7_75t_L g1963 ( 
.A(n_1784),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1805),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1899),
.B(n_1791),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1836),
.B(n_1881),
.Y(n_1966)
);

INVxp67_ASAP7_75t_SL g1967 ( 
.A(n_1791),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1899),
.B(n_1897),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1807),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1897),
.B(n_1873),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1820),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1884),
.B(n_1886),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1897),
.B(n_1868),
.Y(n_1973)
);

OAI21x1_ASAP7_75t_L g1974 ( 
.A1(n_1818),
.A2(n_1895),
.B(n_1893),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1938),
.Y(n_1975)
);

AO31x2_ASAP7_75t_L g1976 ( 
.A1(n_1801),
.A2(n_1889),
.A3(n_1932),
.B(n_1921),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1790),
.B(n_1880),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1904),
.B(n_1911),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1916),
.B(n_1941),
.Y(n_1979)
);

INVxp67_ASAP7_75t_L g1980 ( 
.A(n_1870),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1833),
.B(n_1867),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1939),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1826),
.B(n_1811),
.Y(n_1983)
);

AOI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1929),
.A2(n_1940),
.B1(n_1786),
.B2(n_1934),
.C(n_1792),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1939),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_SL g1986 ( 
.A1(n_1782),
.A2(n_1900),
.B1(n_1914),
.B2(n_1924),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1885),
.B(n_1877),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1887),
.B(n_1890),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1840),
.B(n_1869),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1896),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1832),
.B(n_1817),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1861),
.B(n_1860),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1859),
.B(n_1863),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1907),
.B(n_1813),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1859),
.B(n_1863),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1849),
.B(n_1835),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1813),
.B(n_1822),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1784),
.Y(n_1998)
);

OAI31xp33_ASAP7_75t_L g1999 ( 
.A1(n_1934),
.A2(n_1922),
.A3(n_1928),
.B(n_1901),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1849),
.B(n_1854),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1862),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1808),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1864),
.Y(n_2003)
);

OA21x2_ASAP7_75t_L g2004 ( 
.A1(n_1830),
.A2(n_1845),
.B(n_1831),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1845),
.B(n_1830),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1788),
.B(n_1878),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1857),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1812),
.B(n_1847),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1787),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1894),
.B(n_1918),
.Y(n_2010)
);

OAI221xp5_ASAP7_75t_L g2011 ( 
.A1(n_1786),
.A2(n_1923),
.B1(n_1883),
.B2(n_1879),
.C(n_1909),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1858),
.Y(n_2012)
);

OA21x2_ASAP7_75t_L g2013 ( 
.A1(n_1831),
.A2(n_1853),
.B(n_1815),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1908),
.B(n_1837),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1844),
.B(n_1853),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1931),
.B(n_1936),
.Y(n_2016)
);

AO21x2_ASAP7_75t_L g2017 ( 
.A1(n_1825),
.A2(n_1789),
.B(n_1933),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1804),
.B(n_1855),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1825),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1781),
.B(n_1804),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1794),
.B(n_1838),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_L g2022 ( 
.A1(n_1903),
.A2(n_1912),
.B1(n_1905),
.B2(n_1917),
.Y(n_2022)
);

INVxp67_ASAP7_75t_SL g2023 ( 
.A(n_1821),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1839),
.Y(n_2024)
);

NAND2xp33_ASAP7_75t_R g2025 ( 
.A(n_2014),
.B(n_1834),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1944),
.B(n_1824),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_2016),
.B(n_1780),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1981),
.A2(n_1794),
.B1(n_1875),
.B2(n_1902),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1944),
.B(n_1824),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_1949),
.B(n_1816),
.Y(n_2030)
);

OAI321xp33_ASAP7_75t_L g2031 ( 
.A1(n_1981),
.A2(n_1876),
.A3(n_1935),
.B1(n_1892),
.B2(n_1926),
.C(n_1925),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_2008),
.B(n_1780),
.Y(n_2032)
);

AOI33xp33_ASAP7_75t_L g2033 ( 
.A1(n_1986),
.A2(n_1920),
.A3(n_1883),
.B1(n_1888),
.B2(n_1930),
.B3(n_1926),
.Y(n_2033)
);

INVxp67_ASAP7_75t_L g2034 ( 
.A(n_1990),
.Y(n_2034)
);

OAI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_1984),
.A2(n_1920),
.B1(n_1879),
.B2(n_1930),
.C(n_1925),
.Y(n_2035)
);

AOI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1984),
.A2(n_1910),
.B1(n_1875),
.B2(n_1888),
.C(n_1923),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1949),
.B(n_1819),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1996),
.B(n_1865),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1956),
.B(n_1848),
.Y(n_2039)
);

AO21x2_ASAP7_75t_L g2040 ( 
.A1(n_1967),
.A2(n_1821),
.B(n_1937),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1952),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1981),
.A2(n_2022),
.B1(n_2005),
.B2(n_1992),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_2017),
.A2(n_1909),
.B1(n_1919),
.B2(n_1906),
.Y(n_2043)
);

NAND4xp25_ASAP7_75t_L g2044 ( 
.A(n_1986),
.B(n_1795),
.C(n_1915),
.D(n_1823),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1961),
.B(n_1866),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1996),
.B(n_1977),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1956),
.B(n_1960),
.Y(n_2047)
);

OA21x2_ASAP7_75t_L g2048 ( 
.A1(n_1967),
.A2(n_1848),
.B(n_1823),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_2005),
.A2(n_1795),
.B1(n_1919),
.B2(n_1906),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2017),
.A2(n_1882),
.B1(n_1785),
.B2(n_1829),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1992),
.A2(n_1882),
.B1(n_1802),
.B2(n_1851),
.Y(n_2051)
);

OAI221xp5_ASAP7_75t_L g2052 ( 
.A1(n_1999),
.A2(n_1806),
.B1(n_1852),
.B2(n_1810),
.C(n_1846),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_1992),
.A2(n_1829),
.B1(n_1842),
.B2(n_1918),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1977),
.B(n_1850),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1946),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1946),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1985),
.Y(n_2057)
);

NAND4xp25_ASAP7_75t_L g2058 ( 
.A(n_1980),
.B(n_1987),
.C(n_1999),
.D(n_2011),
.Y(n_2058)
);

NOR3xp33_ASAP7_75t_SL g2059 ( 
.A(n_2006),
.B(n_2011),
.C(n_1987),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_2017),
.A2(n_2004),
.B1(n_1989),
.B2(n_1980),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1978),
.B(n_1979),
.Y(n_2061)
);

BUFx2_ASAP7_75t_L g2062 ( 
.A(n_1951),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_2017),
.A2(n_2004),
.B1(n_1989),
.B2(n_2013),
.Y(n_2063)
);

OAI221xp5_ASAP7_75t_L g2064 ( 
.A1(n_2020),
.A2(n_1966),
.B1(n_1994),
.B2(n_2002),
.C(n_1989),
.Y(n_2064)
);

AO21x2_ASAP7_75t_L g2065 ( 
.A1(n_1959),
.A2(n_1968),
.B(n_1965),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1945),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_2004),
.A2(n_2013),
.B1(n_2019),
.B2(n_1995),
.Y(n_2067)
);

INVx4_ASAP7_75t_L g2068 ( 
.A(n_1950),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2020),
.A2(n_1970),
.B(n_1973),
.Y(n_2069)
);

OAI33xp33_ASAP7_75t_L g2070 ( 
.A1(n_1966),
.A2(n_1994),
.A3(n_1997),
.B1(n_1983),
.B2(n_1988),
.B3(n_1972),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1973),
.B(n_2000),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1973),
.B(n_2000),
.Y(n_2072)
);

OAI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_2002),
.A2(n_1997),
.B1(n_2019),
.B2(n_1970),
.C(n_2015),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_1985),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1950),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1950),
.Y(n_2076)
);

NOR3xp33_ASAP7_75t_L g2077 ( 
.A(n_1958),
.B(n_1970),
.C(n_2007),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2004),
.A2(n_2013),
.B1(n_1993),
.B2(n_1995),
.Y(n_2078)
);

OAI211xp5_ASAP7_75t_L g2079 ( 
.A1(n_2007),
.A2(n_2012),
.B(n_2015),
.C(n_1968),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1945),
.Y(n_2080)
);

NAND2xp33_ASAP7_75t_R g2081 ( 
.A(n_1991),
.B(n_1943),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1943),
.B(n_2001),
.Y(n_2082)
);

NAND4xp25_ASAP7_75t_L g2083 ( 
.A(n_1947),
.B(n_1954),
.C(n_1948),
.D(n_1951),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1954),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1943),
.B(n_2001),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_1963),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2004),
.A2(n_2013),
.B1(n_1993),
.B2(n_1995),
.Y(n_2087)
);

OA21x2_ASAP7_75t_L g2088 ( 
.A1(n_1974),
.A2(n_1959),
.B(n_1965),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1964),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1958),
.B(n_2024),
.Y(n_2090)
);

AOI31xp33_ASAP7_75t_L g2091 ( 
.A1(n_1991),
.A2(n_2021),
.A3(n_2012),
.B(n_2024),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1964),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1969),
.Y(n_2093)
);

OAI31xp33_ASAP7_75t_L g2094 ( 
.A1(n_2021),
.A2(n_1959),
.A3(n_1965),
.B(n_1968),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1969),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1971),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2065),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2071),
.B(n_1948),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2071),
.B(n_1998),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_2074),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_2041),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2055),
.B(n_1976),
.Y(n_2102)
);

NAND2x1_ASAP7_75t_L g2103 ( 
.A(n_2068),
.B(n_1998),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2055),
.B(n_1976),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2072),
.B(n_1982),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2056),
.B(n_1976),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2061),
.B(n_1953),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2056),
.B(n_2069),
.Y(n_2108)
);

AND2x4_ASAP7_75t_L g2109 ( 
.A(n_2077),
.B(n_1942),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2065),
.Y(n_2110)
);

BUFx2_ASAP7_75t_L g2111 ( 
.A(n_2062),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2065),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_2062),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2034),
.B(n_1976),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2066),
.B(n_1976),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2082),
.B(n_2085),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2046),
.B(n_1957),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2080),
.B(n_1976),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2080),
.B(n_1976),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2082),
.B(n_1962),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2084),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2084),
.B(n_1955),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2085),
.B(n_2018),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2042),
.A2(n_2013),
.B1(n_1993),
.B2(n_2003),
.Y(n_2124)
);

INVx1_ASAP7_75t_SL g2125 ( 
.A(n_2057),
.Y(n_2125)
);

AND2x4_ASAP7_75t_L g2126 ( 
.A(n_2086),
.B(n_1942),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2079),
.B(n_1955),
.Y(n_2127)
);

INVxp67_ASAP7_75t_SL g2128 ( 
.A(n_2088),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2038),
.B(n_2018),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2089),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2088),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2088),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2089),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2037),
.B(n_1975),
.Y(n_2134)
);

OR2x6_ASAP7_75t_L g2135 ( 
.A(n_2039),
.B(n_2010),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2058),
.B(n_2027),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2047),
.B(n_2037),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2092),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2054),
.B(n_2009),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_2045),
.B(n_2032),
.Y(n_2140)
);

NAND2x1p5_ASAP7_75t_L g2141 ( 
.A(n_2090),
.B(n_2010),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2131),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2128),
.B(n_2088),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2115),
.B(n_2083),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2116),
.B(n_2054),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2131),
.Y(n_2146)
);

INVxp67_ASAP7_75t_SL g2147 ( 
.A(n_2128),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2134),
.B(n_2093),
.Y(n_2148)
);

BUFx2_ASAP7_75t_L g2149 ( 
.A(n_2109),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2116),
.B(n_2094),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2115),
.B(n_2030),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2116),
.B(n_2026),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2134),
.B(n_2093),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2116),
.B(n_2123),
.Y(n_2154)
);

NAND2x1p5_ASAP7_75t_L g2155 ( 
.A(n_2103),
.B(n_2048),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2123),
.B(n_2026),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2131),
.B(n_2132),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2121),
.Y(n_2158)
);

BUFx2_ASAP7_75t_L g2159 ( 
.A(n_2109),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2118),
.B(n_2091),
.Y(n_2160)
);

BUFx3_ASAP7_75t_L g2161 ( 
.A(n_2111),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2132),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2121),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2099),
.B(n_2029),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2099),
.B(n_2029),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2130),
.Y(n_2166)
);

AND2x4_ASAP7_75t_L g2167 ( 
.A(n_2109),
.B(n_2086),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2130),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2108),
.B(n_2095),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2133),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2132),
.B(n_2098),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2109),
.B(n_2068),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2133),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_2100),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2108),
.B(n_2095),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2097),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2118),
.B(n_2096),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2122),
.B(n_2114),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2097),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2098),
.B(n_2040),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_2119),
.B(n_2114),
.Y(n_2181)
);

INVx3_ASAP7_75t_SL g2182 ( 
.A(n_2126),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2138),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_2101),
.Y(n_2184)
);

NAND2x1p5_ASAP7_75t_L g2185 ( 
.A(n_2103),
.B(n_2048),
.Y(n_2185)
);

INVx3_ASAP7_75t_SL g2186 ( 
.A(n_2126),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2120),
.B(n_2040),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2111),
.B(n_2040),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2122),
.B(n_2096),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2117),
.B(n_2075),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2117),
.B(n_2068),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2097),
.Y(n_2192)
);

INVx1_ASAP7_75t_SL g2193 ( 
.A(n_2174),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2152),
.B(n_2145),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2174),
.Y(n_2195)
);

NOR2x1_ASAP7_75t_L g2196 ( 
.A(n_2161),
.B(n_2136),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2166),
.Y(n_2197)
);

INVx2_ASAP7_75t_SL g2198 ( 
.A(n_2161),
.Y(n_2198)
);

INVx2_ASAP7_75t_SL g2199 ( 
.A(n_2161),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2152),
.B(n_2139),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2166),
.Y(n_2201)
);

OR2x2_ASAP7_75t_L g2202 ( 
.A(n_2151),
.B(n_2137),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_2160),
.B(n_2127),
.Y(n_2203)
);

NOR2x1p5_ASAP7_75t_L g2204 ( 
.A(n_2160),
.B(n_2137),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2166),
.Y(n_2205)
);

INVx1_ASAP7_75t_SL g2206 ( 
.A(n_2160),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2151),
.B(n_2102),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2168),
.Y(n_2208)
);

INVxp33_ASAP7_75t_L g2209 ( 
.A(n_2145),
.Y(n_2209)
);

INVxp67_ASAP7_75t_L g2210 ( 
.A(n_2184),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_2184),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_2145),
.B(n_2140),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_2154),
.B(n_2135),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2143),
.Y(n_2214)
);

INVx2_ASAP7_75t_SL g2215 ( 
.A(n_2161),
.Y(n_2215)
);

AND2x2_ASAP7_75t_L g2216 ( 
.A(n_2152),
.B(n_2139),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2168),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2144),
.A2(n_2070),
.B(n_2127),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2168),
.Y(n_2219)
);

AOI21x1_ASAP7_75t_L g2220 ( 
.A1(n_2188),
.A2(n_2113),
.B(n_2110),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2156),
.B(n_2059),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2156),
.B(n_2169),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2170),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2152),
.B(n_2105),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2156),
.B(n_2169),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2143),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2170),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2156),
.B(n_2060),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2175),
.B(n_2129),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2175),
.B(n_2129),
.Y(n_2230)
);

XNOR2xp5_ASAP7_75t_L g2231 ( 
.A(n_2150),
.B(n_2028),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2170),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_2151),
.B(n_2100),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2173),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2173),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2154),
.B(n_2105),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2143),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2173),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2183),
.Y(n_2239)
);

NOR3xp33_ASAP7_75t_L g2240 ( 
.A(n_2149),
.B(n_2044),
.C(n_2064),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2164),
.B(n_2107),
.Y(n_2241)
);

INVxp67_ASAP7_75t_L g2242 ( 
.A(n_2149),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2183),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2202),
.B(n_2193),
.Y(n_2244)
);

NOR2x1_ASAP7_75t_L g2245 ( 
.A(n_2196),
.B(n_2149),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2194),
.B(n_2164),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2218),
.B(n_2158),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2240),
.A2(n_2063),
.B1(n_2078),
.B2(n_2087),
.Y(n_2248)
);

AOI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2231),
.A2(n_2073),
.B1(n_2124),
.B2(n_2043),
.Y(n_2249)
);

OAI32xp33_ASAP7_75t_L g2250 ( 
.A1(n_2206),
.A2(n_2203),
.A3(n_2221),
.B1(n_2209),
.B2(n_2144),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2231),
.A2(n_2050),
.B1(n_2051),
.B2(n_2067),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_2195),
.Y(n_2252)
);

AOI21xp33_ASAP7_75t_SL g2253 ( 
.A1(n_2212),
.A2(n_2186),
.B(n_2182),
.Y(n_2253)
);

INVxp67_ASAP7_75t_SL g2254 ( 
.A(n_2204),
.Y(n_2254)
);

OAI221xp5_ASAP7_75t_L g2255 ( 
.A1(n_2228),
.A2(n_2144),
.B1(n_2155),
.B2(n_2185),
.C(n_2143),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2211),
.Y(n_2256)
);

NAND3xp33_ASAP7_75t_L g2257 ( 
.A(n_2242),
.B(n_2188),
.C(n_2159),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2197),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2202),
.B(n_2181),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2197),
.Y(n_2260)
);

OAI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2233),
.A2(n_2049),
.B(n_2188),
.Y(n_2261)
);

AOI32xp33_ASAP7_75t_L g2262 ( 
.A1(n_2214),
.A2(n_2180),
.A3(n_2187),
.B1(n_2150),
.B2(n_2147),
.Y(n_2262)
);

A2O1A1Ixp33_ASAP7_75t_L g2263 ( 
.A1(n_2214),
.A2(n_2187),
.B(n_2180),
.C(n_2150),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2222),
.B(n_2158),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2201),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2229),
.A2(n_2187),
.B1(n_2180),
.B2(n_2081),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2201),
.Y(n_2267)
);

OAI322xp33_ASAP7_75t_L g2268 ( 
.A1(n_2207),
.A2(n_2181),
.A3(n_2147),
.B1(n_2178),
.B2(n_2102),
.C1(n_2104),
.C2(n_2106),
.Y(n_2268)
);

INVxp67_ASAP7_75t_L g2269 ( 
.A(n_2198),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2205),
.Y(n_2270)
);

OAI21xp5_ASAP7_75t_L g2271 ( 
.A1(n_2210),
.A2(n_2035),
.B(n_2036),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2205),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2194),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2224),
.B(n_2164),
.Y(n_2274)
);

OAI221xp5_ASAP7_75t_L g2275 ( 
.A1(n_2226),
.A2(n_2155),
.B1(n_2185),
.B2(n_2110),
.C(n_2112),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2224),
.Y(n_2276)
);

OR2x2_ASAP7_75t_L g2277 ( 
.A(n_2230),
.B(n_2181),
.Y(n_2277)
);

NAND2x1_ASAP7_75t_L g2278 ( 
.A(n_2213),
.B(n_2159),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2208),
.Y(n_2279)
);

NAND2xp33_ASAP7_75t_L g2280 ( 
.A(n_2198),
.B(n_2155),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_L g2281 ( 
.A(n_2199),
.B(n_2215),
.C(n_2217),
.Y(n_2281)
);

AND2x4_ASAP7_75t_L g2282 ( 
.A(n_2213),
.B(n_2154),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2225),
.B(n_2158),
.Y(n_2283)
);

NOR3xp33_ASAP7_75t_SL g2284 ( 
.A(n_2241),
.B(n_2025),
.C(n_2076),
.Y(n_2284)
);

NAND4xp25_ASAP7_75t_L g2285 ( 
.A(n_2247),
.B(n_2159),
.C(n_2226),
.D(n_2237),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2258),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2260),
.Y(n_2287)
);

INVx1_ASAP7_75t_SL g2288 ( 
.A(n_2244),
.Y(n_2288)
);

OAI221xp5_ASAP7_75t_L g2289 ( 
.A1(n_2261),
.A2(n_2185),
.B1(n_2155),
.B2(n_2110),
.C(n_2112),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_2282),
.B(n_2213),
.Y(n_2290)
);

OAI22xp33_ASAP7_75t_SL g2291 ( 
.A1(n_2247),
.A2(n_2185),
.B1(n_2155),
.B2(n_2112),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2265),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2267),
.Y(n_2293)
);

OAI211xp5_ASAP7_75t_L g2294 ( 
.A1(n_2250),
.A2(n_2215),
.B(n_2199),
.C(n_2237),
.Y(n_2294)
);

OAI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2245),
.A2(n_2150),
.B(n_2220),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2270),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2272),
.Y(n_2297)
);

INVx1_ASAP7_75t_SL g2298 ( 
.A(n_2278),
.Y(n_2298)
);

O2A1O1Ixp33_ASAP7_75t_L g2299 ( 
.A1(n_2271),
.A2(n_2187),
.B(n_2180),
.C(n_2185),
.Y(n_2299)
);

AOI221xp5_ASAP7_75t_L g2300 ( 
.A1(n_2261),
.A2(n_2178),
.B1(n_2157),
.B2(n_2207),
.C(n_2142),
.Y(n_2300)
);

AOI211xp5_ASAP7_75t_SL g2301 ( 
.A1(n_2255),
.A2(n_2252),
.B(n_2254),
.C(n_2269),
.Y(n_2301)
);

AOI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2271),
.A2(n_2048),
.B1(n_2021),
.B2(n_2142),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2279),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2256),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2263),
.A2(n_2106),
.B(n_2104),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2259),
.Y(n_2306)
);

INVx1_ASAP7_75t_SL g2307 ( 
.A(n_2282),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2273),
.Y(n_2308)
);

OAI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2249),
.A2(n_2052),
.B1(n_2220),
.B2(n_2119),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2246),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2264),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2264),
.Y(n_2312)
);

HB1xp67_ASAP7_75t_L g2313 ( 
.A(n_2257),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_2248),
.A2(n_2251),
.B1(n_2266),
.B2(n_2284),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2283),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2283),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2290),
.B(n_2274),
.Y(n_2317)
);

NOR3xp33_ASAP7_75t_SL g2318 ( 
.A(n_2294),
.B(n_2281),
.C(n_2275),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2288),
.B(n_2276),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2310),
.B(n_2200),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2306),
.Y(n_2321)
);

NOR4xp25_ASAP7_75t_SL g2322 ( 
.A(n_2289),
.B(n_2253),
.C(n_2262),
.D(n_2232),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2290),
.B(n_2200),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2290),
.B(n_2310),
.Y(n_2324)
);

NOR2x1_ASAP7_75t_L g2325 ( 
.A(n_2285),
.B(n_2280),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2313),
.B(n_2216),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2307),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2286),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2287),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2292),
.Y(n_2330)
);

NOR3x1_ASAP7_75t_L g2331 ( 
.A(n_2295),
.B(n_2277),
.C(n_2227),
.Y(n_2331)
);

XNOR2xp5_ASAP7_75t_L g2332 ( 
.A(n_2309),
.B(n_2141),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2293),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2296),
.Y(n_2334)
);

OAI21xp5_ASAP7_75t_SL g2335 ( 
.A1(n_2301),
.A2(n_2172),
.B(n_2216),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2298),
.B(n_2268),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2313),
.B(n_2165),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2308),
.B(n_2236),
.Y(n_2338)
);

NOR3xp33_ASAP7_75t_SL g2339 ( 
.A(n_2304),
.B(n_2076),
.C(n_2208),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_2311),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_SL g2341 ( 
.A1(n_2327),
.A2(n_2299),
.B(n_2291),
.Y(n_2341)
);

NOR5xp2_ASAP7_75t_L g2342 ( 
.A(n_2335),
.B(n_2312),
.C(n_2297),
.D(n_2303),
.E(n_2316),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2317),
.B(n_2236),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2324),
.B(n_2312),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2324),
.B(n_2315),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2327),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2319),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2338),
.B(n_2300),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2331),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2318),
.B(n_2309),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2338),
.B(n_2314),
.Y(n_2351)
);

NAND3xp33_ASAP7_75t_L g2352 ( 
.A(n_2322),
.B(n_2302),
.C(n_2305),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2323),
.B(n_2165),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2321),
.Y(n_2354)
);

AOI221x1_ASAP7_75t_L g2355 ( 
.A1(n_2341),
.A2(n_2321),
.B1(n_2336),
.B2(n_2328),
.C(n_2334),
.Y(n_2355)
);

OAI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_2350),
.A2(n_2325),
.B(n_2332),
.Y(n_2356)
);

AOI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2350),
.A2(n_2302),
.B1(n_2332),
.B2(n_2337),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2352),
.A2(n_2326),
.B(n_2340),
.Y(n_2358)
);

OAI211xp5_ASAP7_75t_L g2359 ( 
.A1(n_2349),
.A2(n_2334),
.B(n_2330),
.C(n_2329),
.Y(n_2359)
);

XNOR2x1_ASAP7_75t_L g2360 ( 
.A(n_2349),
.B(n_2328),
.Y(n_2360)
);

OAI211xp5_ASAP7_75t_SL g2361 ( 
.A1(n_2348),
.A2(n_2339),
.B(n_2330),
.C(n_2329),
.Y(n_2361)
);

AOI221xp5_ASAP7_75t_L g2362 ( 
.A1(n_2346),
.A2(n_2351),
.B1(n_2347),
.B2(n_2344),
.C(n_2354),
.Y(n_2362)
);

AOI222xp33_ASAP7_75t_L g2363 ( 
.A1(n_2344),
.A2(n_2333),
.B1(n_2176),
.B2(n_2179),
.C1(n_2192),
.C2(n_2320),
.Y(n_2363)
);

AOI221xp5_ASAP7_75t_L g2364 ( 
.A1(n_2345),
.A2(n_2317),
.B1(n_2323),
.B2(n_2162),
.C(n_2146),
.Y(n_2364)
);

AOI211xp5_ASAP7_75t_L g2365 ( 
.A1(n_2342),
.A2(n_2353),
.B(n_2343),
.C(n_2031),
.Y(n_2365)
);

AOI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2355),
.A2(n_2243),
.B(n_2227),
.Y(n_2366)
);

O2A1O1Ixp33_ASAP7_75t_L g2367 ( 
.A1(n_2356),
.A2(n_2162),
.B(n_2142),
.C(n_2146),
.Y(n_2367)
);

AOI322xp5_ASAP7_75t_L g2368 ( 
.A1(n_2357),
.A2(n_2146),
.A3(n_2162),
.B1(n_2142),
.B2(n_2157),
.C1(n_2179),
.C2(n_2176),
.Y(n_2368)
);

AND2x2_ASAP7_75t_SL g2369 ( 
.A(n_2362),
.B(n_2033),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2360),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_2361),
.A2(n_2162),
.B1(n_2146),
.B2(n_2176),
.Y(n_2371)
);

INVx5_ASAP7_75t_L g2372 ( 
.A(n_2359),
.Y(n_2372)
);

AOI31xp33_ASAP7_75t_L g2373 ( 
.A1(n_2370),
.A2(n_2365),
.A3(n_2358),
.B(n_2364),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2372),
.B(n_2154),
.Y(n_2374)
);

NAND4xp25_ASAP7_75t_L g2375 ( 
.A(n_2366),
.B(n_2363),
.C(n_2172),
.D(n_2167),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2369),
.A2(n_2157),
.B1(n_2243),
.B2(n_2238),
.Y(n_2376)
);

OAI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2372),
.A2(n_2232),
.B(n_2238),
.Y(n_2377)
);

NAND4xp75_ASAP7_75t_L g2378 ( 
.A(n_2368),
.B(n_2157),
.C(n_2235),
.D(n_2234),
.Y(n_2378)
);

AND2x4_ASAP7_75t_L g2379 ( 
.A(n_2371),
.B(n_2191),
.Y(n_2379)
);

AND3x4_ASAP7_75t_L g2380 ( 
.A(n_2367),
.B(n_2172),
.C(n_2167),
.Y(n_2380)
);

NAND4xp25_ASAP7_75t_L g2381 ( 
.A(n_2374),
.B(n_2172),
.C(n_2167),
.D(n_2234),
.Y(n_2381)
);

NAND4xp25_ASAP7_75t_L g2382 ( 
.A(n_2376),
.B(n_2377),
.C(n_2375),
.D(n_2373),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2380),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2378),
.Y(n_2384)
);

OAI211xp5_ASAP7_75t_SL g2385 ( 
.A1(n_2379),
.A2(n_2235),
.B(n_2239),
.C(n_2223),
.Y(n_2385)
);

AOI22xp33_ASAP7_75t_SL g2386 ( 
.A1(n_2374),
.A2(n_2176),
.B1(n_2192),
.B2(n_2179),
.Y(n_2386)
);

OAI222xp33_ASAP7_75t_L g2387 ( 
.A1(n_2376),
.A2(n_2135),
.B1(n_2219),
.B2(n_2192),
.C1(n_2179),
.C2(n_2141),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2382),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_2383),
.A2(n_2171),
.B1(n_2172),
.B2(n_2192),
.Y(n_2389)
);

NAND3xp33_ASAP7_75t_SL g2390 ( 
.A(n_2384),
.B(n_2141),
.C(n_2171),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2385),
.B(n_2163),
.Y(n_2391)
);

OAI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2388),
.A2(n_2387),
.B(n_2381),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2389),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2393),
.Y(n_2394)
);

OR2x2_ASAP7_75t_L g2395 ( 
.A(n_2392),
.B(n_2390),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2394),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2395),
.Y(n_2397)
);

AOI322xp5_ASAP7_75t_SL g2398 ( 
.A1(n_2394),
.A2(n_2391),
.A3(n_2386),
.B1(n_2165),
.B2(n_2171),
.C1(n_2023),
.C2(n_2190),
.Y(n_2398)
);

AOI21xp5_ASAP7_75t_L g2399 ( 
.A1(n_2397),
.A2(n_2171),
.B(n_2163),
.Y(n_2399)
);

OAI21xp5_ASAP7_75t_L g2400 ( 
.A1(n_2396),
.A2(n_2163),
.B(n_2177),
.Y(n_2400)
);

OAI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2399),
.A2(n_2398),
.B(n_2177),
.Y(n_2401)
);

AOI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2400),
.A2(n_2153),
.B(n_2148),
.Y(n_2402)
);

AOI322xp5_ASAP7_75t_L g2403 ( 
.A1(n_2401),
.A2(n_2172),
.A3(n_2023),
.B1(n_2125),
.B2(n_2053),
.C1(n_2153),
.C2(n_2148),
.Y(n_2403)
);

OAI221xp5_ASAP7_75t_R g2404 ( 
.A1(n_2403),
.A2(n_2402),
.B1(n_2182),
.B2(n_2186),
.C(n_2113),
.Y(n_2404)
);

OAI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2404),
.A2(n_2186),
.B1(n_2182),
.B2(n_2189),
.Y(n_2405)
);


endmodule