module fake_jpeg_22425_n_289 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_18),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_67),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_26),
.B1(n_24),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_57),
.B1(n_62),
.B2(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_28),
.B1(n_24),
.B2(n_19),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_61),
.B1(n_79),
.B2(n_0),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_24),
.B1(n_28),
.B2(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_75),
.B1(n_86),
.B2(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

AND2x4_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_29),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_60),
.A2(n_1),
.B(n_2),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_45),
.B1(n_39),
.B2(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_19),
.B1(n_18),
.B2(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_71),
.Y(n_95)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_73),
.Y(n_108)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_23),
.B1(n_33),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_32),
.B1(n_23),
.B2(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_22),
.B1(n_37),
.B2(n_30),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_22),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_41),
.A2(n_38),
.B1(n_30),
.B2(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_42),
.A2(n_27),
.B1(n_31),
.B2(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_13),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_35),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_42),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_42),
.B1(n_35),
.B2(n_31),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_85),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_115),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_31),
.A3(n_29),
.B1(n_21),
.B2(n_5),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_65),
.B(n_79),
.C(n_62),
.D(n_84),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_104),
.B1(n_109),
.B2(n_66),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_11),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_111),
.C(n_56),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_11),
.B1(n_16),
.B2(n_5),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_1),
.C(n_2),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_17),
.B1(n_12),
.B2(n_6),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_73),
.B(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_52),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_118),
.Y(n_150)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g178 ( 
.A(n_123),
.B(n_128),
.C(n_129),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_134),
.B1(n_92),
.B2(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_127),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_68),
.B1(n_74),
.B2(n_70),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_51),
.B1(n_54),
.B2(n_53),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_144),
.B1(n_153),
.B2(n_91),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_80),
.B1(n_53),
.B2(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_82),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_140),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_81),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_143),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_67),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_100),
.A2(n_51),
.B1(n_50),
.B2(n_68),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_154),
.B1(n_115),
.B2(n_117),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_64),
.Y(n_147)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_64),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_97),
.A2(n_84),
.B1(n_71),
.B2(n_16),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_92),
.A2(n_71),
.B1(n_15),
.B2(n_17),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_156),
.A2(n_167),
.B1(n_175),
.B2(n_176),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_122),
.C(n_106),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_179),
.C(n_135),
.Y(n_191)
);

AOI21x1_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_92),
.B(n_96),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_138),
.B1(n_130),
.B2(n_154),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_163),
.Y(n_187)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_166),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_SL g166 ( 
.A(n_127),
.B(n_114),
.C(n_110),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_114),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_177),
.B(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_91),
.B1(n_119),
.B2(n_122),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_14),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_129),
.B(n_119),
.C(n_105),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_105),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_128),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_137),
.B(n_110),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_183),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_124),
.A2(n_118),
.B(n_14),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_177),
.C(n_171),
.Y(n_227)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_208),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_153),
.B(n_132),
.C(n_144),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_209),
.B(n_165),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_142),
.B1(n_147),
.B2(n_125),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_205),
.B1(n_176),
.B2(n_164),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_202),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_177),
.C(n_166),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_130),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_14),
.Y(n_228)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_206),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_145),
.B1(n_126),
.B2(n_141),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_148),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_152),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_207),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

OAI322xp33_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_178),
.A3(n_169),
.B1(n_182),
.B2(n_180),
.C1(n_157),
.C2(n_158),
.Y(n_210)
);

OA21x2_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_211),
.B(n_223),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_178),
.B(n_184),
.C(n_182),
.D(n_165),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_169),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_168),
.B(n_185),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_190),
.B(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_225),
.B1(n_194),
.B2(n_199),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_175),
.B1(n_181),
.B2(n_174),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_195),
.B1(n_207),
.B2(n_193),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_179),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_200),
.B1(n_201),
.B2(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_202),
.C(n_190),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_209),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_186),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_217),
.B1(n_224),
.B2(n_226),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_239),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_199),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_222),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_228),
.B(n_216),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_189),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_211),
.C(n_214),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_187),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_243),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_204),
.C(n_197),
.Y(n_244)
);

XNOR2x2_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.C(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_235),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_224),
.B(n_218),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_237),
.B(n_244),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_238),
.B(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_222),
.B1(n_213),
.B2(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_246),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_232),
.B1(n_241),
.B2(n_243),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_251),
.Y(n_271)
);

AOI31xp67_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_249),
.A3(n_229),
.B(n_245),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_264),
.B(n_254),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_271),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_248),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_268),
.A2(n_272),
.B(n_261),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_270),
.B1(n_263),
.B2(n_236),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_187),
.Y(n_272)
);

AOI21x1_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_260),
.B(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_277),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_266),
.C(n_245),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_281),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_192),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_276),
.B(n_274),
.Y(n_283)
);

AOI321xp33_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_284),
.A3(n_280),
.B1(n_285),
.B2(n_197),
.C(n_208),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_277),
.Y(n_284)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_287),
.B(n_208),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_171),
.Y(n_289)
);


endmodule