module fake_netlist_1_10_n_698 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_698);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_698;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_9), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_37), .Y(n_80) );
INVx4_ASAP7_75t_R g81 ( .A(n_1), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_74), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_21), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_20), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_39), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_72), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_25), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_6), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_40), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_1), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_69), .Y(n_93) );
BUFx2_ASAP7_75t_L g94 ( .A(n_27), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_15), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_57), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_15), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_44), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_26), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_36), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_75), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_71), .Y(n_103) );
NOR2xp67_ASAP7_75t_L g104 ( .A(n_34), .B(n_70), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_49), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_58), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_62), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_66), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_67), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_64), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_46), .Y(n_113) );
CKINVDCx14_ASAP7_75t_R g114 ( .A(n_60), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_22), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_51), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_30), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_28), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_5), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_45), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_23), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_10), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_55), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_56), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_29), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_10), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_94), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_113), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_94), .B(n_0), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_102), .B(n_0), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_113), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_80), .A2(n_35), .B(n_77), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_126), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_79), .B(n_2), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_91), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_98), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_98), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_79), .B(n_2), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_100), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_117), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_125), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_105), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
OR2x2_ASAP7_75t_L g151 ( .A(n_85), .B(n_3), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_106), .Y(n_152) );
INVxp67_ASAP7_75t_L g153 ( .A(n_101), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_107), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_97), .B(n_119), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_107), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_108), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_108), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
XOR2xp5_ASAP7_75t_L g161 ( .A(n_116), .B(n_3), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_111), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_88), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_111), .B(n_4), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_115), .Y(n_165) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_88), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_115), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_120), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_89), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_120), .B(n_4), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_127), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_127), .B(n_114), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_155), .B(n_96), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_169), .B(n_83), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_169), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_136), .B(n_84), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
OAI221xp5_ASAP7_75t_L g180 ( .A1(n_153), .A2(n_110), .B1(n_90), .B2(n_122), .C(n_112), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_145), .B(n_121), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
NOR2xp67_ASAP7_75t_L g183 ( .A(n_160), .B(n_87), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_133), .B(n_90), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_145), .B(n_121), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_136), .B(n_93), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_137), .B(n_139), .Y(n_188) );
NOR2xp67_ASAP7_75t_L g189 ( .A(n_163), .B(n_110), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_137), .A2(n_104), .B(n_99), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_129), .A2(n_112), .B1(n_122), .B2(n_124), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_139), .B(n_118), .Y(n_196) );
NOR2xp33_ASAP7_75t_R g197 ( .A(n_158), .B(n_123), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_166), .B(n_92), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_158), .B(n_86), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_129), .B(n_81), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_130), .A2(n_82), .B1(n_95), .B2(n_109), .Y(n_201) );
NOR3xp33_ASAP7_75t_L g202 ( .A(n_170), .B(n_6), .C(n_7), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
NOR2x1_ASAP7_75t_L g204 ( .A(n_140), .B(n_7), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_140), .B(n_8), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_142), .B(n_9), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_142), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_165), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_143), .B(n_11), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_143), .B(n_12), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_144), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_148), .A2(n_14), .B(n_16), .C(n_17), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_165), .B(n_48), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
AND2x4_ASAP7_75t_SL g217 ( .A(n_148), .B(n_14), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_150), .B(n_50), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_164), .B(n_17), .C(n_18), .Y(n_219) );
INVx8_ASAP7_75t_L g220 ( .A(n_149), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_150), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
BUFx12f_ASAP7_75t_L g223 ( .A(n_151), .Y(n_223) );
OAI21xp33_ASAP7_75t_L g224 ( .A1(n_154), .A2(n_18), .B(n_19), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_151), .A2(n_24), .B(n_31), .C(n_32), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_154), .B(n_33), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_156), .B(n_38), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_149), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_161), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_221), .B(n_168), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_199), .B(n_168), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_226), .B(n_156), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_171), .A2(n_159), .B1(n_157), .B2(n_134), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_175), .B(n_157), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_194), .B(n_141), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_223), .Y(n_236) );
AND3x1_ASAP7_75t_SL g237 ( .A(n_180), .B(n_159), .C(n_134), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_174), .B(n_167), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_200), .B(n_141), .Y(n_239) );
NOR2xp33_ASAP7_75t_R g240 ( .A(n_177), .B(n_41), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_212), .A2(n_167), .B1(n_162), .B2(n_152), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_191), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_188), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_195), .A2(n_167), .B1(n_162), .B2(n_152), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_200), .B(n_162), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_183), .B(n_152), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_197), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_199), .B(n_135), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_182), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_178), .B(n_135), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_190), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_200), .B(n_147), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_191), .Y(n_253) );
NAND2x1p5_ASAP7_75t_L g254 ( .A(n_204), .B(n_135), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_177), .B(n_147), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_176), .B(n_147), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_193), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_203), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_217), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_189), .B(n_146), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_173), .B(n_146), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_186), .B(n_146), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_223), .B(n_138), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_184), .B(n_138), .Y(n_266) );
CKINVDCx8_ASAP7_75t_R g267 ( .A(n_229), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_217), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_198), .A2(n_138), .B1(n_131), .B2(n_128), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_197), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_196), .B(n_131), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_229), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_205), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_206), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_201), .A2(n_131), .B1(n_128), .B2(n_149), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_220), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_192), .B(n_128), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_181), .B(n_149), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_225), .B(n_202), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_181), .B(n_149), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_185), .Y(n_282) );
BUFx4f_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_207), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_227), .A2(n_132), .B(n_43), .C(n_47), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_185), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_219), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_220), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_227), .B(n_132), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_214), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_214), .Y(n_291) );
BUFx4f_ASAP7_75t_L g292 ( .A(n_220), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_208), .B(n_132), .Y(n_293) );
AND2x2_ASAP7_75t_SL g294 ( .A(n_224), .B(n_132), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_290), .A2(n_218), .B1(n_215), .B2(n_228), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_235), .B(n_228), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_243), .B(n_218), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_291), .A2(n_215), .B1(n_222), .B2(n_210), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_230), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_276), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_267), .Y(n_301) );
BUFx2_ASAP7_75t_SL g302 ( .A(n_236), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_257), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_232), .A2(n_222), .B(n_210), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_259), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_239), .B(n_213), .Y(n_306) );
INVx3_ASAP7_75t_SL g307 ( .A(n_236), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_289), .A2(n_187), .B(n_179), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_283), .B(n_213), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_255), .B(n_187), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_259), .B(n_213), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_272), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_268), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_179), .B(n_172), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_268), .B(n_42), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_239), .B(n_52), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_284), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_249), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_276), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_258), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_274), .B(n_213), .Y(n_324) );
OAI321xp33_ASAP7_75t_L g325 ( .A1(n_280), .A2(n_172), .A3(n_54), .B1(n_59), .B2(n_61), .C(n_63), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_241), .A2(n_53), .B1(n_65), .B2(n_68), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_285), .A2(n_73), .B(n_76), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_232), .A2(n_78), .B(n_238), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_256), .A2(n_248), .B(n_262), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_251), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_250), .A2(n_263), .B(n_273), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_SL g332 ( .A1(n_287), .A2(n_278), .B(n_271), .C(n_279), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_260), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_276), .Y(n_334) );
INVx3_ASAP7_75t_SL g335 ( .A(n_245), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_264), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_266), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_261), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_245), .B(n_252), .Y(n_339) );
OR2x6_ASAP7_75t_L g340 ( .A(n_247), .B(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_274), .B(n_256), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
NOR2x1_ASAP7_75t_SL g343 ( .A(n_277), .B(n_288), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_264), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_241), .A2(n_233), .B1(n_231), .B2(n_262), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_261), .B(n_265), .Y(n_346) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_270), .B(n_292), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_341), .B(n_231), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_300), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_299), .B(n_244), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_339), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_308), .A2(n_254), .B(n_281), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_303), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_327), .A2(n_254), .B(n_269), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_333), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_329), .B(n_248), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_300), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_339), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_303), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_335), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
INVx2_ASAP7_75t_SL g366 ( .A(n_300), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_300), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_313), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_323), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g372 ( .A1(n_345), .A2(n_294), .B(n_234), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_337), .B(n_246), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_321), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_321), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_336), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_318), .B(n_286), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_353), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_348), .B(n_318), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_348), .B(n_318), .Y(n_383) );
AND2x4_ASAP7_75t_SL g384 ( .A(n_380), .B(n_317), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_348), .B(n_297), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_380), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_362), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_355), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_355), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_356), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g393 ( .A1(n_350), .A2(n_315), .B1(n_338), .B2(n_317), .C1(n_347), .C2(n_319), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_380), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_353), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_358), .B(n_344), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_365), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_356), .B(n_340), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_349), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_372), .A2(n_316), .B(n_325), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_340), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_357), .B(n_317), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_365), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_349), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_349), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_382), .A2(n_358), .B1(n_350), .B2(n_351), .Y(n_409) );
AOI21x1_ASAP7_75t_L g410 ( .A1(n_402), .A2(n_372), .B(n_354), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_389), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_389), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_393), .A2(n_358), .B1(n_350), .B2(n_351), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_387), .B(n_349), .Y(n_414) );
AOI31xp33_ASAP7_75t_L g415 ( .A1(n_393), .A2(n_360), .A3(n_270), .B(n_301), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_382), .A2(n_357), .B1(n_360), .B2(n_340), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_381), .B(n_357), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_382), .A2(n_351), .B1(n_361), .B2(n_346), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_385), .A2(n_361), .B1(n_379), .B2(n_275), .C(n_364), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_381), .B(n_369), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_397), .B(n_369), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_383), .A2(n_347), .B1(n_379), .B2(n_373), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_397), .B(n_369), .Y(n_425) );
OAI31xp33_ASAP7_75t_SL g426 ( .A1(n_404), .A2(n_354), .A3(n_326), .B(n_364), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_404), .A2(n_370), .B1(n_378), .B2(n_377), .Y(n_429) );
NAND4xp25_ASAP7_75t_L g430 ( .A(n_400), .B(n_373), .C(n_379), .D(n_306), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_394), .B(n_375), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_401), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_394), .B(n_375), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_401), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_396), .B(n_375), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_400), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_384), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_396), .B(n_375), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_396), .B(n_365), .Y(n_440) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_387), .A2(n_354), .B(n_332), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_401), .Y(n_442) );
NOR3x1_ASAP7_75t_L g443 ( .A(n_430), .B(n_395), .C(n_386), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_417), .B(n_386), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_417), .B(n_395), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_415), .B(n_385), .C(n_373), .Y(n_447) );
OAI21xp33_ASAP7_75t_SL g448 ( .A1(n_430), .A2(n_392), .B(n_403), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_417), .B(n_387), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_419), .A2(n_383), .B(n_388), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_412), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_420), .B(n_403), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_420), .B(n_399), .Y(n_455) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_426), .B(n_384), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_420), .B(n_399), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_442), .B(n_407), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_442), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_423), .B(n_398), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_423), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_422), .B(n_388), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_427), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_428), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_423), .B(n_425), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_435), .B(n_388), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_406), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_431), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_442), .B(n_407), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_437), .B(n_406), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_434), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_437), .B(n_406), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_431), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_433), .B(n_405), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_433), .B(n_436), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_433), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_434), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_436), .B(n_398), .Y(n_487) );
AOI32xp33_ASAP7_75t_L g488 ( .A1(n_416), .A2(n_384), .A3(n_404), .B1(n_305), .B2(n_314), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_439), .B(n_392), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_447), .A2(n_415), .B1(n_416), .B2(n_413), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_445), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_450), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_470), .B(n_429), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_483), .B(n_440), .Y(n_496) );
NOR3xp33_ASAP7_75t_SL g497 ( .A(n_448), .B(n_438), .C(n_419), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_473), .B(n_440), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_452), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_469), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_461), .B(n_440), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_473), .B(n_414), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_462), .B(n_414), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_463), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_454), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_453), .B(n_429), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_487), .B(n_409), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_463), .B(n_414), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_469), .B(n_414), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_460), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_464), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_444), .B(n_409), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_466), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_446), .B(n_432), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_467), .B(n_398), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_468), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_459), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_474), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_447), .B(n_404), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_458), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_449), .B(n_432), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_486), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_475), .B(n_414), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_486), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_479), .B(n_424), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_465), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_465), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_471), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_471), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_458), .B(n_405), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_477), .B(n_432), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_481), .B(n_441), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_449), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_484), .B(n_441), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_455), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_479), .B(n_418), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_478), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_485), .B(n_441), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_457), .B(n_405), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_491), .B(n_408), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_476), .B(n_399), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_480), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_456), .A2(n_237), .B1(n_305), .B2(n_306), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_491), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_489), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_490), .B(n_426), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_488), .B(n_408), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_472), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_482), .B(n_441), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_500), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_535), .B(n_476), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_510), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_516), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_514), .B(n_456), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_497), .B(n_451), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_496), .B(n_451), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_544), .B(n_443), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_533), .B(n_410), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_537), .B(n_410), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_542), .B(n_408), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_501), .B(n_407), .Y(n_562) );
OA21x2_ASAP7_75t_L g563 ( .A1(n_546), .A2(n_352), .B(n_328), .Y(n_563) );
OR2x6_ASAP7_75t_L g564 ( .A(n_530), .B(n_366), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_516), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_518), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_518), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_548), .B(n_402), .Y(n_568) );
NAND2xp33_ASAP7_75t_L g569 ( .A(n_492), .B(n_240), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_517), .B(n_376), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g571 ( .A1(n_519), .A2(n_294), .B(n_240), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_493), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_519), .B(n_376), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_494), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_545), .B(n_402), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_499), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_541), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_526), .B(n_402), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_504), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_528), .B(n_402), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_529), .B(n_378), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_521), .B(n_369), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_505), .B(n_511), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_513), .B(n_378), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_527), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_507), .B(n_377), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_525), .B(n_536), .C(n_522), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_525), .B(n_377), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_503), .B(n_359), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_522), .B(n_307), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_523), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_498), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_539), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_498), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_495), .B(n_370), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_503), .B(n_502), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_503), .B(n_359), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_509), .Y(n_602) );
NAND4xp75_ASAP7_75t_L g603 ( .A(n_556), .B(n_547), .C(n_536), .D(n_543), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_589), .A2(n_512), .B1(n_540), .B2(n_524), .C(n_534), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_597), .B(n_534), .Y(n_605) );
AO221x1_ASAP7_75t_L g606 ( .A1(n_596), .A2(n_520), .B1(n_547), .B2(n_506), .C(n_540), .Y(n_606) );
OAI21xp33_ASAP7_75t_SL g607 ( .A1(n_597), .A2(n_520), .B(n_509), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_600), .B(n_520), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_584), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_573), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_556), .B(n_515), .C(n_549), .Y(n_611) );
BUFx4f_ASAP7_75t_SL g612 ( .A(n_593), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_575), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_577), .Y(n_614) );
BUFx3_ASAP7_75t_L g615 ( .A(n_551), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_569), .A2(n_502), .B1(n_534), .B2(n_508), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_569), .B(n_324), .C(n_370), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_593), .A2(n_508), .B(n_532), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_550), .B(n_538), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_550), .A2(n_538), .B(n_532), .Y(n_620) );
AOI21xp5_ASAP7_75t_SL g621 ( .A1(n_578), .A2(n_343), .B(n_312), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_557), .A2(n_307), .B1(n_312), .B2(n_363), .Y(n_622) );
NOR4xp25_ASAP7_75t_L g623 ( .A(n_558), .B(n_332), .C(n_363), .D(n_371), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_594), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_591), .B(n_324), .C(n_295), .D(n_298), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_578), .B(n_359), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_598), .B(n_367), .Y(n_627) );
AOI221x1_ASAP7_75t_L g628 ( .A1(n_571), .A2(n_359), .B1(n_367), .B2(n_363), .C(n_368), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_574), .A2(n_237), .B1(n_371), .B2(n_368), .Y(n_629) );
OA211x2_ASAP7_75t_L g630 ( .A1(n_570), .A2(n_295), .B(n_298), .C(n_310), .Y(n_630) );
INVxp67_ASAP7_75t_SL g631 ( .A(n_572), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_583), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_595), .B(n_367), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_590), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g635 ( .A(n_570), .B(n_588), .C(n_599), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_586), .B(n_367), .C(n_359), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_602), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_552), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_574), .A2(n_367), .B1(n_374), .B2(n_366), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_587), .B(n_352), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_611), .B(n_560), .C(n_559), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_607), .A2(n_585), .B(n_582), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_615), .B(n_555), .Y(n_643) );
O2A1O1Ixp5_ASAP7_75t_L g644 ( .A1(n_618), .A2(n_561), .B(n_553), .C(n_566), .Y(n_644) );
XOR2xp5_ASAP7_75t_L g645 ( .A(n_603), .B(n_562), .Y(n_645) );
XNOR2xp5_ASAP7_75t_L g646 ( .A(n_608), .B(n_601), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_604), .A2(n_567), .B(n_592), .C(n_554), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_634), .Y(n_648) );
AOI311xp33_ASAP7_75t_L g649 ( .A1(n_611), .A2(n_568), .A3(n_579), .B(n_581), .C(n_576), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_610), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_635), .A2(n_565), .B1(n_554), .B2(n_580), .C(n_572), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_635), .A2(n_565), .A3(n_580), .B1(n_563), .B2(n_564), .C1(n_374), .C2(n_366), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_609), .A2(n_304), .B1(n_374), .B2(n_322), .C(n_296), .Y(n_653) );
INVx2_ASAP7_75t_SL g654 ( .A(n_612), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_624), .B(n_563), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_616), .A2(n_564), .B1(n_563), .B2(n_312), .Y(n_656) );
OAI33xp33_ASAP7_75t_L g657 ( .A1(n_619), .A2(n_234), .A3(n_564), .B1(n_282), .B2(n_344), .B3(n_253), .Y(n_657) );
AOI221xp5_ASAP7_75t_SL g658 ( .A1(n_620), .A2(n_321), .B1(n_342), .B2(n_334), .C(n_322), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_632), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_622), .A2(n_342), .B(n_334), .C(n_321), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_606), .A2(n_342), .B1(n_334), .B2(n_352), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_637), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_630), .A2(n_334), .B1(n_342), .B2(n_309), .Y(n_663) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_661), .B(n_629), .C(n_617), .D(n_628), .Y(n_664) );
NOR2x1p5_ASAP7_75t_L g665 ( .A(n_643), .B(n_605), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_642), .A2(n_622), .B(n_623), .C(n_617), .Y(n_666) );
NOR2x1_ASAP7_75t_L g667 ( .A(n_647), .B(n_621), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_651), .B(n_614), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_644), .B(n_636), .C(n_638), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_650), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_659), .B(n_631), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_648), .B(n_613), .Y(n_672) );
NOR4xp75_ASAP7_75t_L g673 ( .A(n_654), .B(n_626), .C(n_640), .D(n_627), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_645), .A2(n_633), .B1(n_631), .B2(n_639), .Y(n_674) );
NOR2xp67_ASAP7_75t_L g675 ( .A(n_641), .B(n_625), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_642), .B(n_309), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_662), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_675), .B(n_649), .C(n_652), .Y(n_678) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_671), .A2(n_655), .B(n_656), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_667), .A2(n_656), .B1(n_657), .B2(n_646), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_672), .Y(n_681) );
NOR2xp67_ASAP7_75t_L g682 ( .A(n_669), .B(n_663), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_670), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_665), .A2(n_660), .B1(n_653), .B2(n_658), .Y(n_684) );
BUFx2_ASAP7_75t_L g685 ( .A(n_677), .Y(n_685) );
NAND5xp2_ASAP7_75t_L g686 ( .A(n_680), .B(n_666), .C(n_674), .D(n_676), .E(n_668), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_678), .B(n_664), .C(n_676), .Y(n_687) );
XOR2x2_ASAP7_75t_L g688 ( .A(n_682), .B(n_673), .Y(n_688) );
NOR2xp67_ASAP7_75t_SL g689 ( .A(n_685), .B(n_288), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_684), .A2(n_242), .B(n_283), .C(n_292), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_690), .B(n_684), .C(n_679), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_687), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_686), .A2(n_288), .B1(n_681), .B2(n_683), .C(n_689), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g694 ( .A1(n_692), .A2(n_688), .B1(n_691), .B2(n_693), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_692), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_695), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_694), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_697), .B(n_696), .Y(n_698) );
endmodule