module fake_jpeg_14985_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

HB1xp67_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_15),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_14),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

BUFx24_ASAP7_75t_SL g18 ( 
.A(n_16),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_12),
.B(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_21),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_14),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.C(n_25),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_9),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_9),
.B(n_7),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_21),
.B(n_0),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.C(n_3),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_24),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.C(n_31),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AO221x1_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.B(n_4),
.Y(n_37)
);


endmodule