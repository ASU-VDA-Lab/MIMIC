module real_jpeg_29754_n_12 (n_5, n_4, n_8, n_0, n_274, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_274;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g62 ( 
.A(n_0),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_1),
.Y(n_101)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_4),
.A2(n_20),
.B1(n_23),
.B2(n_27),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_4),
.A2(n_27),
.B1(n_60),
.B2(n_61),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_4),
.A2(n_27),
.B1(n_39),
.B2(n_41),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_20),
.B1(n_23),
.B2(n_49),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_6),
.A2(n_39),
.B1(n_41),
.B2(n_49),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_20),
.B1(n_23),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_35),
.B1(n_39),
.B2(n_41),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_7),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_208)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_10),
.A2(n_20),
.B1(n_23),
.B2(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_11),
.A2(n_20),
.B1(n_23),
.B2(n_30),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_20),
.B(n_22),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_11),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_30),
.B1(n_39),
.B2(n_41),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_11),
.B(n_19),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_11),
.A2(n_39),
.B(n_148),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_57),
.B(n_61),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_11),
.B(n_38),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_79),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_78),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_64),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_16),
.B(n_64),
.Y(n_78)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_16),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_33),
.CI(n_45),
.CON(n_16),
.SN(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_24),
.B(n_28),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_18),
.A2(n_28),
.B(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_19),
.A2(n_29),
.B1(n_31),
.B2(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_19),
.B(n_31),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

INVx5_ASAP7_75t_SL g23 ( 
.A(n_20),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_20),
.A2(n_30),
.B(n_40),
.C(n_147),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_21),
.A2(n_26),
.B(n_30),
.C(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_29),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_30),
.A2(n_39),
.B(n_58),
.C(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_30),
.B(n_103),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_30),
.B(n_59),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_38),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_37),
.B(n_90),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_38),
.A2(n_51),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_44),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_52),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_67),
.B1(n_87),
.B2(n_92),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_46),
.B(n_92),
.C(n_93),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_46),
.A2(n_67),
.B1(n_107),
.B2(n_129),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_46),
.B(n_129),
.C(n_224),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_52),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_52),
.A2(n_71),
.B1(n_74),
.B2(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_63),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_111),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_55),
.A2(n_59),
.B1(n_111),
.B2(n_117),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_55),
.A2(n_59),
.B1(n_63),
.B2(n_229),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_59),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_60),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_100),
.Y(n_99)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_72),
.C(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_130),
.Y(n_264)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.C(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_107),
.C(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_72),
.A2(n_130),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_72),
.A2(n_130),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_73),
.B(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_74),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_89),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_255),
.A3(n_265),
.B1(n_270),
.B2(n_271),
.C(n_274),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_237),
.B(n_254),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_218),
.B(n_236),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_140),
.B(n_201),
.C(n_217),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_126),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_84),
.B(n_126),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_104),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_85),
.B(n_105),
.C(n_113),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_93),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_135),
.C(n_138),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_87),
.A2(n_92),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_87),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_87),
.B(n_243),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_97),
.A2(n_133),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_97),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_97),
.B(n_185),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_162),
.C(n_174),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_123),
.B(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_99),
.B(n_100),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_99),
.A2(n_103),
.B1(n_122),
.B2(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_112),
.B2(n_113),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_107),
.A2(n_114),
.B1(n_115),
.B2(n_129),
.Y(n_192)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_114),
.A2(n_115),
.B1(n_169),
.B2(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_114),
.B(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_129),
.C(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_115),
.B(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B(n_119),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.C(n_134),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_127),
.B(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_130),
.B(n_211),
.C(n_213),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_132),
.B(n_134),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_135),
.B(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_200),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_195),
.B(n_199),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_165),
.B(n_194),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_153),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_152),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_162),
.C(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_156),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_162),
.A2(n_164),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_207),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_189),
.B(n_193),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_176),
.B(n_188),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_171),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_169),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B(n_187),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_184),
.B(n_186),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_215),
.B2(n_216),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_210),
.C(n_216),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_219),
.B(n_220),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_235),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_227),
.C(n_235),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_231),
.B1(n_232),
.B2(n_234),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_232),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_246),
.B(n_248),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_252),
.B2(n_253),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_245),
.C(n_253),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_257),
.C(n_261),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_257),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_261),
.A2(n_262),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);


endmodule