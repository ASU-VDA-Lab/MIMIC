module fake_jpeg_6974_n_40 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_40);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_8),
.B1(n_18),
.B2(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_9),
.B1(n_14),
.B2(n_4),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

A2O1A1O1Ixp25_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_20),
.B(n_1),
.C(n_0),
.D(n_22),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_36),
.A3(n_21),
.B1(n_26),
.B2(n_11),
.C1(n_12),
.C2(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_34),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_35),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_5),
.B(n_7),
.Y(n_40)
);


endmodule