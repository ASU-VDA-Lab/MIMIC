module fake_jpeg_31607_n_77 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_9),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AO22x1_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_13),
.B1(n_23),
.B2(n_22),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_48),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_27),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_26),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_3),
.Y(n_60)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_32),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_18),
.C(n_17),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_4),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_2),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_59),
.C(n_4),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_48),
.B(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_61),
.B1(n_5),
.B2(n_11),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_24),
.B1(n_15),
.B2(n_6),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_65),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_62),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_53),
.Y(n_73)
);

OAI321xp33_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_54),
.A3(n_68),
.B1(n_71),
.B2(n_63),
.C(n_16),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_69),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_58),
.Y(n_77)
);


endmodule