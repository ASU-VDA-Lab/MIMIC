module real_jpeg_16906_n_23 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_23);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_23;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_51;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_0),
.B(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_0),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_1),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_10),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI222xp33_ASAP7_75t_L g23 ( 
.A1(n_3),
.A2(n_24),
.B1(n_63),
.B2(n_66),
.C1(n_83),
.C2(n_86),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_5),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_6),
.C(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_32),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_7),
.B(n_15),
.C(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_9),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_47),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_9),
.B(n_14),
.C(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_13),
.B(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_16),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_25),
.B1(n_61),
.B2(n_62),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_18),
.A2(n_61),
.B1(n_67),
.B2(n_82),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_19),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_58),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_43),
.C(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

AOI31xp33_ASAP7_75t_L g54 ( 
.A1(n_22),
.A2(n_35),
.A3(n_51),
.B(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_60),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_57),
.B(n_59),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B(n_56),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_50),
.B(n_53),
.C(n_54),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B(n_49),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_75),
.C(n_79),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_48),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_77),
.C(n_78),
.Y(n_76)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_55),
.C(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_71),
.C(n_80),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_81),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);


endmodule