module fake_jpeg_19753_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_41),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_47),
.B1(n_54),
.B2(n_22),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_47)
);

NAND2xp67_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_18),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_21),
.B1(n_23),
.B2(n_32),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_42),
.A3(n_16),
.B1(n_33),
.B2(n_28),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_28),
.B1(n_33),
.B2(n_19),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_69),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_22),
.B1(n_19),
.B2(n_25),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_67),
.B1(n_83),
.B2(n_62),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_53),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_85),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_82),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_27),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_84),
.B(n_37),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_22),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_38),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_59),
.B1(n_18),
.B2(n_30),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_106),
.B1(n_108),
.B2(n_113),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_59),
.C(n_34),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_117),
.C(n_34),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_80),
.B1(n_79),
.B2(n_89),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_84),
.B1(n_71),
.B2(n_72),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_30),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_68),
.B1(n_64),
.B2(n_34),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_75),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_18),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_90),
.B(n_76),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_144),
.B1(n_97),
.B2(n_88),
.Y(n_167)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_130),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_30),
.B(n_18),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_127),
.A2(n_31),
.B(n_26),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_128),
.B(n_134),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_86),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_132),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_91),
.B1(n_60),
.B2(n_77),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_138),
.B1(n_115),
.B2(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_70),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_60),
.B1(n_68),
.B2(n_64),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

AO21x2_ASAP7_75t_L g144 ( 
.A1(n_96),
.A2(n_36),
.B(n_35),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_36),
.B1(n_35),
.B2(n_12),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_98),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_36),
.B1(n_35),
.B2(n_12),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_94),
.A2(n_118),
.B1(n_117),
.B2(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_112),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_112),
.B1(n_109),
.B2(n_114),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_143),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_114),
.B1(n_118),
.B2(n_103),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_146),
.A2(n_118),
.B1(n_122),
.B2(n_100),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_122),
.B1(n_121),
.B2(n_97),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_172),
.B1(n_176),
.B2(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_121),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_171),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_167),
.B(n_170),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_97),
.B1(n_88),
.B2(n_15),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_170),
.A2(n_173),
.B1(n_164),
.B2(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_24),
.B1(n_17),
.B2(n_30),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_30),
.B1(n_26),
.B2(n_14),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_175),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_124),
.B1(n_123),
.B2(n_130),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_123),
.A2(n_24),
.B1(n_17),
.B2(n_31),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_180),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_123),
.A2(n_24),
.B1(n_17),
.B2(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_140),
.A2(n_24),
.B1(n_26),
.B2(n_13),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_149),
.C(n_141),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_187),
.C(n_201),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_136),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_206),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_159),
.C(n_152),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_189),
.A2(n_191),
.B1(n_194),
.B2(n_198),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_167),
.B1(n_152),
.B2(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_142),
.B1(n_144),
.B2(n_135),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_135),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_144),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_124),
.B1(n_126),
.B2(n_2),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_205),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_0),
.C(n_1),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_4),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_0),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_212),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_168),
.B(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_157),
.B(n_3),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_160),
.B(n_3),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_181),
.B(n_4),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_169),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_171),
.CI(n_180),
.CON(n_221),
.SN(n_221)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_226),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_179),
.B(n_166),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_166),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_184),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_177),
.B(n_182),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_163),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_204),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_4),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_211),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_215),
.B1(n_194),
.B2(n_199),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_244),
.A2(n_239),
.B1(n_202),
.B2(n_222),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_248),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_189),
.B1(n_188),
.B2(n_202),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_227),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_253),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_210),
.C(n_200),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_221),
.C(n_227),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_219),
.B(n_210),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_255),
.A2(n_238),
.B1(n_231),
.B2(n_236),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_205),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_212),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_261),
.Y(n_263)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_203),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_239),
.B1(n_225),
.B2(n_220),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_276),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_268),
.C(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_270),
.B1(n_274),
.B2(n_235),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_244),
.A2(n_260),
.B1(n_250),
.B2(n_251),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_221),
.C(n_240),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_250),
.A2(n_257),
.B1(n_255),
.B2(n_218),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_254),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_237),
.C(n_236),
.Y(n_284)
);

XOR2x2_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_218),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_233),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_240),
.B(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_285),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_234),
.Y(n_283)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_287),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_230),
.B1(n_248),
.B2(n_229),
.Y(n_286)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_4),
.C(n_5),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_269),
.B(n_5),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_290),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_5),
.C(n_6),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_5),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_7),
.C(n_8),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_272),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_267),
.B1(n_278),
.B2(n_263),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_7),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_263),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_292),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_281),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_281),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_271),
.C(n_275),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_310),
.A2(n_313),
.B(n_8),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_271),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_314),
.B(n_302),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_294),
.B(n_8),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_303),
.B(n_295),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_316),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_305),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_306),
.C(n_310),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_8),
.B(n_9),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_323),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_320),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_319),
.B(n_322),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_10),
.B(n_11),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_10),
.B1(n_11),
.B2(n_305),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_10),
.B(n_11),
.Y(n_329)
);


endmodule