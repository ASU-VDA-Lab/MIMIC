module fake_jpeg_16968_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_41),
.B1(n_44),
.B2(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_47),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_2),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_22),
.B(n_23),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_13),
.B(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_2),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_44),
.B1(n_43),
.B2(n_39),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_67),
.B1(n_53),
.B2(n_3),
.Y(n_76)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_73),
.B1(n_70),
.B2(n_5),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_19),
.B1(n_34),
.B2(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_6),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_26),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_56),
.B1(n_57),
.B2(n_21),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_87),
.B(n_68),
.C(n_7),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_58),
.B1(n_10),
.B2(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_8),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_8),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_98),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_95),
.B1(n_83),
.B2(n_93),
.Y(n_102)
);

OAI321xp33_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_103),
.A3(n_99),
.B1(n_82),
.B2(n_88),
.C(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_91),
.C(n_89),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_101),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_9),
.CI(n_25),
.CON(n_106),
.SN(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_27),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_38),
.Y(n_110)
);


endmodule