module fake_ariane_74_n_863 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_863);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_863;

wire n_295;
wire n_556;
wire n_356;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_600;
wire n_433;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_590;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_429;
wire n_654;
wire n_365;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_571;
wire n_680;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_650;
wire n_258;
wire n_364;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_98),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_105),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_91),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_108),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_23),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_10),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_21),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_14),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_96),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_57),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_128),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_106),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_119),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_177),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_79),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_16),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_9),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_83),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_84),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_82),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_10),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_31),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_114),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_143),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_3),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_169),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_53),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_168),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_80),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_111),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_1),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_116),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_127),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_170),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_155),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_94),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_42),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_134),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_42),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_176),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_99),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_156),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_120),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_27),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_181),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_130),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_121),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_124),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_72),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_25),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_193),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_126),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_47),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_64),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_178),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_102),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_44),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_54),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_208),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_88),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_118),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_81),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_152),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_74),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_22),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_203),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_112),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_72),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_140),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_189),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_149),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_198),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_199),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_97),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_74),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_44),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_192),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_207),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_179),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_184),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_150),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_138),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_71),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_142),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_147),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_50),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_185),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_48),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_46),
.Y(n_320)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_63),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_75),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_204),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_161),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_110),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_202),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_117),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_113),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_43),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_62),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_78),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_194),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_28),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_58),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_195),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_0),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_0),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_85),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_210),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_210),
.Y(n_344)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_235),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_302),
.B(n_1),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_216),
.B(n_2),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_216),
.B(n_3),
.Y(n_348)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_235),
.Y(n_350)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_210),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_4),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_239),
.B(n_5),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_295),
.B(n_5),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_6),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_210),
.Y(n_356)
);

BUFx8_ASAP7_75t_SL g357 ( 
.A(n_288),
.Y(n_357)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_236),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_264),
.B(n_8),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_218),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_213),
.B(n_8),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_217),
.B(n_9),
.Y(n_362)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_236),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_218),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_218),
.Y(n_365)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_236),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_222),
.B(n_11),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_218),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_86),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_247),
.Y(n_371)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_211),
.B(n_87),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_264),
.B(n_12),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_282),
.B(n_12),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g375 ( 
.A(n_251),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_220),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_247),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_247),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_251),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_247),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_229),
.B(n_13),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_234),
.B(n_14),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_15),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_259),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_265),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_259),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_238),
.B(n_16),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_259),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_294),
.B(n_17),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_240),
.B(n_18),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_265),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_241),
.B(n_18),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_259),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_282),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_244),
.B(n_19),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_322),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_249),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_248),
.B(n_20),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_223),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_20),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_253),
.B(n_21),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_294),
.B(n_22),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_256),
.B(n_24),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_260),
.B(n_25),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_277),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_320),
.B(n_26),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_263),
.B(n_27),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_331),
.B(n_29),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_322),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_215),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_299),
.B(n_30),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_297),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_219),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_297),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_268),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_299),
.B(n_228),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_225),
.B(n_257),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_286),
.B(n_32),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_211),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_331),
.B(n_246),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_281),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_305),
.Y(n_427)
);

BUFx8_ASAP7_75t_L g428 ( 
.A(n_246),
.Y(n_428)
);

NAND2x1_ASAP7_75t_L g429 ( 
.A(n_269),
.B(n_274),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_230),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_231),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_232),
.B(n_33),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_289),
.B(n_34),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_237),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_274),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_243),
.B(n_35),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_280),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_280),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_291),
.B(n_293),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_250),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_254),
.B(n_36),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_315),
.B(n_318),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_290),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_312),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_242),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_284),
.B(n_37),
.Y(n_446)
);

AO22x2_ASAP7_75t_L g447 ( 
.A1(n_374),
.A2(n_323),
.B1(n_330),
.B2(n_307),
.Y(n_447)
);

AO22x2_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_334),
.B1(n_332),
.B2(n_283),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_338),
.Y(n_449)
);

AND2x2_ASAP7_75t_SL g450 ( 
.A(n_422),
.B(n_312),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_338),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_346),
.A2(n_262),
.B1(n_267),
.B2(n_245),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_R g453 ( 
.A1(n_347),
.A2(n_255),
.B1(n_258),
.B2(n_252),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_415),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_411),
.A2(n_333),
.B1(n_313),
.B2(n_266),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_345),
.B(n_349),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_399),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_395),
.A2(n_272),
.B1(n_279),
.B2(n_278),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

AO22x2_ASAP7_75t_L g460 ( 
.A1(n_354),
.A2(n_373),
.B1(n_390),
.B2(n_359),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_L g461 ( 
.A1(n_413),
.A2(n_292),
.B1(n_298),
.B2(n_287),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_376),
.A2(n_317),
.B1(n_319),
.B2(n_314),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_342),
.Y(n_463)
);

NAND3x1_ASAP7_75t_L g464 ( 
.A(n_348),
.B(n_325),
.C(n_324),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_425),
.A2(n_439),
.B1(n_361),
.B2(n_367),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_350),
.B(n_327),
.Y(n_467)
);

INVx8_ASAP7_75t_L g468 ( 
.A(n_375),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_342),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_424),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_358),
.B(n_209),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_403),
.A2(n_316),
.B1(n_212),
.B2(n_214),
.Y(n_472)
);

AO22x2_ASAP7_75t_L g473 ( 
.A1(n_373),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_434),
.A2(n_224),
.B1(n_226),
.B2(n_221),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_417),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_363),
.B(n_227),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_363),
.Y(n_478)
);

NAND3x1_ASAP7_75t_L g479 ( 
.A(n_353),
.B(n_38),
.C(n_39),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_366),
.B(n_233),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_380),
.B(n_386),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_357),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_342),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_344),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_392),
.B(n_261),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_392),
.B(n_270),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_435),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_406),
.A2(n_273),
.B1(n_275),
.B2(n_271),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_409),
.B(n_276),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_340),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_445),
.A2(n_329),
.B1(n_328),
.B2(n_326),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_362),
.A2(n_391),
.B1(n_393),
.B2(n_384),
.Y(n_493)
);

AO22x2_ASAP7_75t_L g494 ( 
.A1(n_406),
.A2(n_416),
.B1(n_421),
.B2(n_432),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_416),
.A2(n_311),
.B1(n_310),
.B2(n_309),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_382),
.A2(n_308),
.B1(n_304),
.B2(n_301),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_343),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_419),
.Y(n_499)
);

AO22x2_ASAP7_75t_L g500 ( 
.A1(n_432),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_436),
.A2(n_285),
.B1(n_300),
.B2(n_296),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_344),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_344),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_454),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_490),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_449),
.A2(n_429),
.B(n_339),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_491),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_459),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_497),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_451),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_460),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_436),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_468),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_483),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_457),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_465),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_420),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_468),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_463),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_466),
.B(n_426),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_474),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_488),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_498),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_476),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_450),
.B(n_428),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_460),
.B(n_400),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_504),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_463),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_489),
.B(n_426),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_426),
.Y(n_535)
);

XNOR2x2_ASAP7_75t_L g536 ( 
.A(n_452),
.B(n_401),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_469),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_469),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_484),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_501),
.B(n_427),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_467),
.B(n_427),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_473),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_456),
.B(n_441),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_485),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_467),
.B(n_478),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_455),
.B(n_431),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_471),
.B(n_427),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_477),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_462),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_502),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_481),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_480),
.B(n_417),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_486),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_448),
.Y(n_556)
);

AOI21x1_ASAP7_75t_L g557 ( 
.A1(n_487),
.A2(n_352),
.B(n_337),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_448),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_473),
.B(n_446),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_511),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_508),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_506),
.B(n_472),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_514),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_550),
.B(n_475),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_512),
.B(n_341),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_509),
.B(n_518),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_530),
.B(n_500),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_553),
.Y(n_569)
);

BUFx4f_ASAP7_75t_SL g570 ( 
.A(n_514),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_492),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_559),
.A2(n_453),
.B1(n_479),
.B2(n_442),
.Y(n_572)
);

AND2x2_ASAP7_75t_SL g573 ( 
.A(n_543),
.B(n_529),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_531),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_531),
.Y(n_576)
);

OAI21xp33_ASAP7_75t_L g577 ( 
.A1(n_505),
.A2(n_355),
.B(n_383),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_559),
.B(n_458),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_528),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_430),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_526),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_519),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_554),
.B(n_440),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_516),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

INVx3_ASAP7_75t_SL g588 ( 
.A(n_515),
.Y(n_588)
);

AND2x2_ASAP7_75t_SL g589 ( 
.A(n_522),
.B(n_388),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_544),
.B(n_341),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_521),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_513),
.B(n_549),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_552),
.B(n_341),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_549),
.B(n_443),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_524),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_552),
.B(n_370),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_525),
.Y(n_599)
);

NAND2x1p5_ASAP7_75t_L g600 ( 
.A(n_556),
.B(n_443),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_558),
.B(n_370),
.Y(n_601)
);

AND2x2_ASAP7_75t_SL g602 ( 
.A(n_541),
.B(n_397),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_527),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_555),
.B(n_437),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_546),
.B(n_444),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_534),
.B(n_461),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_546),
.B(n_444),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_541),
.B(n_405),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_520),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_532),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_535),
.B(n_496),
.Y(n_612)
);

AND2x2_ASAP7_75t_SL g613 ( 
.A(n_540),
.B(n_407),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_540),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_570),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_581),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_566),
.B(n_536),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_560),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_604),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_569),
.B(n_548),
.Y(n_620)
);

NAND2x1_ASAP7_75t_L g621 ( 
.A(n_584),
.B(n_520),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_592),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_588),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_563),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_571),
.B(n_557),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_589),
.B(n_542),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_576),
.Y(n_627)
);

CKINVDCx6p67_ASAP7_75t_R g628 ( 
.A(n_588),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_584),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_593),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_589),
.B(n_542),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_582),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_584),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_600),
.B(n_464),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_582),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_610),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_561),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_564),
.B(n_607),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_600),
.B(n_533),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_610),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_578),
.B(n_537),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_600),
.B(n_538),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_578),
.B(n_568),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_583),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_589),
.B(n_539),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_580),
.B(n_408),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_594),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_610),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_609),
.B(n_423),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_573),
.B(n_433),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_602),
.B(n_545),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_610),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_601),
.B(n_551),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_596),
.B(n_412),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_594),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_602),
.B(n_372),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_630),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_639),
.B(n_573),
.Y(n_660)
);

INVx6_ASAP7_75t_L g661 ( 
.A(n_615),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_618),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_623),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_643),
.B(n_574),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_617),
.B(n_651),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_628),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_640),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_646),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_630),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_616),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_640),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_645),
.B(n_596),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_630),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_624),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_627),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_616),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_634),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_634),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_629),
.Y(n_679)
);

INVx6_ASAP7_75t_L g680 ( 
.A(n_633),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_655),
.Y(n_681)
);

NAND2x1p5_ASAP7_75t_L g682 ( 
.A(n_633),
.B(n_601),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_631),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_655),
.Y(n_684)
);

NAND2x1p5_ASAP7_75t_L g685 ( 
.A(n_636),
.B(n_601),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_638),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_642),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_631),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_640),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_642),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_652),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_644),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_649),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_654),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_654),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_637),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_657),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_641),
.Y(n_698)
);

BUFx4_ASAP7_75t_R g699 ( 
.A(n_666),
.Y(n_699)
);

INVxp67_ASAP7_75t_SL g700 ( 
.A(n_683),
.Y(n_700)
);

INVxp67_ASAP7_75t_SL g701 ( 
.A(n_683),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_668),
.Y(n_702)
);

INVx6_ASAP7_75t_L g703 ( 
.A(n_661),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_665),
.B(n_622),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_662),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_675),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_661),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_675),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_660),
.A2(n_612),
.B1(n_572),
.B2(n_562),
.Y(n_709)
);

OAI22xp33_ASAP7_75t_L g710 ( 
.A1(n_691),
.A2(n_626),
.B1(n_632),
.B2(n_635),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_679),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_686),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_686),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_693),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_697),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_663),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_664),
.B(n_648),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_688),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_698),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_664),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_L g721 ( 
.A1(n_672),
.A2(n_620),
.B1(n_619),
.B2(n_656),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_672),
.A2(n_591),
.B1(n_603),
.B2(n_599),
.Y(n_722)
);

INVx6_ASAP7_75t_L g723 ( 
.A(n_661),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_667),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_709),
.A2(n_577),
.B1(n_579),
.B2(n_597),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_709),
.A2(n_608),
.B1(n_605),
.B2(n_586),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_702),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_710),
.A2(n_608),
.B1(n_605),
.B2(n_587),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_699),
.Y(n_729)
);

BUFx5_ASAP7_75t_L g730 ( 
.A(n_705),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_704),
.B(n_674),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_700),
.B(n_653),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_717),
.A2(n_689),
.B1(n_692),
.B2(n_671),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_701),
.A2(n_692),
.B1(n_670),
.B2(n_676),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_706),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_708),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_716),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_SL g738 ( 
.A1(n_721),
.A2(n_685),
.B(n_682),
.Y(n_738)
);

OAI222xp33_ASAP7_75t_L g739 ( 
.A1(n_722),
.A2(n_647),
.B1(n_658),
.B2(n_644),
.C1(n_625),
.C2(n_575),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_724),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_714),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_711),
.A2(n_613),
.B1(n_565),
.B2(n_681),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_715),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_712),
.A2(n_565),
.B1(n_684),
.B2(n_601),
.Y(n_744)
);

BUFx12f_ASAP7_75t_L g745 ( 
.A(n_707),
.Y(n_745)
);

OAI21xp33_ASAP7_75t_L g746 ( 
.A1(n_718),
.A2(n_379),
.B(n_369),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_703),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_713),
.A2(n_585),
.B1(n_614),
.B2(n_611),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_719),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_720),
.A2(n_606),
.B1(n_680),
.B2(n_438),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_730),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_728),
.A2(n_723),
.B1(n_690),
.B2(n_694),
.Y(n_752)
);

OAI221xp5_ASAP7_75t_SL g753 ( 
.A1(n_725),
.A2(n_590),
.B1(n_595),
.B2(n_598),
.C(n_687),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_729),
.A2(n_650),
.B1(n_637),
.B2(n_696),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_726),
.A2(n_695),
.B1(n_678),
.B2(n_677),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_742),
.A2(n_567),
.B1(n_678),
.B2(n_677),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_731),
.B(n_659),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_730),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_725),
.A2(n_695),
.B1(n_673),
.B2(n_669),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_733),
.A2(n_673),
.B1(n_669),
.B2(n_659),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_735),
.A2(n_381),
.B1(n_414),
.B2(n_410),
.Y(n_761)
);

OAI221xp5_ASAP7_75t_L g762 ( 
.A1(n_727),
.A2(n_621),
.B1(n_351),
.B2(n_49),
.C(n_50),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_746),
.A2(n_414),
.B1(n_410),
.B2(n_402),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_736),
.A2(n_414),
.B1(n_410),
.B2(n_402),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_738),
.A2(n_402),
.B1(n_394),
.B2(n_389),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_732),
.B(n_51),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_730),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_749),
.A2(n_377),
.B1(n_394),
.B2(n_389),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_744),
.A2(n_371),
.B1(n_387),
.B2(n_385),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_741),
.B(n_360),
.C(n_356),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_748),
.A2(n_371),
.B1(n_387),
.B2(n_385),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_730),
.A2(n_371),
.B1(n_387),
.B2(n_381),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_730),
.Y(n_773)
);

AOI221x1_ASAP7_75t_L g774 ( 
.A1(n_734),
.A2(n_356),
.B1(n_360),
.B2(n_364),
.C(n_365),
.Y(n_774)
);

AOI222xp33_ASAP7_75t_L g775 ( 
.A1(n_739),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.C1(n_57),
.C2(n_59),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_743),
.B(n_60),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_747),
.A2(n_378),
.B1(n_368),
.B2(n_365),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_737),
.B(n_61),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_750),
.A2(n_368),
.B1(n_364),
.B2(n_398),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_757),
.B(n_740),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_758),
.B(n_740),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_766),
.B(n_745),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_775),
.B(n_65),
.C(n_66),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_778),
.B(n_67),
.Y(n_784)
);

NAND3xp33_ASAP7_75t_L g785 ( 
.A(n_762),
.B(n_69),
.C(n_70),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_758),
.B(n_73),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_767),
.B(n_773),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_776),
.B(n_751),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_751),
.B(n_76),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_759),
.B(n_77),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_SL g791 ( 
.A1(n_765),
.A2(n_82),
.B(n_83),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_755),
.B(n_89),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_753),
.B(n_92),
.C(n_93),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_760),
.B(n_95),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_756),
.B(n_752),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_754),
.B(n_100),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_777),
.B(n_101),
.C(n_103),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_SL g798 ( 
.A1(n_770),
.A2(n_104),
.B1(n_107),
.B2(n_109),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_788),
.B(n_772),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_785),
.B(n_763),
.C(n_774),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_781),
.B(n_761),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_783),
.A2(n_779),
.B1(n_771),
.B2(n_769),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_793),
.B(n_768),
.C(n_764),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_786),
.B(n_115),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_782),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_787),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_780),
.B(n_122),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_789),
.B(n_123),
.Y(n_808)
);

AND2x2_ASAP7_75t_SL g809 ( 
.A(n_790),
.B(n_125),
.Y(n_809)
);

BUFx4f_ASAP7_75t_SL g810 ( 
.A(n_784),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_809),
.B(n_790),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_806),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_806),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_810),
.Y(n_814)
);

XNOR2x2_ASAP7_75t_L g815 ( 
.A(n_805),
.B(n_795),
.Y(n_815)
);

NAND4xp75_ASAP7_75t_L g816 ( 
.A(n_808),
.B(n_796),
.C(n_794),
.D(n_792),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_799),
.B(n_791),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_799),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_817),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_818),
.Y(n_820)
);

AO22x1_ASAP7_75t_L g821 ( 
.A1(n_815),
.A2(n_810),
.B1(n_800),
.B2(n_807),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_814),
.Y(n_822)
);

AO22x2_ASAP7_75t_L g823 ( 
.A1(n_811),
.A2(n_801),
.B1(n_803),
.B2(n_807),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_822),
.Y(n_824)
);

OA22x2_ASAP7_75t_L g825 ( 
.A1(n_819),
.A2(n_816),
.B1(n_813),
.B2(n_812),
.Y(n_825)
);

OA22x2_ASAP7_75t_L g826 ( 
.A1(n_821),
.A2(n_813),
.B1(n_804),
.B2(n_807),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_820),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_827),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_824),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_829),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_828),
.A2(n_826),
.B1(n_823),
.B2(n_825),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_828),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_832),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_830),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_831),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_834),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_833),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_836),
.B(n_835),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_837),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_838),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_839),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_841),
.Y(n_842)
);

AOI22x1_ASAP7_75t_L g843 ( 
.A1(n_841),
.A2(n_798),
.B1(n_797),
.B2(n_802),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_SL g844 ( 
.A1(n_840),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_840),
.Y(n_845)
);

AOI22x1_ASAP7_75t_L g846 ( 
.A1(n_845),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_846)
);

OAI22x1_ASAP7_75t_L g847 ( 
.A1(n_843),
.A2(n_139),
.B1(n_141),
.B2(n_144),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_842),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_844),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_845),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_850),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_848),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_847),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_853),
.A2(n_849),
.B1(n_846),
.B2(n_159),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_L g855 ( 
.A1(n_851),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_855),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_854),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_857),
.A2(n_852),
.B1(n_165),
.B2(n_171),
.Y(n_858)
);

AO22x2_ASAP7_75t_L g859 ( 
.A1(n_856),
.A2(n_164),
.B1(n_172),
.B2(n_173),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_859),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_858),
.Y(n_861)
);

AOI221xp5_ASAP7_75t_L g862 ( 
.A1(n_861),
.A2(n_174),
.B1(n_182),
.B2(n_186),
.C(n_191),
.Y(n_862)
);

AOI211xp5_ASAP7_75t_L g863 ( 
.A1(n_862),
.A2(n_860),
.B(n_196),
.C(n_197),
.Y(n_863)
);


endmodule