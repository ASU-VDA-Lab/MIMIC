module fake_jpeg_29039_n_540 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_540);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_434;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

CKINVDCx6p67_ASAP7_75t_R g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_68),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_15),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_69),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_31),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_84),
.B(n_85),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_15),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_21),
.B(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_104),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_21),
.B(n_40),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_109),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_0),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_32),
.B1(n_40),
.B2(n_36),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_150),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_116),
.A2(n_119),
.B1(n_143),
.B2(n_73),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_56),
.A2(n_42),
.B1(n_43),
.B2(n_38),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_32),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_135),
.B(n_160),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_65),
.A2(n_43),
.B1(n_42),
.B2(n_45),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_53),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_145),
.B(n_108),
.C(n_48),
.Y(n_228)
);

NAND2x1_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_53),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_83),
.B(n_20),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_154),
.B(n_164),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_89),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_67),
.B(n_20),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_61),
.A2(n_53),
.B1(n_48),
.B2(n_45),
.Y(n_168)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_81),
.B1(n_80),
.B2(n_70),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_57),
.B(n_19),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_48),
.Y(n_183)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_174),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_175),
.A2(n_196),
.B1(n_226),
.B2(n_142),
.Y(n_263)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

INVx5_ASAP7_75t_SL g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx6p67_ASAP7_75t_R g238 ( 
.A(n_178),
.Y(n_238)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_179),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_188),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_87),
.B1(n_102),
.B2(n_100),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_181),
.A2(n_197),
.B1(n_201),
.B2(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_187),
.Y(n_235)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

OR2x2_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_53),
.Y(n_185)
);

OR2x2_ASAP7_75t_SL g245 ( 
.A(n_185),
.B(n_161),
.Y(n_245)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_49),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_46),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_200),
.Y(n_241)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_192),
.Y(n_267)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_121),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_121),
.A2(n_91),
.B1(n_96),
.B2(n_19),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_133),
.B(n_76),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_213),
.C(n_228),
.Y(n_237)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_123),
.A2(n_34),
.B1(n_30),
.B2(n_51),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_131),
.Y(n_203)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_149),
.A2(n_34),
.B1(n_51),
.B2(n_49),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_30),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_208),
.Y(n_260)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_27),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_137),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_217),
.Y(n_246)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_211),
.Y(n_272)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_212),
.B(n_214),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_48),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_145),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_123),
.A2(n_27),
.B1(n_39),
.B2(n_47),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_220),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_166),
.A2(n_47),
.B1(n_39),
.B2(n_38),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_221),
.B1(n_115),
.B2(n_120),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_129),
.A2(n_45),
.B1(n_93),
.B2(n_103),
.Y(n_221)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_223),
.Y(n_251)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_113),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_124),
.B(n_93),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_134),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_158),
.B1(n_157),
.B2(n_117),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_117),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_183),
.B(n_159),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_233),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

CKINVDCx12_ASAP7_75t_R g236 ( 
.A(n_178),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_236),
.Y(n_291)
);

OA22x2_ASAP7_75t_SL g242 ( 
.A1(n_185),
.A2(n_116),
.B1(n_119),
.B2(n_171),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_242),
.B(n_263),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_245),
.B(n_180),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_198),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_264),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_212),
.A2(n_158),
.B1(n_142),
.B2(n_126),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_270),
.A2(n_130),
.B1(n_128),
.B2(n_229),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_187),
.B(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_206),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_224),
.B(n_46),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_210),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_194),
.B1(n_213),
.B2(n_214),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_274),
.A2(n_282),
.B1(n_237),
.B2(n_264),
.Y(n_312)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_194),
.B(n_228),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_277),
.A2(n_304),
.B(n_256),
.Y(n_332)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_309),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_212),
.B1(n_151),
.B2(n_146),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_280),
.A2(n_257),
.B1(n_177),
.B2(n_195),
.Y(n_313)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_194),
.B1(n_213),
.B2(n_198),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_284),
.A2(n_300),
.B1(n_301),
.B2(n_247),
.Y(n_331)
);

NOR2x1_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_208),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_285),
.B(n_287),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_230),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_286),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_260),
.B(n_225),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_290),
.A2(n_231),
.B(n_268),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_245),
.A2(n_223),
.B1(n_184),
.B2(n_125),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_308),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_293),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_241),
.B(n_174),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_299),
.Y(n_329)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

BUFx4f_ASAP7_75t_SL g299 ( 
.A(n_238),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_263),
.A2(n_130),
.B1(n_128),
.B2(n_125),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_235),
.A2(n_199),
.B1(n_186),
.B2(n_227),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_238),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_302),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_260),
.B(n_190),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_303),
.B(n_307),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_237),
.A2(n_193),
.B(n_192),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_265),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_232),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_235),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_311),
.B(n_320),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_328),
.B1(n_340),
.B2(n_301),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_313),
.A2(n_325),
.B1(n_331),
.B2(n_293),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_271),
.C(n_233),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_297),
.C(n_276),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_233),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_324),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_277),
.A2(n_268),
.B(n_251),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_327),
.B(n_330),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_232),
.C(n_240),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_242),
.B1(n_240),
.B2(n_222),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_242),
.B(n_249),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_289),
.A2(n_266),
.B1(n_176),
.B2(n_255),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_285),
.A2(n_272),
.B(n_265),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_332),
.A2(n_291),
.B(n_281),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_289),
.A2(n_247),
.B1(n_255),
.B2(n_230),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_272),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_292),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_344),
.A2(n_367),
.B(n_373),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_357),
.Y(n_381)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_331),
.A2(n_288),
.B1(n_274),
.B2(n_282),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_347),
.A2(n_317),
.B1(n_286),
.B2(n_250),
.Y(n_392)
);

INVx13_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_330),
.A2(n_288),
.B(n_290),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_250),
.B(n_253),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_351),
.A2(n_354),
.B1(n_369),
.B2(n_327),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_336),
.B1(n_337),
.B2(n_333),
.Y(n_378)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_340),
.A2(n_328),
.B1(n_322),
.B2(n_300),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_319),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_356),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_309),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_359),
.Y(n_384)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_334),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_361),
.Y(n_401)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_311),
.B(n_299),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_275),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_365),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_316),
.B(n_291),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_364),
.B(n_366),
.Y(n_398)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_299),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_259),
.C(n_269),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_284),
.B1(n_278),
.B2(n_306),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_308),
.B(n_307),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_370),
.A2(n_310),
.B(n_252),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_286),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_372),
.B(n_295),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_332),
.A2(n_252),
.B(n_256),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_374),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_375),
.A2(n_376),
.B1(n_382),
.B2(n_385),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_354),
.A2(n_315),
.B1(n_336),
.B2(n_326),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_378),
.A2(n_392),
.B1(n_356),
.B2(n_361),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_351),
.A2(n_326),
.B1(n_324),
.B2(n_312),
.Y(n_382)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_364),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_383),
.B(n_355),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_363),
.A2(n_318),
.B1(n_338),
.B2(n_342),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_320),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_387),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_370),
.A2(n_342),
.B1(n_318),
.B2(n_333),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_389),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_333),
.B1(n_321),
.B2(n_317),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_390),
.A2(n_400),
.B(n_343),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_396),
.C(n_405),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_259),
.C(n_269),
.Y(n_396)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_344),
.B(n_253),
.Y(n_399)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_358),
.B(n_243),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_374),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_243),
.C(n_207),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_344),
.A2(n_347),
.B1(n_357),
.B2(n_349),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_406),
.A2(n_367),
.B1(n_372),
.B2(n_350),
.Y(n_415)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_382),
.B(n_350),
.CI(n_371),
.CON(n_408),
.SN(n_408)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_414),
.Y(n_442)
);

AO22x1_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_349),
.B1(n_355),
.B2(n_373),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_411),
.A2(n_420),
.B1(n_400),
.B2(n_399),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_415),
.A2(n_417),
.B1(n_422),
.B2(n_377),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_353),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_433),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_406),
.A2(n_359),
.B1(n_365),
.B2(n_346),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_262),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_419),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_398),
.B(n_360),
.Y(n_419)
);

INVx11_ASAP7_75t_L g421 ( 
.A(n_380),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_395),
.B(n_262),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_428),
.Y(n_447)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_387),
.B(n_348),
.Y(n_426)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_393),
.B(n_202),
.C(n_248),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_391),
.C(n_388),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_381),
.B(n_295),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_381),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_430),
.Y(n_456)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_431),
.A2(n_432),
.B1(n_434),
.B2(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_405),
.B(n_170),
.Y(n_433)
);

BUFx12_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_1),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_439),
.B(n_443),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_444),
.C(n_452),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_411),
.B(n_375),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_389),
.C(n_402),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_407),
.A2(n_378),
.B1(n_392),
.B2(n_391),
.Y(n_445)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_445),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_453),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_417),
.A2(n_385),
.B1(n_397),
.B2(n_404),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_450),
.A2(n_409),
.B1(n_432),
.B2(n_431),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_411),
.A2(n_399),
.B(n_401),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_420),
.B(n_413),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_390),
.C(n_401),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_415),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_407),
.B(n_394),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_455),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_394),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_403),
.C(n_386),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_458),
.C(n_410),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_408),
.B(n_403),
.C(n_386),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_436),
.B1(n_148),
.B2(n_3),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_442),
.A2(n_409),
.B(n_413),
.Y(n_462)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_441),
.Y(n_479)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_448),
.Y(n_466)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_467),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_439),
.A2(n_412),
.B(n_430),
.Y(n_468)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_408),
.C(n_412),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_471),
.C(n_473),
.Y(n_490)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_456),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_472),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_410),
.C(n_425),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_458),
.B(n_379),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_379),
.C(n_434),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_455),
.C(n_453),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_474),
.B(n_477),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_449),
.A2(n_421),
.B1(n_434),
.B2(n_151),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_475),
.A2(n_446),
.B1(n_450),
.B2(n_447),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_437),
.A2(n_1),
.B(n_2),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_487),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_465),
.B1(n_476),
.B2(n_475),
.Y(n_500)
);

INVx6_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_483),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_441),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_489),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_464),
.A2(n_438),
.B1(n_443),
.B2(n_454),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_491),
.Y(n_498)
);

MAJx2_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_1),
.C(n_2),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_148),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_45),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_465),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_1),
.Y(n_493)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_493),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_463),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_501),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_478),
.A2(n_476),
.B1(n_468),
.B2(n_473),
.Y(n_499)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_499),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_500),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_479),
.B(n_459),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_7),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_45),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_505),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_3),
.C(n_4),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_508),
.C(n_489),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_4),
.C(n_6),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_494),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_493),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_505),
.A2(n_486),
.B(n_485),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_511),
.A2(n_497),
.B(n_508),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_514),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_480),
.C(n_492),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_520),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_495),
.A2(n_491),
.B1(n_8),
.B2(n_10),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_500),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_507),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_7),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_519),
.B(n_11),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_522),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_524),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_507),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_527),
.C(n_512),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_521),
.A2(n_513),
.B(n_526),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_529),
.A2(n_531),
.B(n_517),
.Y(n_534)
);

AOI21xp33_ASAP7_75t_L g532 ( 
.A1(n_530),
.A2(n_521),
.B(n_510),
.Y(n_532)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_533),
.B(n_534),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_SL g533 ( 
.A1(n_528),
.A2(n_526),
.B(n_515),
.C(n_499),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_498),
.B(n_13),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_14),
.B(n_12),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_537),
.A2(n_12),
.B(n_13),
.Y(n_538)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_538),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_12),
.Y(n_540)
);


endmodule