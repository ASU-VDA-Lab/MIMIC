module fake_ariane_838_n_1126 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1126);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1126;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_586;
wire n_443;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_958;
wire n_702;
wire n_905;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_821;
wire n_928;
wire n_1099;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_1026;
wire n_951;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1102;
wire n_975;
wire n_1101;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_976;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_SL g216 ( 
.A(n_16),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_169),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_115),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_12),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_12),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_70),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_94),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_69),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_101),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_48),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_143),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_138),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_105),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_56),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_76),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_161),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_53),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_81),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_43),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_191),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_16),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_86),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_120),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_124),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_66),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_99),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_167),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_104),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_10),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_23),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_78),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_90),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_156),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_150),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_17),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_193),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_51),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_35),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_2),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_203),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_168),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_122),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_20),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_153),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_83),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_95),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_28),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_221),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_226),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_233),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_226),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_272),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_216),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_243),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_260),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_236),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_237),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_241),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_231),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_231),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_283),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

BUFx2_ASAP7_75t_SL g324 ( 
.A(n_246),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_283),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_277),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_218),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_245),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_253),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_219),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_258),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_304),
.B(n_238),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_262),
.B(n_259),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_335),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_295),
.B1(n_333),
.B2(n_334),
.Y(n_339)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_267),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_302),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_284),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_274),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_301),
.B(n_276),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_320),
.A2(n_322),
.B1(n_333),
.B2(n_324),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_223),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_288),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_279),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_286),
.B(n_223),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g365 ( 
.A(n_305),
.B(n_282),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_310),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_331),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_222),
.B(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_291),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_287),
.B(n_223),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_225),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_315),
.A2(n_269),
.B(n_230),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_316),
.B(n_323),
.Y(n_379)
);

AND2x2_ASAP7_75t_SL g380 ( 
.A(n_307),
.B(n_269),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_290),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_294),
.Y(n_382)
);

AOI22x1_ASAP7_75t_SL g383 ( 
.A1(n_322),
.A2(n_280),
.B1(n_278),
.B2(n_275),
.Y(n_383)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_306),
.A2(n_235),
.B(n_228),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_312),
.B(n_239),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_298),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_328),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_309),
.B(n_247),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_300),
.A2(n_250),
.B(n_248),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_327),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_380),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

NOR2x1p5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_292),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_338),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_362),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_339),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

INVx11_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_390),
.B(n_327),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_387),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_366),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_368),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_349),
.B(n_319),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_366),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_345),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_324),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_317),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_338),
.B(n_252),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_348),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_342),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_348),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_390),
.B(n_292),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

OR2x6_ASAP7_75t_L g439 ( 
.A(n_338),
.B(n_293),
.Y(n_439)
);

INVx11_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_352),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_390),
.B(n_293),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_347),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_353),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_353),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_390),
.B(n_256),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_370),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_370),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_390),
.B(n_257),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_354),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_388),
.B(n_261),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_SL g456 ( 
.A(n_369),
.B(n_263),
.Y(n_456)
);

NOR2x1p5_ASAP7_75t_L g457 ( 
.A(n_386),
.B(n_264),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_354),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_347),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_345),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_337),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_354),
.Y(n_463)
);

INVx8_ASAP7_75t_L g464 ( 
.A(n_338),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_369),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_402),
.A2(n_380),
.B(n_378),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_398),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_402),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_393),
.B(n_359),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_437),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_391),
.B(n_359),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_405),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_415),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_415),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_393),
.B(n_344),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_383),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_420),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_420),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_427),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_441),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_427),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_360),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_433),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_433),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_344),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_435),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_424),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_464),
.B(n_389),
.Y(n_490)
);

XNOR2x2_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_336),
.Y(n_491)
);

XNOR2x2_ASAP7_75t_L g492 ( 
.A(n_404),
.B(n_365),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_421),
.B(n_383),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_435),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_464),
.B(n_389),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_438),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_444),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_389),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_361),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_456),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_450),
.Y(n_503)
);

XNOR2x2_ASAP7_75t_L g504 ( 
.A(n_404),
.B(n_365),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_449),
.B(n_388),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_450),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_461),
.A2(n_378),
.B(n_371),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_452),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_445),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_452),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_426),
.B(n_363),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_429),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_454),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_454),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_R g516 ( 
.A(n_439),
.B(n_389),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_458),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_417),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_426),
.B(n_379),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_458),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_462),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_461),
.B(n_449),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_462),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_439),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_463),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_464),
.B(n_344),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_456),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_463),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_439),
.B(n_379),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_448),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_392),
.A2(n_371),
.B(n_384),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_423),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_430),
.B(n_344),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_425),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_425),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_392),
.A2(n_371),
.B(n_384),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_394),
.B(n_355),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_417),
.B(n_379),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_425),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_411),
.B(n_388),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_466),
.A2(n_371),
.B(n_395),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_513),
.B(n_417),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_500),
.B(n_455),
.Y(n_552)
);

NOR2xp67_ASAP7_75t_L g553 ( 
.A(n_512),
.B(n_436),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

NOR3x1_ASAP7_75t_L g555 ( 
.A(n_489),
.B(n_442),
.C(n_519),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_467),
.A2(n_384),
.B1(n_457),
.B2(n_355),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_468),
.B(n_408),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_470),
.B(n_388),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_470),
.B(n_379),
.Y(n_560)
);

OAI221xp5_ASAP7_75t_L g561 ( 
.A1(n_520),
.A2(n_357),
.B1(n_372),
.B2(n_382),
.C(n_381),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_466),
.A2(n_399),
.B(n_397),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_474),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_396),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_475),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g567 ( 
.A(n_483),
.B(n_451),
.C(n_447),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_478),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_472),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_487),
.A2(n_403),
.B(n_401),
.Y(n_570)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_548),
.A2(n_487),
.B(n_479),
.C(n_482),
.Y(n_571)
);

AND2x6_ASAP7_75t_SL g572 ( 
.A(n_477),
.B(n_382),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_548),
.B(n_355),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_545),
.B(n_355),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_481),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_476),
.B(n_446),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_528),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_505),
.A2(n_385),
.B1(n_446),
.B2(n_384),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_467),
.A2(n_446),
.B1(n_372),
.B2(n_399),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_480),
.B(n_397),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_502),
.A2(n_468),
.B1(n_527),
.B2(n_525),
.Y(n_582)
);

BUFx8_ASAP7_75t_L g583 ( 
.A(n_484),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_485),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_509),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_488),
.B(n_400),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_494),
.B(n_400),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_496),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_527),
.B(n_408),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_497),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_539),
.B(n_375),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_498),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_511),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_507),
.A2(n_403),
.B(n_401),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_476),
.B(n_350),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_539),
.B(n_350),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_501),
.B(n_350),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_543),
.B(n_440),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_503),
.B(n_350),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_523),
.B(n_406),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_506),
.B(n_375),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_518),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_508),
.B(n_375),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_510),
.B(n_364),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_514),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_490),
.B(n_495),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_490),
.B(n_364),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_538),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_492),
.A2(n_381),
.B1(n_337),
.B2(n_376),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_502),
.B(n_376),
.Y(n_610)
);

OR2x2_ASAP7_75t_SL g611 ( 
.A(n_504),
.B(n_440),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_491),
.B(n_414),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_516),
.A2(n_495),
.B1(n_499),
.B2(n_523),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_523),
.B(n_414),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_523),
.B(n_406),
.Y(n_615)
);

NAND2x1p5_ASAP7_75t_L g616 ( 
.A(n_499),
.B(n_407),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_516),
.A2(n_412),
.B1(n_410),
.B2(n_409),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_581),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_572),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_610),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_614),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_562),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_551),
.B(n_493),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_554),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_552),
.B(n_515),
.Y(n_626)
);

BUFx4f_ASAP7_75t_L g627 ( 
.A(n_589),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_589),
.B(n_543),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_571),
.A2(n_542),
.B(n_532),
.C(n_517),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_577),
.Y(n_630)
);

AND2x4_ASAP7_75t_SL g631 ( 
.A(n_565),
.B(n_521),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_557),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_SL g633 ( 
.A(n_567),
.B(n_270),
.C(n_265),
.Y(n_633)
);

AOI22x1_ASAP7_75t_L g634 ( 
.A1(n_564),
.A2(n_536),
.B1(n_537),
.B2(n_535),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_583),
.Y(n_635)
);

OR2x2_ASAP7_75t_SL g636 ( 
.A(n_611),
.B(n_337),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_558),
.B(n_337),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_553),
.B(n_569),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_SL g639 ( 
.A(n_561),
.B(n_541),
.C(n_540),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_581),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_559),
.A2(n_542),
.B(n_532),
.C(n_522),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_575),
.A2(n_523),
.B1(n_531),
.B2(n_534),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_614),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_566),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_568),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_579),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_583),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_560),
.B(n_524),
.Y(n_648)
);

AND2x6_ASAP7_75t_SL g649 ( 
.A(n_565),
.B(n_526),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_584),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_598),
.Y(n_651)
);

OR2x2_ASAP7_75t_SL g652 ( 
.A(n_588),
.B(n_529),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_589),
.Y(n_653)
);

NOR3xp33_ASAP7_75t_SL g654 ( 
.A(n_582),
.B(n_590),
.C(n_612),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_585),
.A2(n_533),
.B1(n_547),
.B2(n_549),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_598),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_586),
.Y(n_658)
);

BUFx12f_ASAP7_75t_L g659 ( 
.A(n_616),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_SL g660 ( 
.A(n_592),
.B(n_555),
.C(n_574),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_SL g661 ( 
.A(n_591),
.B(n_546),
.C(n_271),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_596),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_605),
.B(n_431),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_573),
.B(n_407),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_556),
.B(n_431),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_580),
.B(n_409),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_593),
.B(n_410),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_602),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_608),
.B(n_412),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_586),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_618),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_606),
.A2(n_418),
.B1(n_413),
.B2(n_419),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_607),
.B(n_413),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_613),
.B(n_418),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_604),
.B(n_609),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_SL g676 ( 
.A(n_587),
.B(n_507),
.C(n_0),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_587),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_601),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_603),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_616),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_578),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_600),
.B(n_419),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_595),
.B(n_422),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_600),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_657),
.B(n_615),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_621),
.B(n_597),
.Y(n_686)
);

NOR3xp33_ASAP7_75t_L g687 ( 
.A(n_633),
.B(n_550),
.C(n_563),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_676),
.B(n_550),
.C(n_563),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_626),
.B(n_576),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_639),
.A2(n_599),
.B1(n_617),
.B2(n_570),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_648),
.A2(n_594),
.B(n_615),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_625),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_634),
.A2(n_594),
.B(n_422),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_619),
.A2(n_432),
.B1(n_434),
.B2(n_2),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_654),
.B(n_459),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_630),
.B(n_432),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_662),
.B(n_434),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_671),
.B(n_459),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_641),
.A2(n_443),
.B(n_416),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_677),
.B(n_459),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_683),
.A2(n_459),
.B(n_443),
.Y(n_702)
);

NOR2x1_ASAP7_75t_SL g703 ( 
.A(n_628),
.B(n_459),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_673),
.A2(n_443),
.B(n_416),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_623),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_629),
.A2(n_443),
.B(n_416),
.Y(n_706)
);

OAI21x1_ASAP7_75t_SL g707 ( 
.A1(n_675),
.A2(n_346),
.B(n_0),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_622),
.B(n_416),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_624),
.B(n_346),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_619),
.B(n_1),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_631),
.B(n_1),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_SL g712 ( 
.A(n_660),
.B(n_3),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_657),
.B(n_653),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_622),
.B(n_643),
.Y(n_714)
);

INVx6_ASAP7_75t_L g715 ( 
.A(n_649),
.Y(n_715)
);

NAND2x1p5_ASAP7_75t_L g716 ( 
.A(n_643),
.B(n_416),
.Y(n_716)
);

AOI21x1_ASAP7_75t_L g717 ( 
.A1(n_674),
.A2(n_340),
.B(n_443),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_640),
.A2(n_269),
.B(n_340),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_640),
.A2(n_347),
.B(n_34),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_658),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_SL g721 ( 
.A(n_627),
.B(n_269),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_656),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_658),
.B(n_670),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_670),
.A2(n_347),
.B(n_269),
.C(n_5),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_627),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_664),
.A2(n_347),
.B(n_36),
.Y(n_726)
);

AO31x2_ASAP7_75t_L g727 ( 
.A1(n_679),
.A2(n_269),
.A3(n_340),
.B(n_109),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_632),
.B(n_3),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_679),
.A2(n_628),
.B(n_678),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_657),
.B(n_33),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_644),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_652),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_674),
.A2(n_40),
.B(n_38),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_661),
.A2(n_269),
.B(n_5),
.C(n_6),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_643),
.B(n_4),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_672),
.A2(n_44),
.B(n_42),
.Y(n_736)
);

BUFx4f_ASAP7_75t_SL g737 ( 
.A(n_635),
.Y(n_737)
);

OAI21x1_ASAP7_75t_SL g738 ( 
.A1(n_645),
.A2(n_4),
.B(n_6),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_642),
.A2(n_46),
.B(n_45),
.Y(n_739)
);

OAI21x1_ASAP7_75t_SL g740 ( 
.A1(n_650),
.A2(n_655),
.B(n_646),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_665),
.A2(n_340),
.B(n_49),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_667),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_689),
.A2(n_682),
.B(n_666),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_692),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_723),
.B(n_651),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_734),
.A2(n_638),
.B(n_637),
.C(n_663),
.Y(n_746)
);

OAI21xp33_ASAP7_75t_L g747 ( 
.A1(n_724),
.A2(n_647),
.B(n_656),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_718),
.A2(n_681),
.B(n_636),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_720),
.B(n_656),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_737),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_721),
.B(n_699),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_700),
.A2(n_682),
.B(n_666),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_731),
.B(n_686),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_732),
.B(n_620),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_713),
.B(n_680),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_722),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_705),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_721),
.B(n_680),
.Y(n_758)
);

CKINVDCx11_ASAP7_75t_R g759 ( 
.A(n_713),
.Y(n_759)
);

AO31x2_ASAP7_75t_L g760 ( 
.A1(n_690),
.A2(n_681),
.A3(n_684),
.B(n_680),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_SL g761 ( 
.A(n_696),
.B(n_659),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_735),
.A2(n_667),
.B(n_669),
.C(n_9),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_725),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_694),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_710),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_700),
.A2(n_684),
.B(n_669),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_694),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_711),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_740),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_704),
.A2(n_693),
.B(n_741),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_715),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_712),
.A2(n_684),
.B1(n_668),
.B2(n_9),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_717),
.A2(n_668),
.B(n_50),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_SL g774 ( 
.A(n_715),
.B(n_733),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_706),
.A2(n_52),
.B(n_47),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_714),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_688),
.A2(n_709),
.B1(n_728),
.B2(n_695),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_695),
.A2(n_730),
.B1(n_685),
.B2(n_690),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_688),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_779)
);

AOI221x1_ASAP7_75t_L g780 ( 
.A1(n_687),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.C(n_13),
.Y(n_780)
);

OAI21xp33_ASAP7_75t_L g781 ( 
.A1(n_729),
.A2(n_11),
.B(n_13),
.Y(n_781)
);

AO22x2_ASAP7_75t_L g782 ( 
.A1(n_707),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_782)
);

AO32x2_ASAP7_75t_L g783 ( 
.A1(n_727),
.A2(n_14),
.A3(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_783)
);

AOI221x1_ASAP7_75t_L g784 ( 
.A1(n_738),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_702),
.A2(n_127),
.B(n_213),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_691),
.A2(n_21),
.B(n_22),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_697),
.Y(n_787)
);

AO31x2_ASAP7_75t_L g788 ( 
.A1(n_726),
.A2(n_129),
.A3(n_212),
.B(n_210),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_698),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_742),
.B(n_730),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_701),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_SL g792 ( 
.A1(n_736),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_739),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_719),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_703),
.A2(n_28),
.B(n_29),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_708),
.A2(n_134),
.B(n_209),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_SL g797 ( 
.A1(n_685),
.A2(n_29),
.B(n_30),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_716),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_727),
.A2(n_135),
.B(n_208),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_727),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_689),
.A2(n_31),
.B(n_32),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_712),
.B(n_54),
.C(n_55),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_689),
.A2(n_57),
.B(n_58),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_715),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_689),
.B(n_215),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_713),
.Y(n_806)
);

OAI21x1_ASAP7_75t_L g807 ( 
.A1(n_718),
.A2(n_62),
.B(n_63),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_725),
.B(n_64),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_689),
.A2(n_205),
.B(n_67),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_689),
.B(n_204),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_797),
.A2(n_65),
.B1(n_68),
.B2(n_71),
.Y(n_811)
);

BUFx8_ASAP7_75t_L g812 ( 
.A(n_771),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_744),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_SL g814 ( 
.A1(n_800),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_814)
);

BUFx2_ASAP7_75t_SL g815 ( 
.A(n_750),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_753),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_757),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_774),
.B(n_75),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_787),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_759),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_745),
.B(n_82),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_806),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_778),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_806),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_747),
.A2(n_772),
.B1(n_781),
.B2(n_808),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_791),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_763),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_808),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_SL g829 ( 
.A1(n_768),
.A2(n_92),
.B1(n_93),
.B2(n_96),
.Y(n_829)
);

CKINVDCx11_ASAP7_75t_R g830 ( 
.A(n_806),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_756),
.Y(n_831)
);

BUFx10_ASAP7_75t_L g832 ( 
.A(n_765),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_780),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_833)
);

OAI22xp33_ASAP7_75t_L g834 ( 
.A1(n_798),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_754),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_SL g836 ( 
.A1(n_782),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_777),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_755),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_767),
.Y(n_839)
);

INVx6_ASAP7_75t_L g840 ( 
.A(n_790),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_SL g841 ( 
.A1(n_782),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_841)
);

NAND2x1p5_ASAP7_75t_L g842 ( 
.A(n_761),
.B(n_119),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_789),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_793),
.A2(n_126),
.B1(n_131),
.B2(n_133),
.Y(n_844)
);

CKINVDCx6p67_ASAP7_75t_R g845 ( 
.A(n_805),
.Y(n_845)
);

INVx6_ASAP7_75t_L g846 ( 
.A(n_776),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_760),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_749),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_764),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_769),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_779),
.A2(n_136),
.B1(n_137),
.B2(n_140),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_794),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_743),
.B(n_146),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_810),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_801),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_752),
.B(n_151),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_751),
.B(n_152),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_SL g858 ( 
.A1(n_802),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_858)
);

INVx6_ASAP7_75t_L g859 ( 
.A(n_758),
.Y(n_859)
);

INVx3_ASAP7_75t_SL g860 ( 
.A(n_762),
.Y(n_860)
);

INVx8_ASAP7_75t_L g861 ( 
.A(n_795),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_784),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_748),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_786),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_746),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_760),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_804),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_867)
);

BUFx8_ASAP7_75t_L g868 ( 
.A(n_783),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_760),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_796),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_773),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_868),
.A2(n_766),
.B1(n_809),
.B2(n_803),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_SL g873 ( 
.A1(n_865),
.A2(n_811),
.B(n_818),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_813),
.Y(n_874)
);

NAND4xp25_ASAP7_75t_L g875 ( 
.A(n_850),
.B(n_792),
.C(n_783),
.D(n_788),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_832),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_817),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_847),
.B(n_783),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_826),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_866),
.A2(n_770),
.B(n_799),
.Y(n_880)
);

NAND2x1p5_ASAP7_75t_L g881 ( 
.A(n_871),
.B(n_775),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_816),
.B(n_788),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_863),
.B(n_785),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_839),
.B(n_788),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_869),
.Y(n_885)
);

NAND2x1p5_ASAP7_75t_L g886 ( 
.A(n_853),
.B(n_807),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_847),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_840),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_848),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_870),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_856),
.A2(n_166),
.B(n_170),
.Y(n_891)
);

OAI21xp33_ASAP7_75t_SL g892 ( 
.A1(n_825),
.A2(n_171),
.B(n_173),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_822),
.B(n_174),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_870),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_859),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_859),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_861),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_831),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_861),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_827),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_821),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_838),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_845),
.B(n_854),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_849),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_857),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_822),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_824),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_862),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_846),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_846),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_860),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_835),
.Y(n_912)
);

INVx4_ASAP7_75t_SL g913 ( 
.A(n_829),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_830),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_836),
.B(n_841),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_837),
.Y(n_916)
);

OA21x2_ASAP7_75t_L g917 ( 
.A1(n_880),
.A2(n_843),
.B(n_855),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_878),
.B(n_844),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_901),
.B(n_833),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_897),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_883),
.Y(n_921)
);

AO21x2_ASAP7_75t_L g922 ( 
.A1(n_882),
.A2(n_823),
.B(n_852),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_897),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_878),
.B(n_815),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_883),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_885),
.Y(n_926)
);

INVxp67_ASAP7_75t_SL g927 ( 
.A(n_887),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_883),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_885),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_877),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_887),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_894),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_874),
.B(n_828),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_880),
.B(n_814),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_884),
.B(n_842),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_875),
.A2(n_819),
.B(n_851),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_904),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_901),
.B(n_812),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_879),
.B(n_864),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_899),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_886),
.B(n_858),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_886),
.B(n_820),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_873),
.B(n_867),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_886),
.B(n_178),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_890),
.B(n_180),
.Y(n_945)
);

NAND2x1p5_ASAP7_75t_L g946 ( 
.A(n_894),
.B(n_834),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_924),
.B(n_900),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_924),
.B(n_900),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_924),
.B(n_925),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_926),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_926),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_937),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_937),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_931),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_926),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_920),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_931),
.B(n_902),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_942),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_931),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_940),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_929),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_929),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_929),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_920),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_925),
.B(n_908),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_928),
.B(n_899),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_930),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_927),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_918),
.B(n_908),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_930),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_953),
.B(n_919),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_952),
.B(n_969),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_967),
.Y(n_973)
);

AO21x2_ASAP7_75t_L g974 ( 
.A1(n_959),
.A2(n_919),
.B(n_934),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_959),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_968),
.B(n_927),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_967),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_958),
.B(n_942),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_958),
.B(n_942),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_970),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_960),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_964),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_958),
.B(n_928),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_970),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_949),
.B(n_928),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_949),
.B(n_921),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_978),
.B(n_965),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_973),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_971),
.B(n_903),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_972),
.B(n_957),
.Y(n_990)
);

AND2x4_ASAP7_75t_SL g991 ( 
.A(n_978),
.B(n_965),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_982),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_981),
.Y(n_993)
);

NAND2x1_ASAP7_75t_L g994 ( 
.A(n_979),
.B(n_956),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_979),
.B(n_947),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_985),
.B(n_947),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_977),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_975),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_991),
.B(n_985),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_998),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_988),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_992),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_997),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_993),
.B(n_974),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_993),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_1005),
.B(n_994),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1002),
.Y(n_1007)
);

AO221x2_ASAP7_75t_L g1008 ( 
.A1(n_1001),
.A2(n_898),
.B1(n_912),
.B2(n_938),
.C(n_914),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_999),
.B(n_987),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1002),
.B(n_992),
.Y(n_1010)
);

NAND2xp33_ASAP7_75t_SL g1011 ( 
.A(n_1004),
.B(n_987),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1010),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1007),
.B(n_1003),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1009),
.B(n_991),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_1006),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1008),
.Y(n_1016)
);

AOI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_1011),
.A2(n_974),
.B1(n_1000),
.B2(n_989),
.C(n_998),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1010),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1009),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1009),
.B(n_995),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1009),
.B(n_996),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1013),
.Y(n_1023)
);

NOR4xp25_ASAP7_75t_L g1024 ( 
.A(n_1012),
.B(n_1000),
.C(n_989),
.D(n_938),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1020),
.B(n_1018),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_1019),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_1017),
.B(n_913),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_1015),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_1017),
.A2(n_943),
.B(n_873),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1026),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1024),
.B(n_1021),
.Y(n_1031)
);

OAI31xp33_ASAP7_75t_L g1032 ( 
.A1(n_1027),
.A2(n_1016),
.A3(n_915),
.B(n_1014),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_974),
.B1(n_936),
.B2(n_915),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_990),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1029),
.A2(n_936),
.B1(n_913),
.B2(n_943),
.Y(n_1035)
);

AOI321xp33_ASAP7_75t_L g1036 ( 
.A1(n_1022),
.A2(n_934),
.A3(n_941),
.B1(n_872),
.B2(n_918),
.C(n_944),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1023),
.B(n_980),
.Y(n_1037)
);

OAI222xp33_ASAP7_75t_L g1038 ( 
.A1(n_1033),
.A2(n_1025),
.B1(n_943),
.B2(n_914),
.C1(n_934),
.C2(n_911),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1030),
.B(n_984),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1034),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1037),
.Y(n_1041)
);

NAND4xp25_ASAP7_75t_SL g1042 ( 
.A(n_1031),
.B(n_983),
.C(n_976),
.D(n_986),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1032),
.A2(n_1036),
.B(n_1035),
.C(n_943),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1040),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1041),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1039),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1043),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1042),
.B(n_976),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1038),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_1040),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1040),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1050),
.B(n_892),
.C(n_889),
.Y(n_1052)
);

NOR2x1_ASAP7_75t_L g1053 ( 
.A(n_1051),
.B(n_1044),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1046),
.Y(n_1054)
);

AND4x1_ASAP7_75t_L g1055 ( 
.A(n_1046),
.B(n_983),
.C(n_944),
.D(n_909),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1045),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1047),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_L g1058 ( 
.A(n_1049),
.B(n_944),
.C(n_943),
.Y(n_1058)
);

OAI211xp5_ASAP7_75t_SL g1059 ( 
.A1(n_1053),
.A2(n_1048),
.B(n_876),
.C(n_956),
.Y(n_1059)
);

OAI211xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1054),
.A2(n_876),
.B(n_921),
.C(n_916),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1056),
.Y(n_1061)
);

OAI22xp33_ASAP7_75t_SL g1062 ( 
.A1(n_1057),
.A2(n_975),
.B1(n_943),
.B2(n_910),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1058),
.B(n_986),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1061),
.B(n_1055),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_1059),
.B(n_1052),
.Y(n_1065)
);

OAI211xp5_ASAP7_75t_SL g1066 ( 
.A1(n_1063),
.A2(n_921),
.B(n_916),
.C(n_910),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_1060),
.B(n_891),
.C(n_893),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1062),
.B(n_959),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1059),
.A2(n_936),
.B1(n_935),
.B2(n_913),
.Y(n_1069)
);

AOI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1059),
.A2(n_891),
.B(n_941),
.C(n_935),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_1061),
.B(n_893),
.C(n_905),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_SL g1072 ( 
.A(n_1064),
.B(n_895),
.Y(n_1072)
);

NAND4xp75_ASAP7_75t_L g1073 ( 
.A(n_1065),
.B(n_936),
.C(n_941),
.D(n_935),
.Y(n_1073)
);

NAND4xp75_ASAP7_75t_L g1074 ( 
.A(n_1068),
.B(n_936),
.C(n_945),
.D(n_948),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_1069),
.B(n_940),
.Y(n_1075)
);

AND3x4_ASAP7_75t_L g1076 ( 
.A(n_1067),
.B(n_966),
.C(n_893),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_L g1077 ( 
.A(n_1071),
.B(n_945),
.C(n_894),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1070),
.A2(n_1066),
.B(n_948),
.Y(n_1078)
);

AO21x1_ASAP7_75t_L g1079 ( 
.A1(n_1064),
.A2(n_966),
.B(n_946),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1070),
.B(n_954),
.Y(n_1080)
);

XOR2xp5_ASAP7_75t_L g1081 ( 
.A(n_1073),
.B(n_946),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1078),
.B(n_966),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_1080),
.B(n_913),
.C(n_950),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1072),
.B(n_961),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_1077),
.B(n_966),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_1076),
.B(n_932),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1079),
.B(n_962),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_1075),
.B(n_923),
.Y(n_1088)
);

AND4x1_ASAP7_75t_L g1089 ( 
.A(n_1074),
.B(n_933),
.C(n_945),
.D(n_918),
.Y(n_1089)
);

XOR2x1_ASAP7_75t_L g1090 ( 
.A(n_1072),
.B(n_946),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1072),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_1080),
.B(n_906),
.C(n_896),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_1080),
.B(n_957),
.Y(n_1093)
);

NAND5xp2_ASAP7_75t_L g1094 ( 
.A(n_1091),
.B(n_946),
.C(n_933),
.D(n_881),
.E(n_888),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1087),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1089),
.B(n_962),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1083),
.A2(n_950),
.B(n_963),
.C(n_955),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1088),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1090),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1082),
.A2(n_939),
.B1(n_921),
.B2(n_961),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1092),
.A2(n_922),
.B1(n_933),
.B2(n_917),
.Y(n_1101)
);

OAI22x1_ASAP7_75t_L g1102 ( 
.A1(n_1081),
.A2(n_1086),
.B1(n_1085),
.B2(n_1093),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_1098),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1096),
.A2(n_1084),
.B1(n_939),
.B2(n_963),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1097),
.A2(n_955),
.B1(n_951),
.B2(n_932),
.Y(n_1105)
);

INVxp67_ASAP7_75t_SL g1106 ( 
.A(n_1095),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_1099),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1102),
.A2(n_922),
.B1(n_917),
.B2(n_951),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1100),
.A2(n_932),
.B1(n_881),
.B2(n_923),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1106),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1103),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1107),
.A2(n_1101),
.B1(n_1094),
.B2(n_932),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_SL g1113 ( 
.A1(n_1111),
.A2(n_1112),
.B(n_1110),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1113),
.B(n_1104),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1114),
.A2(n_1105),
.B(n_1109),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1114),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_1108),
.B1(n_922),
.B2(n_923),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_922),
.B1(n_917),
.B2(n_907),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1116),
.A2(n_907),
.B1(n_890),
.B2(n_917),
.Y(n_1119)
);

OA21x2_ASAP7_75t_L g1120 ( 
.A1(n_1117),
.A2(n_181),
.B(n_182),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1118),
.A2(n_183),
.B(n_184),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1119),
.A2(n_185),
.B(n_186),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_194),
.B(n_195),
.Y(n_1123)
);

AO221x2_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_196),
.B1(n_197),
.B2(n_199),
.C(n_200),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1124),
.A2(n_1120),
.B1(n_907),
.B2(n_917),
.Y(n_1125)
);

AOI211xp5_ASAP7_75t_L g1126 ( 
.A1(n_1125),
.A2(n_1123),
.B(n_201),
.C(n_202),
.Y(n_1126)
);


endmodule