module real_aes_2342_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_0), .B(n_497), .Y(n_511) );
AOI22xp5_ASAP7_75t_SL g790 ( .A1(n_1), .A2(n_791), .B1(n_794), .B2(n_795), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_1), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_2), .A2(n_496), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_3), .B(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_4), .B(n_286), .Y(n_522) );
INVx1_ASAP7_75t_L g160 ( .A(n_5), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_6), .B(n_179), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_7), .B(n_286), .Y(n_551) );
INVx1_ASAP7_75t_L g188 ( .A(n_8), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_9), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_10), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g592 ( .A(n_11), .B(n_283), .Y(n_592) );
INVx2_ASAP7_75t_L g149 ( .A(n_12), .Y(n_149) );
AOI221x1_ASAP7_75t_L g495 ( .A1(n_13), .A2(n_26), .B1(n_496), .B2(n_497), .C(n_498), .Y(n_495) );
AND3x1_ASAP7_75t_L g113 ( .A(n_14), .B(n_40), .C(n_114), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_14), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_15), .B(n_497), .Y(n_588) );
INVx1_ASAP7_75t_L g284 ( .A(n_16), .Y(n_284) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_17), .A2(n_185), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_18), .B(n_231), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_19), .B(n_286), .Y(n_575) );
AO21x1_ASAP7_75t_L g517 ( .A1(n_20), .A2(n_497), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_21), .Y(n_130) );
INVx1_ASAP7_75t_L g111 ( .A(n_22), .Y(n_111) );
INVx1_ASAP7_75t_L g281 ( .A(n_23), .Y(n_281) );
INVx1_ASAP7_75t_SL g246 ( .A(n_24), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_25), .B(n_166), .Y(n_267) );
AOI33xp33_ASAP7_75t_L g217 ( .A1(n_27), .A2(n_57), .A3(n_155), .B1(n_164), .B2(n_218), .B3(n_219), .Y(n_217) );
NAND2x1_ASAP7_75t_L g509 ( .A(n_28), .B(n_286), .Y(n_509) );
NAND2x1_ASAP7_75t_L g550 ( .A(n_29), .B(n_283), .Y(n_550) );
INVx1_ASAP7_75t_L g197 ( .A(n_30), .Y(n_197) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_31), .A2(n_89), .B(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g180 ( .A(n_31), .B(n_89), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_32), .B(n_174), .Y(n_243) );
INVxp33_ASAP7_75t_L g797 ( .A(n_33), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_34), .B(n_283), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_35), .A2(n_94), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_35), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_36), .B(n_286), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_37), .B(n_283), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_38), .A2(n_496), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g154 ( .A(n_39), .Y(n_154) );
AND2x2_ASAP7_75t_L g172 ( .A(n_39), .B(n_160), .Y(n_172) );
AND2x2_ASAP7_75t_L g178 ( .A(n_39), .B(n_157), .Y(n_178) );
OR2x6_ASAP7_75t_L g129 ( .A(n_40), .B(n_110), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_41), .A2(n_770), .B1(n_775), .B2(n_780), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_42), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_43), .A2(n_54), .B1(n_792), .B2(n_793), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_43), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_44), .B(n_497), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_45), .B(n_174), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_46), .A2(n_147), .B1(n_179), .B2(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_47), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_48), .B(n_166), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_49), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_50), .B(n_283), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_51), .B(n_185), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_52), .B(n_166), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_53), .A2(n_496), .B(n_549), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_54), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_55), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_56), .B(n_283), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_58), .B(n_166), .Y(n_229) );
INVx1_ASAP7_75t_L g159 ( .A(n_59), .Y(n_159) );
INVx1_ASAP7_75t_L g168 ( .A(n_59), .Y(n_168) );
AND2x2_ASAP7_75t_L g230 ( .A(n_60), .B(n_231), .Y(n_230) );
AOI221xp5_ASAP7_75t_L g186 ( .A1(n_61), .A2(n_77), .B1(n_152), .B2(n_174), .C(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_62), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_63), .B(n_286), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_64), .B(n_147), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g151 ( .A1(n_65), .A2(n_152), .B(n_161), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_66), .A2(n_496), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g278 ( .A(n_67), .Y(n_278) );
AO21x1_ASAP7_75t_L g519 ( .A1(n_68), .A2(n_496), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_69), .B(n_497), .Y(n_540) );
INVx1_ASAP7_75t_L g228 ( .A(n_70), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_71), .B(n_497), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_72), .A2(n_152), .B(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g533 ( .A(n_73), .B(n_232), .Y(n_533) );
INVx1_ASAP7_75t_L g157 ( .A(n_74), .Y(n_157) );
INVx1_ASAP7_75t_L g170 ( .A(n_74), .Y(n_170) );
AND2x2_ASAP7_75t_L g553 ( .A(n_75), .B(n_146), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_76), .B(n_174), .Y(n_220) );
AND2x2_ASAP7_75t_L g248 ( .A(n_78), .B(n_146), .Y(n_248) );
INVx1_ASAP7_75t_L g279 ( .A(n_79), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_80), .A2(n_152), .B(n_245), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_81), .A2(n_152), .B(n_212), .C(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g112 ( .A(n_82), .Y(n_112) );
AND2x2_ASAP7_75t_L g538 ( .A(n_83), .B(n_146), .Y(n_538) );
AND2x2_ASAP7_75t_SL g145 ( .A(n_84), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_85), .B(n_497), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_86), .A2(n_152), .B1(n_215), .B2(n_216), .Y(n_214) );
XNOR2xp5_ASAP7_75t_L g770 ( .A(n_87), .B(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g518 ( .A(n_88), .B(n_179), .Y(n_518) );
AND2x2_ASAP7_75t_L g512 ( .A(n_90), .B(n_146), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_91), .B(n_283), .Y(n_576) );
INVx1_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_93), .B(n_286), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_94), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_95), .B(n_283), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_96), .A2(n_496), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g221 ( .A(n_97), .B(n_146), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_98), .B(n_286), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_99), .A2(n_195), .B(n_196), .C(n_199), .Y(n_194) );
BUFx2_ASAP7_75t_L g133 ( .A(n_100), .Y(n_133) );
BUFx2_ASAP7_75t_SL g786 ( .A(n_100), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_101), .A2(n_496), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_102), .B(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_117), .B(n_796), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g798 ( .A(n_107), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_113), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_134), .B(n_784), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_131), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_121), .A2(n_788), .B(n_789), .Y(n_787) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_130), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_125), .Y(n_788) );
BUFx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
OR2x6_ASAP7_75t_SL g483 ( .A(n_127), .B(n_128), .Y(n_483) );
AND2x6_ASAP7_75t_SL g487 ( .A(n_127), .B(n_129), .Y(n_487) );
OR2x2_ASAP7_75t_L g783 ( .A(n_127), .B(n_129), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI21xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_770), .B(n_774), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_481), .B1(n_484), .B2(n_488), .Y(n_136) );
INVx2_ASAP7_75t_L g779 ( .A(n_137), .Y(n_779) );
BUFx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND3x1_ASAP7_75t_L g138 ( .A(n_139), .B(n_371), .C(n_436), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_325), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_270), .B(n_298), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_233), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_181), .Y(n_142) );
AOI21xp33_ASAP7_75t_L g372 ( .A1(n_143), .A2(n_373), .B(n_384), .Y(n_372) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_143), .B(n_314), .Y(n_407) );
AND2x2_ASAP7_75t_L g422 ( .A(n_143), .B(n_423), .Y(n_422) );
OR2x6_ASAP7_75t_L g432 ( .A(n_143), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g434 ( .A(n_143), .B(n_424), .Y(n_434) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g308 ( .A(n_144), .Y(n_308) );
AND2x2_ASAP7_75t_L g321 ( .A(n_144), .B(n_322), .Y(n_321) );
INVx4_ASAP7_75t_L g340 ( .A(n_144), .Y(n_340) );
AND2x2_ASAP7_75t_L g343 ( .A(n_144), .B(n_259), .Y(n_343) );
NOR2x1_ASAP7_75t_SL g346 ( .A(n_144), .B(n_274), .Y(n_346) );
AND2x4_ASAP7_75t_L g358 ( .A(n_144), .B(n_356), .Y(n_358) );
OR2x2_ASAP7_75t_L g368 ( .A(n_144), .B(n_240), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_144), .B(n_380), .Y(n_385) );
OR2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_150), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_146), .A2(n_194), .B1(n_200), .B2(n_201), .Y(n_193) );
INVx3_ASAP7_75t_L g201 ( .A(n_146), .Y(n_201) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_147), .B(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx4f_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
AND2x4_ASAP7_75t_L g179 ( .A(n_149), .B(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_149), .B(n_180), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_173), .B(n_179), .Y(n_150) );
INVxp67_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_158), .Y(n_152) );
NOR2x1p5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx1_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OR2x6_ASAP7_75t_L g163 ( .A(n_156), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x6_ASAP7_75t_L g283 ( .A(n_157), .B(n_167), .Y(n_283) );
AND2x6_ASAP7_75t_L g496 ( .A(n_158), .B(n_178), .Y(n_496) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx2_ASAP7_75t_L g164 ( .A(n_159), .Y(n_164) );
AND2x4_ASAP7_75t_L g286 ( .A(n_159), .B(n_169), .Y(n_286) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_165), .C(n_171), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_SL g187 ( .A1(n_163), .A2(n_171), .B(n_188), .C(n_189), .Y(n_187) );
INVxp67_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_163), .A2(n_171), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g245 ( .A1(n_163), .A2(n_171), .B(n_246), .C(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g269 ( .A(n_163), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_163), .A2(n_198), .B1(n_278), .B2(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g175 ( .A(n_164), .B(n_176), .Y(n_175) );
INVxp33_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
INVx1_ASAP7_75t_L g198 ( .A(n_166), .Y(n_198) );
AND2x4_ASAP7_75t_L g497 ( .A(n_166), .B(n_172), .Y(n_497) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_169), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g215 ( .A(n_171), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_171), .A2(n_267), .B(n_268), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_171), .B(n_179), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_171), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_171), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_171), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_171), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_171), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_171), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_171), .A2(n_575), .B(n_576), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_171), .A2(n_591), .B(n_592), .Y(n_590) );
INVx5_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_172), .Y(n_199) );
INVx1_ASAP7_75t_L g208 ( .A(n_174), .Y(n_208) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g262 ( .A(n_175), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_177), .Y(n_263) );
BUFx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_179), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_SL g571 ( .A(n_179), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_179), .A2(n_588), .B(n_589), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_181), .A2(n_314), .B1(n_409), .B2(n_410), .Y(n_408) );
INVx1_ASAP7_75t_SL g452 ( .A(n_181), .Y(n_452) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_209), .Y(n_181) );
INVx2_ASAP7_75t_L g383 ( .A(n_182), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_182), .B(n_329), .Y(n_455) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_191), .Y(n_182) );
BUFx3_ASAP7_75t_L g301 ( .A(n_183), .Y(n_301) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g294 ( .A(n_184), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_184), .B(n_211), .Y(n_316) );
AND2x4_ASAP7_75t_L g333 ( .A(n_184), .B(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g349 ( .A(n_184), .Y(n_349) );
INVx2_ASAP7_75t_L g406 ( .A(n_184), .Y(n_406) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_190), .Y(n_184) );
INVx2_ASAP7_75t_SL g212 ( .A(n_185), .Y(n_212) );
AND2x2_ASAP7_75t_L g324 ( .A(n_191), .B(n_290), .Y(n_324) );
NOR2xp67_ASAP7_75t_L g370 ( .A(n_191), .B(n_293), .Y(n_370) );
AND2x2_ASAP7_75t_L g389 ( .A(n_191), .B(n_293), .Y(n_389) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g251 ( .A(n_192), .Y(n_251) );
INVx1_ASAP7_75t_L g332 ( .A(n_192), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_192), .B(n_223), .Y(n_351) );
AND2x4_ASAP7_75t_L g405 ( .A(n_192), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_202), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_201), .A2(n_224), .B(n_230), .Y(n_223) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_201), .A2(n_224), .B(n_230), .Y(n_293) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_201), .A2(n_506), .B(n_512), .Y(n_505) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_201), .A2(n_527), .B(n_533), .Y(n_526) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_201), .A2(n_527), .B(n_533), .Y(n_560) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_201), .A2(n_506), .B(n_512), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g364 ( .A(n_209), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_209), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_222), .Y(n_209) );
AND2x2_ASAP7_75t_L g348 ( .A(n_210), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g388 ( .A(n_210), .Y(n_388) );
AND2x2_ASAP7_75t_L g393 ( .A(n_210), .B(n_293), .Y(n_393) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_211), .B(n_223), .Y(n_253) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_221), .Y(n_211) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_212), .A2(n_213), .B(n_221), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_214), .B(n_220), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g329 ( .A(n_222), .Y(n_329) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_222), .B(n_301), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_222), .B(n_251), .Y(n_468) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_223), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_231), .Y(n_241) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_231), .A2(n_495), .B(n_501), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_231), .A2(n_540), .B(n_541), .Y(n_539) );
OA21x2_ASAP7_75t_L g640 ( .A1(n_231), .A2(n_495), .B(n_501), .Y(n_640) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OAI21xp33_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_249), .B(n_254), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_236), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g306 ( .A(n_237), .Y(n_306) );
AND2x2_ASAP7_75t_L g320 ( .A(n_237), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g354 ( .A(n_237), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g420 ( .A(n_237), .B(n_338), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_237), .B(n_467), .C(n_468), .Y(n_466) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_238), .Y(n_297) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
AND2x2_ASAP7_75t_L g319 ( .A(n_240), .B(n_274), .Y(n_319) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_240), .Y(n_330) );
AND2x2_ASAP7_75t_L g375 ( .A(n_240), .B(n_273), .Y(n_375) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_240), .Y(n_398) );
INVx1_ASAP7_75t_L g415 ( .A(n_240), .Y(n_415) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_248), .Y(n_240) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_241), .A2(n_547), .B(n_553), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g457 ( .A(n_249), .Y(n_457) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_250), .B(n_328), .Y(n_429) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g291 ( .A(n_251), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI211x1_ASAP7_75t_L g325 ( .A1(n_255), .A2(n_326), .B(n_335), .C(n_352), .Y(n_325) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_256), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g378 ( .A(n_256), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g314 ( .A(n_258), .B(n_273), .Y(n_314) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g272 ( .A(n_259), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_259), .Y(n_339) );
INVx1_ASAP7_75t_L g356 ( .A(n_259), .Y(n_356) );
AND2x2_ASAP7_75t_L g424 ( .A(n_259), .B(n_274), .Y(n_424) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_265), .Y(n_259) );
NOR3xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .C(n_264), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_288), .B(n_295), .Y(n_270) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_271), .B(n_340), .Y(n_443) );
INVx2_ASAP7_75t_L g475 ( .A(n_271), .Y(n_475) );
INVx4_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g307 ( .A(n_272), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g380 ( .A(n_273), .Y(n_380) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g322 ( .A(n_274), .Y(n_322) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_287), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_284), .B2(n_285), .Y(n_280) );
INVxp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
OR2x2_ASAP7_75t_L g382 ( .A(n_289), .B(n_383), .Y(n_382) );
NAND2x1_ASAP7_75t_SL g404 ( .A(n_289), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g304 ( .A(n_290), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
INVx1_ASAP7_75t_L g458 ( .A(n_291), .Y(n_458) );
AND2x2_ASAP7_75t_L g323 ( .A(n_292), .B(n_324), .Y(n_323) );
NOR2x1_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g305 ( .A(n_293), .Y(n_305) );
INVxp33_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g362 ( .A(n_297), .B(n_355), .Y(n_362) );
OAI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B(n_309), .C(n_317), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g386 ( .A(n_300), .B(n_387), .Y(n_386) );
NOR2xp67_ASAP7_75t_SL g391 ( .A(n_300), .B(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_301), .B(n_388), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_303), .B(n_307), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
AND2x2_ASAP7_75t_L g435 ( .A(n_304), .B(n_405), .Y(n_435) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_307), .A2(n_454), .B1(n_456), .B2(n_459), .C1(n_460), .C2(n_463), .Y(n_453) );
INVx1_ASAP7_75t_L g417 ( .A(n_308), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_315), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_313), .Y(n_344) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_313), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g433 ( .A(n_314), .Y(n_433) );
AND2x2_ASAP7_75t_L g478 ( .A(n_314), .B(n_330), .Y(n_478) );
AND2x2_ASAP7_75t_L g359 ( .A(n_315), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g472 ( .A(n_316), .B(n_351), .Y(n_472) );
OAI21xp33_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_320), .B(n_323), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_318), .A2(n_338), .B(n_379), .Y(n_439) );
AND2x2_ASAP7_75t_L g463 ( .A(n_319), .B(n_340), .Y(n_463) );
NOR2xp33_ASAP7_75t_SL g473 ( .A(n_319), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g411 ( .A(n_322), .Y(n_411) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_322), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g446 ( .A(n_324), .Y(n_446) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_331), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g449 ( .A(n_329), .B(n_333), .Y(n_449) );
BUFx2_ASAP7_75t_L g337 ( .A(n_330), .Y(n_337) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g360 ( .A(n_332), .Y(n_360) );
INVx2_ASAP7_75t_L g366 ( .A(n_332), .Y(n_366) );
AND2x2_ASAP7_75t_L g402 ( .A(n_332), .B(n_393), .Y(n_402) );
AND2x4_ASAP7_75t_L g369 ( .A(n_333), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g409 ( .A(n_333), .B(n_366), .Y(n_409) );
AND2x2_ASAP7_75t_L g460 ( .A(n_333), .B(n_461), .Y(n_460) );
AOI31xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_341), .A3(n_345), .B(n_347), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
AND2x2_ASAP7_75t_L g357 ( .A(n_337), .B(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_SL g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x4_ASAP7_75t_L g355 ( .A(n_340), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_343), .A2(n_395), .B1(n_426), .B2(n_429), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_343), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g480 ( .A(n_343), .B(n_396), .Y(n_480) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g395 ( .A(n_346), .B(n_396), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AND2x2_ASAP7_75t_L g418 ( .A(n_348), .B(n_389), .Y(n_418) );
INVx1_ASAP7_75t_L g428 ( .A(n_350), .Y(n_428) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_361), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g451 ( .A(n_354), .Y(n_451) );
AND2x2_ASAP7_75t_L g459 ( .A(n_355), .B(n_411), .Y(n_459) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_355), .Y(n_465) );
AND2x2_ASAP7_75t_L g410 ( .A(n_358), .B(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_363), .B1(n_367), .B2(n_369), .Y(n_361) );
NOR2xp33_ASAP7_75t_SL g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_364), .A2(n_383), .B1(n_477), .B2(n_479), .Y(n_476) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g376 ( .A(n_369), .Y(n_376) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_399), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
OAI21xp33_ASAP7_75t_L g377 ( .A1(n_375), .A2(n_378), .B(n_381), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_378), .A2(n_402), .B1(n_403), .B2(n_407), .Y(n_401) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_390), .B2(n_394), .Y(n_384) );
INVx1_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2xp67_ASAP7_75t_L g399 ( .A(n_400), .B(n_412), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_408), .Y(n_400) );
INVx2_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
NAND2xp33_ASAP7_75t_SL g454 ( .A(n_404), .B(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g427 ( .A(n_405), .Y(n_427) );
INVx3_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
INVxp67_ASAP7_75t_L g470 ( .A(n_410), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_413), .B(n_421), .C(n_425), .D(n_430), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
AND2x2_ASAP7_75t_L g423 ( .A(n_415), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g471 ( .A(n_419), .Y(n_471) );
NAND2xp33_ASAP7_75t_SL g426 ( .A(n_427), .B(n_428), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B(n_435), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND3x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_453), .C(n_464), .Y(n_436) );
AOI221x1_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_442), .B2(n_444), .C(n_450), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp33_ASAP7_75t_SL g444 ( .A(n_445), .B(n_448), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NAND2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_469), .C(n_476), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_469) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_482), .Y(n_778) );
CKINVDCx11_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
CKINVDCx6p67_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
CKINVDCx11_ASAP7_75t_R g776 ( .A(n_485), .Y(n_776) );
INVx3_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g777 ( .A(n_488), .Y(n_777) );
XNOR2x2_ASAP7_75t_SL g789 ( .A(n_488), .B(n_790), .Y(n_789) );
NAND4xp75_ASAP7_75t_L g488 ( .A(n_489), .B(n_680), .C(n_720), .D(n_749), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_642), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_599), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_534), .B(n_554), .Y(n_491) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_493), .B(n_502), .Y(n_492) );
AND2x4_ASAP7_75t_L g598 ( .A(n_493), .B(n_559), .Y(n_598) );
INVx1_ASAP7_75t_SL g651 ( .A(n_493), .Y(n_651) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_493), .A2(n_687), .B(n_690), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_SL g690 ( .A1(n_493), .A2(n_691), .B(n_692), .C(n_693), .Y(n_690) );
NAND2x1_ASAP7_75t_L g731 ( .A(n_493), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_493), .B(n_692), .Y(n_753) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g557 ( .A(n_494), .Y(n_557) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_494), .Y(n_630) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_513), .Y(n_502) );
AND2x2_ASAP7_75t_L g622 ( .A(n_503), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g703 ( .A(n_503), .B(n_559), .Y(n_703) );
INVx1_ASAP7_75t_L g763 ( .A(n_503), .Y(n_763) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g607 ( .A(n_504), .B(n_525), .Y(n_607) );
AND2x2_ASAP7_75t_L g732 ( .A(n_504), .B(n_526), .Y(n_732) );
AND2x2_ASAP7_75t_L g737 ( .A(n_504), .B(n_697), .Y(n_737) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVxp67_ASAP7_75t_L g613 ( .A(n_505), .Y(n_613) );
BUFx3_ASAP7_75t_L g646 ( .A(n_505), .Y(n_646) );
AND2x2_ASAP7_75t_L g692 ( .A(n_505), .B(n_526), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
AND2x2_ASAP7_75t_L g677 ( .A(n_513), .B(n_556), .Y(n_677) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_525), .Y(n_513) );
AND2x4_ASAP7_75t_L g559 ( .A(n_514), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g669 ( .A(n_514), .B(n_653), .Y(n_669) );
AND2x2_ASAP7_75t_SL g712 ( .A(n_514), .B(n_640), .Y(n_712) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g648 ( .A(n_515), .Y(n_648) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g609 ( .A(n_516), .Y(n_609) );
OAI21x1_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_519), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g524 ( .A(n_518), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_525), .B(n_609), .Y(n_612) );
AND2x2_ASAP7_75t_L g697 ( .A(n_525), .B(n_640), .Y(n_697) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g694 ( .A(n_526), .B(n_557), .Y(n_694) );
AND2x2_ASAP7_75t_L g714 ( .A(n_526), .B(n_640), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_528), .B(n_532), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_534), .B(n_603), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_534), .A2(n_726), .B1(n_727), .B2(n_728), .C(n_730), .Y(n_725) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI332xp33_ASAP7_75t_L g759 ( .A1(n_535), .A2(n_619), .A3(n_626), .B1(n_685), .B2(n_760), .B3(n_761), .C1(n_762), .C2(n_764), .Y(n_759) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_536), .B(n_545), .Y(n_535) );
AND2x2_ASAP7_75t_L g565 ( .A(n_536), .B(n_546), .Y(n_565) );
AND2x2_ASAP7_75t_L g582 ( .A(n_536), .B(n_583), .Y(n_582) );
INVx4_ASAP7_75t_L g594 ( .A(n_536), .Y(n_594) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_536), .B(n_595), .Y(n_654) );
INVx5_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR2x1_ASAP7_75t_SL g616 ( .A(n_537), .B(n_583), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_537), .B(n_545), .Y(n_620) );
AND2x2_ASAP7_75t_L g627 ( .A(n_537), .B(n_546), .Y(n_627) );
BUFx2_ASAP7_75t_L g662 ( .A(n_537), .Y(n_662) );
AND2x2_ASAP7_75t_L g717 ( .A(n_537), .B(n_586), .Y(n_717) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OR2x2_ASAP7_75t_L g585 ( .A(n_545), .B(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g595 ( .A(n_545), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g635 ( .A(n_545), .Y(n_635) );
AND2x2_ASAP7_75t_L g705 ( .A(n_545), .B(n_604), .Y(n_705) );
AND2x2_ASAP7_75t_L g718 ( .A(n_545), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_545), .B(n_719), .Y(n_736) );
INVx4_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_546), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
OAI32xp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_561), .A3(n_566), .B1(n_580), .B2(n_597), .Y(n_554) );
INVx2_ASAP7_75t_L g663 ( .A(n_555), .Y(n_663) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g674 ( .A(n_556), .Y(n_674) );
BUFx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g608 ( .A(n_557), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g741 ( .A(n_557), .B(n_646), .Y(n_741) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g653 ( .A(n_560), .Y(n_653) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx2_ASAP7_75t_L g641 ( .A(n_563), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_563), .B(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x4_ASAP7_75t_SL g652 ( .A(n_564), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g729 ( .A(n_564), .Y(n_729) );
AND2x2_ASAP7_75t_L g747 ( .A(n_564), .B(n_609), .Y(n_747) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp67_ASAP7_75t_SL g691 ( .A(n_567), .B(n_620), .Y(n_691) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_568), .B(n_602), .Y(n_689) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g765 ( .A(n_569), .B(n_635), .Y(n_765) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g596 ( .A(n_570), .Y(n_596) );
INVx2_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B(n_578), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_571), .B(n_579), .Y(n_578) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_571), .A2(n_572), .B(n_578), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_577), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_593), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_581), .B(n_639), .Y(n_724) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND3x2_ASAP7_75t_L g679 ( .A(n_582), .B(n_626), .C(n_635), .Y(n_679) );
AND2x2_ASAP7_75t_L g603 ( .A(n_583), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_583), .B(n_586), .Y(n_660) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g614 ( .A(n_585), .B(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g604 ( .A(n_586), .Y(n_604) );
INVx1_ASAP7_75t_L g619 ( .A(n_586), .Y(n_619) );
BUFx3_ASAP7_75t_L g626 ( .A(n_586), .Y(n_626) );
AND2x2_ASAP7_75t_L g636 ( .A(n_586), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x4_ASAP7_75t_L g645 ( .A(n_594), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_594), .B(n_604), .Y(n_688) );
AND2x2_ASAP7_75t_L g644 ( .A(n_595), .B(n_619), .Y(n_644) );
INVx2_ASAP7_75t_L g671 ( .A(n_595), .Y(n_671) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_605), .B(n_610), .C(n_631), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g751 ( .A1(n_600), .A2(n_727), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_603), .B(n_662), .Y(n_661) );
AOI211xp5_ASAP7_75t_SL g681 ( .A1(n_603), .A2(n_682), .B(n_686), .C(n_695), .Y(n_681) );
AND2x2_ASAP7_75t_L g667 ( .A(n_604), .B(n_627), .Y(n_667) );
OR2x2_ASAP7_75t_L g670 ( .A(n_604), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_607), .B(n_712), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_608), .B(n_653), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_608), .A2(n_634), .B1(n_714), .B2(n_717), .C(n_723), .Y(n_722) );
AND2x4_ASAP7_75t_L g639 ( .A(n_609), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g685 ( .A(n_609), .B(n_640), .Y(n_685) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_614), .B1(n_617), .B2(n_621), .C(n_624), .Y(n_610) );
AND2x2_ASAP7_75t_L g756 ( .A(n_611), .B(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g623 ( .A(n_612), .Y(n_623) );
INVx1_ASAP7_75t_L g709 ( .A(n_613), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_614), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g628 ( .A(n_616), .B(n_619), .Y(n_628) );
AND2x2_ASAP7_75t_L g704 ( .A(n_616), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g629 ( .A(n_623), .B(n_630), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_628), .B(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g748 ( .A(n_625), .Y(n_748) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g727 ( .A(n_626), .B(n_654), .Y(n_727) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_627), .B(n_636), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_638), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_632), .A2(n_666), .B1(n_669), .B2(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g738 ( .A(n_632), .Y(n_738) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g658 ( .A(n_635), .Y(n_658) );
INVx1_ASAP7_75t_L g719 ( .A(n_637), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_639), .B(n_641), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_639), .B(n_709), .Y(n_760) );
AND2x2_ASAP7_75t_L g728 ( .A(n_640), .B(n_729), .Y(n_728) );
OAI211xp5_ASAP7_75t_L g721 ( .A1(n_641), .A2(n_722), .B(n_725), .C(n_733), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_664), .Y(n_642) );
AOI322xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .A3(n_647), .B1(n_649), .B2(n_654), .C1(n_655), .C2(n_663), .Y(n_643) );
CKINVDCx16_ASAP7_75t_R g761 ( .A(n_645), .Y(n_761) );
AND2x2_ASAP7_75t_L g711 ( .A(n_646), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g745 ( .A(n_646), .Y(n_745) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_SL g696 ( .A(n_648), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_SL g702 ( .A(n_648), .B(n_694), .Y(n_702) );
AND2x2_ASAP7_75t_L g726 ( .A(n_648), .B(n_692), .Y(n_726) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g698 ( .A(n_652), .Y(n_698) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_661), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI221xp5_ASAP7_75t_SL g701 ( .A1(n_657), .A2(n_702), .B1(n_703), .B2(n_704), .C(n_706), .Y(n_701) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g768 ( .A(n_660), .Y(n_768) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B(n_668), .C(n_672), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g743 ( .A(n_667), .Y(n_743) );
INVx1_ASAP7_75t_L g675 ( .A(n_669), .Y(n_675) );
OR2x2_ASAP7_75t_L g762 ( .A(n_669), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_SL g758 ( .A(n_670), .Y(n_758) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B(n_678), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_674), .B(n_692), .Y(n_769) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_701), .Y(n_680) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_684), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
OR2x2_ASAP7_75t_L g735 ( .A(n_688), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI21xp33_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_698), .B(n_699), .Y(n_695) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
AOI31xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .A3(n_713), .B(n_715), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_712), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_737), .B1(n_738), .B2(n_739), .C(n_742), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_746), .B2(n_748), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_759), .C(n_766), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_751), .B(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_758), .Y(n_754) );
INVxp67_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI22x1_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g794 ( .A(n_791), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
endmodule