module fake_jpeg_10762_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_62),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_59),
.Y(n_74)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_22),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_47),
.C(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_2),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_49),
.B(n_37),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_43),
.B1(n_44),
.B2(n_39),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_57),
.B1(n_40),
.B2(n_61),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_43),
.B1(n_37),
.B2(n_49),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_71),
.B1(n_72),
.B2(n_6),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_51),
.B1(n_39),
.B2(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_51),
.B1(n_45),
.B2(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_52),
.B1(n_50),
.B2(n_42),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_75),
.A3(n_66),
.B1(n_74),
.B2(n_69),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_88),
.B1(n_85),
.B2(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_5),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_5),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_89),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_87),
.B1(n_9),
.B2(n_10),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_6),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_8),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_9),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_103),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_90),
.B1(n_78),
.B2(n_83),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_104),
.B(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_26),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_30),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_20),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_11),
.B(n_13),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_10),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_32),
.B(n_12),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.C(n_115),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_11),
.B(n_14),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_15),
.B(n_17),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_105),
.B1(n_97),
.B2(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

AO221x1_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_102),
.B1(n_96),
.B2(n_113),
.C(n_33),
.Y(n_121)
);

AOI21x1_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_118),
.B(n_119),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_119),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_122),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_109),
.B1(n_94),
.B2(n_111),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_99),
.Y(n_128)
);


endmodule