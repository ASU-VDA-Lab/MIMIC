module fake_jpeg_27593_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_14),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_19),
.C(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_58),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_32),
.C(n_33),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_63),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_34),
.B1(n_28),
.B2(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_57),
.B1(n_46),
.B2(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_64),
.Y(n_76)
);

AOI22x1_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_28),
.B1(n_34),
.B2(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_62),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_30),
.B(n_14),
.C(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_36),
.C(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_41),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_70),
.B(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_38),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_38),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_44),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_15),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_57),
.B(n_63),
.C(n_44),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_52),
.C(n_61),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_91),
.C(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_92),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_75),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_61),
.B1(n_46),
.B2(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_82),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_44),
.C(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_38),
.B(n_44),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_30),
.B(n_36),
.C(n_27),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_101),
.C(n_91),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_93),
.B(n_88),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_104),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_73),
.C(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_107),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_82),
.B(n_77),
.C(n_27),
.D(n_24),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_87),
.A3(n_23),
.B1(n_96),
.B2(n_84),
.C1(n_88),
.C2(n_90),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_97),
.C(n_98),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_94),
.B(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_101),
.B1(n_103),
.B2(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_110),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_112),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_11),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_6),
.B(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_8),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_121),
.B1(n_117),
.B2(n_122),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_123),
.A3(n_124),
.B1(n_7),
.B2(n_6),
.C1(n_1),
.C2(n_4),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_1),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_132),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_133),
.B1(n_2),
.B2(n_3),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_136),
.Y(n_138)
);


endmodule