module real_aes_7224_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_55;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_53;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_54;
wire n_51;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_50;
wire n_38;
wire n_23;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR2xp33_ASAP7_75t_R g21 ( .A(n_0), .B(n_22), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g43 ( .A(n_0), .Y(n_43) );
NAND2xp33_ASAP7_75t_SL g49 ( .A(n_0), .B(n_50), .Y(n_49) );
NAND2xp33_ASAP7_75t_SL g18 ( .A(n_1), .B(n_19), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g29 ( .A(n_1), .B(n_30), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g35 ( .A(n_1), .B(n_36), .Y(n_35) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_1), .B(n_15), .Y(n_42) );
CKINVDCx20_ASAP7_75t_R g54 ( .A(n_1), .Y(n_54) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_2), .Y(n_27) );
NOR3xp33_ASAP7_75t_SL g25 ( .A(n_3), .B(n_9), .C(n_26), .Y(n_25) );
AOI221xp5_ASAP7_75t_SL g32 ( .A1(n_4), .A2(n_6), .B1(n_33), .B2(n_37), .C(n_44), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_5), .B(n_20), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_5), .Y(n_31) );
NAND2xp33_ASAP7_75t_SL g38 ( .A(n_5), .B(n_39), .Y(n_38) );
CKINVDCx20_ASAP7_75t_R g55 ( .A(n_7), .Y(n_55) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_8), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_10), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_11), .Y(n_17) );
INVx1_ASAP7_75t_L g52 ( .A(n_12), .Y(n_52) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_13), .Y(n_23) );
NOR4xp25_ASAP7_75t_SL g37 ( .A(n_13), .B(n_38), .C(n_41), .D(n_43), .Y(n_37) );
NOR2xp33_ASAP7_75t_R g46 ( .A(n_13), .B(n_47), .Y(n_46) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_14), .Y(n_22) );
NAND4xp25_ASAP7_75t_SL g20 ( .A(n_15), .B(n_21), .C(n_23), .D(n_24), .Y(n_20) );
OAI221xp5_ASAP7_75t_R g16 ( .A1(n_17), .A2(n_18), .B1(n_28), .B2(n_29), .C(n_32), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g36 ( .A(n_19), .Y(n_36) );
NOR2xp33_ASAP7_75t_R g30 ( .A(n_20), .B(n_31), .Y(n_30) );
NAND2xp33_ASAP7_75t_SL g40 ( .A(n_22), .B(n_24), .Y(n_40) );
AND2x2_ASAP7_75t_L g24 ( .A(n_25), .B(n_27), .Y(n_24) );
NAND2xp33_ASAP7_75t_SL g53 ( .A(n_30), .B(n_54), .Y(n_53) );
NAND2xp33_ASAP7_75t_SL g51 ( .A(n_31), .B(n_39), .Y(n_51) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_35), .Y(n_34) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g41 ( .A(n_42), .Y(n_41) );
NAND2xp33_ASAP7_75t_SL g47 ( .A(n_42), .B(n_48), .Y(n_47) );
OAI22xp33_ASAP7_75t_SL g44 ( .A1(n_45), .A2(n_52), .B1(n_53), .B2(n_55), .Y(n_44) );
CKINVDCx16_ASAP7_75t_R g45 ( .A(n_46), .Y(n_45) );
CKINVDCx5p33_ASAP7_75t_R g48 ( .A(n_49), .Y(n_48) );
CKINVDCx20_ASAP7_75t_R g50 ( .A(n_51), .Y(n_50) );
endmodule