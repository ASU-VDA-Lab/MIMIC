module fake_jpeg_17174_n_189 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_33),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_0),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_27),
.C(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_27),
.B(n_16),
.C(n_26),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_38),
.A2(n_18),
.B1(n_15),
.B2(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_20),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_55),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_36),
.C(n_32),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_75),
.C(n_15),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_66),
.B(n_0),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_26),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_36),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_32),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_70),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_31),
.B1(n_21),
.B2(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_37),
.B(n_18),
.C(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_24),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_19),
.B1(n_18),
.B2(n_15),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_82),
.B1(n_83),
.B2(n_69),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_66),
.B(n_63),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_7),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_91),
.B1(n_96),
.B2(n_99),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_1),
.B(n_4),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_90),
.B(n_75),
.C(n_72),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_73),
.B1(n_51),
.B2(n_69),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_118),
.B1(n_119),
.B2(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_50),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_120),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_110),
.B(n_111),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_78),
.B1(n_79),
.B2(n_98),
.Y(n_126)
);

AO221x1_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_58),
.B1(n_74),
.B2(n_66),
.C(n_76),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_69),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_114),
.B(n_119),
.C(n_104),
.D(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_115),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_66),
.B(n_67),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_78),
.B(n_79),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_6),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_66),
.B1(n_10),
.B2(n_11),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_126),
.B(n_108),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_79),
.B1(n_78),
.B2(n_98),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_137),
.B1(n_83),
.B2(n_77),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_81),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_132),
.B(n_97),
.C(n_84),
.D(n_82),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_95),
.C(n_87),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.C(n_96),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_116),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_143),
.C(n_134),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_122),
.C(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_84),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_145),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_130),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_97),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_150),
.B1(n_133),
.B2(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_146),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_149),
.B(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_138),
.B1(n_143),
.B2(n_147),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_142),
.C(n_134),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_124),
.B1(n_156),
.B2(n_150),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_153),
.B(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_164),
.B(n_165),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_123),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_127),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_158),
.C(n_161),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_130),
.B(n_136),
.Y(n_169)
);

NAND4xp25_ASAP7_75t_SL g171 ( 
.A(n_165),
.B(n_160),
.C(n_151),
.D(n_124),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_176),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_131),
.B(n_168),
.C(n_85),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_127),
.B(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_180),
.C(n_113),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_133),
.Y(n_180)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_173),
.B(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_184),
.B(n_178),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_181),
.B(n_102),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_186),
.B(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_11),
.Y(n_189)
);


endmodule