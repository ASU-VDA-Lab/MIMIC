module fake_jpeg_29727_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_20),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_62),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_15),
.B1(n_40),
.B2(n_38),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_47),
.B1(n_46),
.B2(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_48),
.B1(n_53),
.B2(n_50),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_78),
.B1(n_53),
.B2(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_86),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_96),
.B1(n_8),
.B2(n_9),
.Y(n_112)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_52),
.A3(n_54),
.B1(n_45),
.B2(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_41),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_1),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_7),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_2),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_97),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_19),
.B1(n_36),
.B2(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_3),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_101),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_23),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_5),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_31),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_7),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_111),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_117),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_12),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_13),
.B1(n_14),
.B2(n_21),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_22),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_120),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_32),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_106),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_125),
.A2(n_99),
.B1(n_117),
.B2(n_120),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_121),
.B1(n_127),
.B2(n_109),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_135),
.CI(n_121),
.CON(n_139),
.SN(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_136),
.B1(n_139),
.B2(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_128),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_126),
.C(n_124),
.Y(n_143)
);

AOI21x1_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_119),
.B(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);


endmodule