module fake_jpeg_15353_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_21),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_0),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_52),
.B(n_45),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_74),
.C(n_5),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_53),
.B1(n_55),
.B2(n_49),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_73),
.B1(n_77),
.B2(n_6),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_58),
.B1(n_51),
.B2(n_50),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_54),
.A3(n_46),
.B1(n_22),
.B2(n_24),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_4),
.Y(n_88)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_64),
.B1(n_54),
.B2(n_46),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_86),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_89),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_91),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_44),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_92),
.Y(n_105)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_4),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_8),
.C(n_10),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_7),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_101),
.B1(n_83),
.B2(n_15),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_109),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_80),
.B1(n_81),
.B2(n_16),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_111),
.B1(n_103),
.B2(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_112),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_83),
.B(n_17),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_13),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_99),
.B1(n_19),
.B2(n_20),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_116),
.B1(n_113),
.B2(n_99),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_120),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_115),
.B(n_120),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_18),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_23),
.C(n_25),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_27),
.C(n_28),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_30),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_42),
.C(n_35),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_33),
.CI(n_36),
.CON(n_129),
.SN(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_41),
.B(n_37),
.C(n_38),
.Y(n_130)
);


endmodule