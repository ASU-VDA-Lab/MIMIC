module fake_jpeg_18909_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_9),
.B(n_0),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_3),
.Y(n_21)
);

AND2x6_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_17),
.B1(n_19),
.B2(n_18),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_14),
.B1(n_20),
.B2(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_31),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_17),
.B1(n_19),
.B2(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_20),
.Y(n_47)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_37),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_10),
.CI(n_16),
.CON(n_45),
.SN(n_45)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_47),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_23),
.C(n_21),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.C(n_45),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_32),
.C(n_37),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_41),
.C(n_42),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_36),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_52),
.C(n_53),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_5),
.C(n_6),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_8),
.C(n_9),
.Y(n_53)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_46),
.C(n_43),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_61),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_41),
.C(n_44),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_38),
.B(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_61),
.C(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_59),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_44),
.A3(n_57),
.B1(n_59),
.B2(n_60),
.C1(n_62),
.C2(n_67),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_70),
.CI(n_57),
.CON(n_71),
.SN(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_66),
.Y(n_72)
);


endmodule