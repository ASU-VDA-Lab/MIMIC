module real_jpeg_8559_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_288, n_6, n_7, n_289, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_288;
input n_6;
input n_7;
input n_289;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_215;
wire n_83;
wire n_221;
wire n_166;
wire n_176;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_278;
wire n_130;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_279;
wire n_59;
wire n_88;
wire n_128;
wire n_244;
wire n_202;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_1),
.A2(n_11),
.B1(n_18),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_29),
.B1(n_39),
.B2(n_41),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_1),
.A2(n_29),
.B1(n_63),
.B2(n_64),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_2),
.A2(n_9),
.B(n_26),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_62)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_5),
.A2(n_39),
.B(n_62),
.C(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_5),
.B(n_39),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_5),
.A2(n_9),
.B(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_11),
.B1(n_18),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_8),
.A2(n_39),
.B1(n_41),
.B2(n_58),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_58),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_9),
.A2(n_11),
.B1(n_18),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_39),
.B1(n_41),
.B2(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_9),
.B(n_36),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_50),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_25),
.B(n_38),
.C(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_9),
.B(n_27),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_10),
.A2(n_11),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_10),
.A2(n_19),
.B1(n_63),
.B2(n_64),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_10),
.A2(n_19),
.B1(n_39),
.B2(n_41),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_22),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_22),
.B(n_50),
.C(n_169),
.Y(n_168)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_281),
.B(n_284),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_71),
.B(n_280),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_30),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_15),
.B(n_30),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_15),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_15),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_27),
.B2(n_28),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_24),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_21),
.A2(n_24),
.B1(n_49),
.B2(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_21),
.B(n_24),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_37),
.B(n_38),
.C(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_48),
.B(n_57),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_28),
.B(n_238),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_31),
.B(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_31),
.B(n_278),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_46),
.CI(n_51),
.CON(n_31),
.SN(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_36),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_35),
.B(n_129),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_43),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_36),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_36),
.A2(n_43),
.B1(n_127),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_37),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_39),
.A2(n_42),
.B(n_50),
.Y(n_133)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_41),
.A2(n_50),
.B(n_67),
.C(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_44),
.B(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_49),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_50),
.B(n_62),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.C(n_59),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_52),
.A2(n_59),
.B1(n_258),
.B2(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_52),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_53),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_54),
.A2(n_55),
.B1(n_143),
.B2(n_149),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_54),
.B(n_143),
.C(n_186),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_54),
.A2(n_55),
.B1(n_126),
.B2(n_130),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_54),
.B(n_126),
.C(n_215),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_54),
.A2(n_55),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_59),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_59),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_70),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_61),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_62),
.A2(n_68),
.B1(n_92),
.B2(n_95),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_62),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_62),
.A2(n_68),
.B1(n_70),
.B2(n_221),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_63),
.B(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_277),
.B(n_279),
.Y(n_71)
);

OAI321xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_250),
.A3(n_270),
.B1(n_275),
.B2(n_276),
.C(n_288),
.Y(n_72)
);

AOI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_205),
.A3(n_225),
.B1(n_244),
.B2(n_249),
.C(n_289),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_174),
.C(n_202),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_154),
.B(n_173),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_139),
.B(n_153),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_121),
.B(n_138),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_110),
.B(n_120),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_100),
.B(n_109),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_89),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_81),
.A2(n_102),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_81),
.B(n_143),
.C(n_148),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_84),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_84),
.A2(n_136),
.B1(n_181),
.B2(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_85),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_86),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_87),
.A2(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_97),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_99),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_126),
.C(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_90),
.A2(n_99),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_94),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_95),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_99),
.B(n_179),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_108),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_106),
.B(n_107),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_107),
.A2(n_113),
.B1(n_114),
.B2(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_115),
.C(n_118),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_107),
.A2(n_119),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_112),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_118),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_117),
.A2(n_118),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_117),
.B(n_193),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_142),
.C(n_152),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_123),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_131),
.B2(n_137),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_130),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_160),
.C(n_164),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_128),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_135),
.B(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_150),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_149),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_149),
.B(n_231),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_155),
.B(n_156),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_166),
.C(n_172),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_164),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_163),
.A2(n_164),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_163),
.A2(n_164),
.B1(n_264),
.B2(n_268),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_163),
.B(n_258),
.C(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_163),
.B(n_268),
.C(n_269),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_197),
.C(n_199),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_166),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_187),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_176),
.B(n_187),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_183),
.CI(n_184),
.CON(n_176),
.SN(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_201),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_196),
.C(n_201),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_245),
.B(n_248),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_207),
.B(n_208),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_224),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_216),
.B2(n_217),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_217),
.C(n_224),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_223),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_218),
.A2(n_219),
.B1(n_236),
.B2(n_239),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_220),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_234),
.B(n_236),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_220),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_227),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_242),
.B2(n_243),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_233),
.B1(n_240),
.B2(n_241),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_241),
.C(n_243),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_252),
.C(n_260),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_252),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_233),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_262),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_255),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_261),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);


endmodule