module fake_ariane_931_n_3785 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_541, n_499, n_12, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_363, n_720, n_354, n_41, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_733, n_761, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_738, n_758, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_753, n_566, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_721, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_510, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_769, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_3785);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_363;
input n_720;
input n_354;
input n_41;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_510;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_769;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_3785;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_3765;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_2238;
wire n_1503;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_3416;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_829;
wire n_1062;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_795;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_3315;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_2650;
wire n_863;
wire n_1254;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2391;
wire n_2332;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_1013;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1840;
wire n_1230;
wire n_2739;
wire n_3739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_2956;
wire n_2382;
wire n_1213;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_3458;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_2909;
wire n_1121;
wire n_1416;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_1594;
wire n_2806;
wire n_1935;
wire n_3191;
wire n_1716;
wire n_3777;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_851;
wire n_1590;
wire n_3280;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_3698;
wire n_3716;
wire n_1179;
wire n_3284;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_1884;
wire n_912;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_3678;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_2970;
wire n_3159;
wire n_992;
wire n_966;
wire n_955;
wire n_3549;
wire n_3624;
wire n_2855;
wire n_794;
wire n_1182;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_3538;
wire n_1376;
wire n_1292;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1178;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_3530;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3629;
wire n_3666;
wire n_3372;
wire n_1623;
wire n_990;
wire n_3559;
wire n_1903;
wire n_867;
wire n_2147;
wire n_3479;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3724;
wire n_1920;
wire n_2083;
wire n_815;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_3046;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_3741;
wire n_2388;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_3496;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_976;
wire n_3567;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3127;
wire n_1731;
wire n_799;
wire n_2829;
wire n_1147;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_965;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3397;
wire n_1111;
wire n_1689;
wire n_970;
wire n_2535;
wire n_3467;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3179;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_2558;
wire n_2996;
wire n_1496;
wire n_1217;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3615;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_3642;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3513;
wire n_3498;
wire n_3682;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_2067;
wire n_1134;
wire n_3374;
wire n_3471;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_3508;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_3477;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_1726;
wire n_2075;
wire n_3263;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3569;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1614;
wire n_1162;
wire n_2031;
wire n_3260;
wire n_3349;
wire n_3761;
wire n_2118;
wire n_3222;
wire n_1740;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_2802;
wire n_1963;
wire n_1104;
wire n_3653;
wire n_3035;
wire n_887;
wire n_3403;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_1202;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_3602;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3501;
wire n_3492;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2949;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_3766;
wire n_1711;
wire n_1219;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_1791;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_3417;
wire n_2449;
wire n_890;
wire n_842;
wire n_3626;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1373;
wire n_1975;
wire n_1081;
wire n_1388;
wire n_2119;
wire n_1540;
wire n_1719;
wire n_1266;
wire n_2742;
wire n_3671;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_2623;
wire n_3392;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_3065;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_3367;
wire n_3669;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_3024;
wire n_951;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3208;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1714;
wire n_1044;
wire n_2696;
wire n_3340;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_3302;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_2489;
wire n_1161;
wire n_3685;
wire n_811;
wire n_3097;
wire n_3507;
wire n_791;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_2622;
wire n_3447;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_1318;
wire n_854;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3422;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1873;
wire n_1137;
wire n_1733;
wire n_1856;
wire n_1258;
wire n_1476;
wire n_1524;
wire n_2723;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_3167;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3746;
wire n_961;
wire n_1807;
wire n_1046;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_1784;
wire n_3110;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_3753;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_2936;
wire n_1154;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_3718;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_2329;
wire n_979;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_3455;
wire n_807;
wire n_3736;
wire n_891;
wire n_3313;
wire n_1659;
wire n_885;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_3317;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_3605;
wire n_3345;
wire n_2170;
wire n_3560;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_3654;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_2605;
wire n_2796;
wire n_1201;
wire n_858;
wire n_2804;
wire n_2475;
wire n_1185;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_2665;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_3769;
wire n_825;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_914;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_1197;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3731;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_3444;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_2343;
wire n_1048;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_2935;
wire n_889;
wire n_3255;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1534;
wire n_1948;
wire n_1065;
wire n_3006;
wire n_2767;
wire n_810;
wire n_3376;
wire n_3381;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_3770;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_1968;
wire n_918;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_3288;
wire n_3251;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_3405;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_1749;
wire n_820;
wire n_872;
wire n_1653;
wire n_3409;
wire n_3522;
wire n_3583;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3241;
wire n_1584;
wire n_1157;
wire n_848;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3553;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_3751;
wire n_3402;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_2951;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_932;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2503;
wire n_2270;
wire n_3470;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_2865;
wire n_1204;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3677;
wire n_1564;
wire n_2010;
wire n_3676;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3576;
wire n_3558;
wire n_3782;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3658;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_3521;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_1663;
wire n_919;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_956;
wire n_3360;
wire n_1930;
wire n_3687;
wire n_1809;
wire n_2787;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_3575;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3633;
wire n_898;
wire n_857;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_2012;
wire n_1937;
wire n_3182;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_3316;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_3776;
wire n_2775;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_2351;
wire n_1619;
wire n_3303;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_2206;
wire n_997;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3232;
wire n_3001;
wire n_3188;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1136;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_3094;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3441;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_865;
wire n_1983;
wire n_1273;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_1923;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_3763;
wire n_1946;
wire n_2148;
wire n_933;
wire n_3244;
wire n_3499;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_1821;
wire n_1168;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3593;
wire n_2673;
wire n_2585;
wire n_1591;
wire n_3293;
wire n_2995;
wire n_3361;
wire n_1683;
wire n_1229;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_3707;
wire n_2052;
wire n_2485;
wire n_1091;
wire n_3779;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2275;
wire n_2183;
wire n_2205;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_3058;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_2792;
wire n_1146;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3592;
wire n_3725;
wire n_2269;
wire n_1474;
wire n_2081;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_2361;
wire n_1001;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3075;
wire n_3030;
wire n_3505;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_3547;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_2239;
wire n_1252;
wire n_1129;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_3041;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g782 ( 
.A(n_166),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_520),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_557),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_491),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_636),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_602),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_57),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_768),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_561),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_694),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_315),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_464),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_658),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_386),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_442),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_374),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_274),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_35),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_27),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_745),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_180),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_212),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_655),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_411),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_73),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_95),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_302),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_240),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_590),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_694),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_71),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_38),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_413),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_625),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_2),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_157),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_718),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_758),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_612),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_492),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_539),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_467),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_448),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_370),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_738),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_327),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_83),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_171),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_348),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_232),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_257),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_375),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_45),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_602),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_729),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_696),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_205),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_24),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_382),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_603),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_384),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_69),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_261),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_775),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_415),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_123),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_737),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_50),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_672),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_35),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_448),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_536),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_132),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_8),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_102),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_538),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_688),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_746),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_258),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_105),
.Y(n_861)
);

BUFx2_ASAP7_75t_SL g862 ( 
.A(n_387),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_321),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_734),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_138),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_256),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_581),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_768),
.Y(n_868)
);

BUFx10_ASAP7_75t_L g869 ( 
.A(n_420),
.Y(n_869)
);

BUFx10_ASAP7_75t_L g870 ( 
.A(n_350),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_24),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_410),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_215),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_723),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_605),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_331),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_212),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_624),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_684),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_646),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_535),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_473),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_250),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_700),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_394),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_570),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_690),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_766),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_432),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_8),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_184),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_705),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_643),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_390),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_264),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_670),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_763),
.Y(n_897)
);

BUFx5_ASAP7_75t_L g898 ( 
.A(n_214),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_106),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_732),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_269),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_586),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_320),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_387),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_546),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_13),
.Y(n_906)
);

CKINVDCx14_ASAP7_75t_R g907 ( 
.A(n_720),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_117),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_56),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_381),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_713),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_310),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_95),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_699),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_305),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_2),
.Y(n_916)
);

CKINVDCx14_ASAP7_75t_R g917 ( 
.A(n_750),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_246),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_67),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_720),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_439),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_728),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_630),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_287),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_709),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_131),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_571),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_700),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_93),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_124),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_323),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_583),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_43),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_675),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_238),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_402),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_452),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_742),
.Y(n_938)
);

BUFx10_ASAP7_75t_L g939 ( 
.A(n_326),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_735),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_0),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_31),
.Y(n_942)
);

CKINVDCx16_ASAP7_75t_R g943 ( 
.A(n_759),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_208),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_497),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_274),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_320),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_244),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_117),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_776),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_318),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_749),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_688),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_7),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_475),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_315),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_138),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_619),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_211),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_266),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_735),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_697),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_718),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_457),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_41),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_96),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_593),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_46),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_288),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_540),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_748),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_738),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_730),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_211),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_498),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_299),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_3),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_253),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_538),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_414),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_518),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_601),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_708),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_490),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_73),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_484),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_526),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_692),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_719),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_365),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_397),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_189),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_423),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_69),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_151),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_46),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_15),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_473),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_730),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_74),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_668),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_486),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_617),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_582),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_659),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_409),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_507),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_524),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_617),
.Y(n_1009)
);

CKINVDCx16_ASAP7_75t_R g1010 ( 
.A(n_398),
.Y(n_1010)
);

CKINVDCx16_ASAP7_75t_R g1011 ( 
.A(n_186),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_163),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_37),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_306),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_469),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_725),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_254),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_740),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_726),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_301),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_686),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_594),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_733),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_422),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_5),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_283),
.Y(n_1026)
);

BUFx5_ASAP7_75t_L g1027 ( 
.A(n_392),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_660),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_158),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_124),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_251),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_169),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_754),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_471),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_23),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_353),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_769),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_103),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_352),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_399),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_685),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_200),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_755),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_295),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_97),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_301),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_668),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_392),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_528),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_442),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_102),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_83),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_699),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_386),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_479),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_619),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_775),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_550),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_79),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_134),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_178),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_224),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_466),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_194),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_696),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_778),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_563),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_371),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_166),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_390),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_743),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_280),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_134),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_49),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_241),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_376),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_533),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_487),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_728),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_512),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_633),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_754),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_457),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_623),
.Y(n_1084)
);

CKINVDCx14_ASAP7_75t_R g1085 ( 
.A(n_234),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_552),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_466),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_667),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_220),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_553),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_547),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_736),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_372),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_407),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_36),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_294),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_549),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_519),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_155),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_219),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_145),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_597),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_645),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_344),
.Y(n_1104)
);

CKINVDCx14_ASAP7_75t_R g1105 ( 
.A(n_756),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_724),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_436),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_610),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_27),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_584),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_571),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_183),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_45),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_519),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_354),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_639),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_343),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_348),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_37),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_743),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_593),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_176),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_133),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_498),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_366),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_631),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_49),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_370),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_377),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_492),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_472),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_268),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_611),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_558),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_243),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_373),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_733),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_618),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_384),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_205),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_625),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_172),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_496),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_481),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_406),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_418),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_271),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_582),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_76),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_741),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_218),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_249),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_476),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_225),
.Y(n_1154)
);

INVxp33_ASAP7_75t_R g1155 ( 
.A(n_643),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_488),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_533),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_221),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_72),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_542),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_237),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_635),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_616),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_373),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_177),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_31),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_329),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_399),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_488),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_400),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_330),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_344),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_136),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_567),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_747),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_707),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_57),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_25),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_731),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_125),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_769),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_601),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_716),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_34),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_477),
.Y(n_1185)
);

INVxp33_ASAP7_75t_SL g1186 ( 
.A(n_118),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_19),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_751),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_416),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_54),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_493),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_255),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_232),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_650),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_749),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_722),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_137),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_299),
.Y(n_1198)
);

INVx4_ASAP7_75t_R g1199 ( 
.A(n_355),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_368),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_610),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_368),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_761),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_744),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_250),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_258),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_779),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_441),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_647),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_613),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_757),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_115),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_452),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_159),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_337),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_272),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_123),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_722),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_243),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_714),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_482),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_105),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_389),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_254),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_673),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_47),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_106),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_692),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_396),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_213),
.Y(n_1230)
);

BUFx10_ASAP7_75t_L g1231 ( 
.A(n_774),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_142),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_752),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_739),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_70),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_188),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_729),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_676),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_750),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_675),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_627),
.Y(n_1241)
);

BUFx5_ASAP7_75t_L g1242 ( 
.A(n_424),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_494),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_514),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_187),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_358),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_361),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_744),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_624),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_103),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_136),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_505),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_239),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_760),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_113),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_302),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_268),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_633),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_753),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_704),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_11),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_18),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_674),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_721),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_737),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_408),
.Y(n_1266)
);

CKINVDCx16_ASAP7_75t_R g1267 ( 
.A(n_411),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_42),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_686),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_99),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_195),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_359),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_229),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_660),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_539),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_724),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_717),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_61),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_291),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_266),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_152),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_441),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_603),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_727),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_424),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_453),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_284),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_676),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_147),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_209),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_162),
.Y(n_1291)
);

CKINVDCx14_ASAP7_75t_R g1292 ( 
.A(n_80),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_459),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_563),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_284),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_428),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_404),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_200),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_558),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_396),
.Y(n_1300)
);

INVxp67_ASAP7_75t_SL g1301 ( 
.A(n_803),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_803),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_868),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_848),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_848),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1066),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_865),
.Y(n_1307)
);

INVxp33_ASAP7_75t_SL g1308 ( 
.A(n_856),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_865),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_946),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_809),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_946),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_943),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_996),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_996),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1006),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_817),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1010),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_907),
.B(n_0),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1006),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1016),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1016),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_902),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_917),
.Y(n_1324)
);

CKINVDCx14_ASAP7_75t_R g1325 ( 
.A(n_1085),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_847),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1058),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_914),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_1058),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1090),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1011),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1099),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_1090),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_898),
.Y(n_1334)
);

CKINVDCx14_ASAP7_75t_R g1335 ( 
.A(n_1105),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_1102),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1102),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1117),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1115),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1115),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1126),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1263),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1126),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1128),
.Y(n_1344)
);

INVxp33_ASAP7_75t_L g1345 ( 
.A(n_1082),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1128),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1267),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1292),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1169),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_873),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1169),
.Y(n_1351)
);

CKINVDCx16_ASAP7_75t_R g1352 ( 
.A(n_869),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_869),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1239),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_898),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1239),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_853),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1249),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_871),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1249),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_898),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_898),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_898),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_898),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_898),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_898),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_991),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_875),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1027),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1027),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1027),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_879),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1027),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1027),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1027),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1027),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1027),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1242),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_880),
.Y(n_1379)
);

INVxp33_ASAP7_75t_L g1380 ( 
.A(n_1084),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1242),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_800),
.Y(n_1382)
);

INVxp33_ASAP7_75t_SL g1383 ( 
.A(n_785),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1242),
.Y(n_1384)
);

BUFx8_ASAP7_75t_SL g1385 ( 
.A(n_889),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1242),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1242),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_897),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1242),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1242),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_800),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1207),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1242),
.Y(n_1393)
);

CKINVDCx16_ASAP7_75t_R g1394 ( 
.A(n_869),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_782),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_783),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_881),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_784),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_800),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_800),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_789),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_800),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_791),
.Y(n_1403)
);

CKINVDCx16_ASAP7_75t_R g1404 ( 
.A(n_870),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_792),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_838),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_802),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_838),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_804),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_807),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_814),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_816),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_818),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_823),
.Y(n_1414)
);

INVxp33_ASAP7_75t_L g1415 ( 
.A(n_1153),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_882),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_909),
.Y(n_1417)
);

INVxp67_ASAP7_75t_SL g1418 ( 
.A(n_838),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1175),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_838),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_825),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_838),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_827),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_842),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_844),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_845),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_849),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_851),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_855),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_857),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_874),
.Y(n_1431)
);

INVxp33_ASAP7_75t_SL g1432 ( 
.A(n_785),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_877),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_866),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_866),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_878),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_883),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1361),
.A2(n_876),
.B(n_813),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1406),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1382),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1362),
.A2(n_876),
.B(n_813),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1406),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1406),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1303),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1402),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1402),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1334),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1334),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1350),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1355),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1406),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1391),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1392),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1399),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1366),
.A2(n_1025),
.B(n_994),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1355),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1400),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1323),
.B(n_1297),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1408),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1313),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1363),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1399),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1325),
.B(n_870),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1363),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1434),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1301),
.B(n_1186),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1418),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1434),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1364),
.Y(n_1469)
);

BUFx8_ASAP7_75t_SL g1470 ( 
.A(n_1385),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1369),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1364),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1365),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1370),
.A2(n_1025),
.B(n_994),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1379),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1365),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1311),
.A2(n_974),
.B1(n_1007),
.B2(n_929),
.Y(n_1477)
);

AND2x6_ASAP7_75t_L g1478 ( 
.A(n_1378),
.B(n_1037),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1378),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1420),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1371),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1373),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1374),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1353),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1375),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1376),
.A2(n_1052),
.B(n_1037),
.Y(n_1486)
);

INVx5_ASAP7_75t_L g1487 ( 
.A(n_1392),
.Y(n_1487)
);

INVx5_ASAP7_75t_L g1488 ( 
.A(n_1324),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1325),
.B(n_870),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1311),
.A2(n_1019),
.B1(n_1050),
.B2(n_1012),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1422),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1328),
.Y(n_1492)
);

NOR2x1_ASAP7_75t_L g1493 ( 
.A(n_1306),
.B(n_1069),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1397),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1306),
.B(n_830),
.Y(n_1495)
);

CKINVDCx8_ASAP7_75t_R g1496 ( 
.A(n_1352),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1305),
.Y(n_1497)
);

AND2x6_ASAP7_75t_L g1498 ( 
.A(n_1377),
.B(n_1052),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1335),
.B(n_939),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1416),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1329),
.B(n_830),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1437),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1333),
.B(n_1186),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1308),
.A2(n_1079),
.B1(n_1096),
.B2(n_1063),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1381),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1384),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1335),
.B(n_939),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1386),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1387),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1394),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1435),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1389),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1317),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1390),
.B(n_1393),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1302),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1319),
.B(n_866),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1336),
.B(n_1112),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1395),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1396),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1319),
.B(n_1348),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1304),
.Y(n_1521)
);

CKINVDCx6p67_ASAP7_75t_R g1522 ( 
.A(n_1404),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1398),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1401),
.A2(n_1073),
.B(n_1069),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1318),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1403),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1368),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1405),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1351),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1407),
.Y(n_1530)
);

INVx5_ASAP7_75t_L g1531 ( 
.A(n_1409),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1415),
.B(n_939),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1307),
.Y(n_1533)
);

OAI22x1_ASAP7_75t_L g1534 ( 
.A1(n_1326),
.A2(n_1155),
.B1(n_837),
.B2(n_859),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1410),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1309),
.B(n_866),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1367),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1310),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1411),
.Y(n_1539)
);

AND2x6_ASAP7_75t_L g1540 ( 
.A(n_1312),
.B(n_1073),
.Y(n_1540)
);

AOI22x1_ASAP7_75t_SL g1541 ( 
.A1(n_1317),
.A2(n_1187),
.B1(n_1188),
.B2(n_1114),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1368),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1412),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1413),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1414),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1314),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1419),
.B(n_1315),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1421),
.Y(n_1548)
);

AND2x6_ASAP7_75t_L g1549 ( 
.A(n_1316),
.B(n_1078),
.Y(n_1549)
);

CKINVDCx11_ASAP7_75t_R g1550 ( 
.A(n_1357),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1423),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1424),
.Y(n_1552)
);

OAI22x1_ASAP7_75t_SL g1553 ( 
.A1(n_1357),
.A2(n_1215),
.B1(n_1222),
.B2(n_1194),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1415),
.B(n_1075),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1425),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1426),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1427),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1428),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1429),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1320),
.Y(n_1560)
);

INVx6_ASAP7_75t_L g1561 ( 
.A(n_1321),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1430),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1514),
.B(n_1322),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1514),
.B(n_1327),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1345),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1446),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1515),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1446),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1445),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1546),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1469),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1562),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1562),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1453),
.B(n_1501),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1538),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1538),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1518),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1476),
.Y(n_1578)
);

BUFx8_ASAP7_75t_L g1579 ( 
.A(n_1525),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1453),
.B(n_1354),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1486),
.A2(n_1337),
.B(n_1330),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1487),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1476),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1519),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1469),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1510),
.B(n_862),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1523),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1530),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1449),
.Y(n_1589)
);

CKINVDCx11_ASAP7_75t_R g1590 ( 
.A(n_1550),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1449),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1481),
.B(n_1372),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1539),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1492),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1476),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1543),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1554),
.B(n_1345),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1479),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1544),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1445),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1479),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1545),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1492),
.B(n_1537),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1438),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1454),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1454),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1454),
.Y(n_1607)
);

OA21x2_ASAP7_75t_L g1608 ( 
.A1(n_1472),
.A2(n_1340),
.B(n_1339),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1479),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1548),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1551),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1552),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1555),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1556),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1472),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1473),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1473),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1447),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1558),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1559),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1521),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1501),
.B(n_1341),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1481),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1517),
.B(n_1343),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1481),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1471),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1537),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1547),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1482),
.B(n_1344),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1517),
.B(n_1346),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1521),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1533),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1506),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1506),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1506),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1533),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1483),
.A2(n_1356),
.B(n_1349),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1508),
.B(n_1358),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1509),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1509),
.B(n_1512),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1494),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1471),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1448),
.B(n_1360),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1560),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1495),
.B(n_1431),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1560),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1526),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1450),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1526),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1526),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1444),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1438),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1528),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1528),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1456),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1528),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1461),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1535),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1494),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1535),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1535),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1509),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1557),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1512),
.B(n_1372),
.Y(n_1664)
);

NAND2xp33_ASAP7_75t_SL g1665 ( 
.A(n_1527),
.B(n_1112),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1460),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1557),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1512),
.B(n_1383),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1464),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1557),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1463),
.B(n_1380),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1440),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1462),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_L g1674 ( 
.A(n_1475),
.B(n_866),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1452),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1542),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1489),
.B(n_1380),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1457),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1459),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1485),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1467),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1480),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1466),
.A2(n_1308),
.B1(n_1232),
.B2(n_1273),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1491),
.Y(n_1684)
);

BUFx8_ASAP7_75t_L g1685 ( 
.A(n_1502),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1511),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1524),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1462),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1495),
.B(n_1433),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1439),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1524),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1499),
.B(n_1331),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1439),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1561),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_SL g1695 ( 
.A(n_1500),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1561),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1561),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1465),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1668),
.B(n_1542),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1672),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1571),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1666),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1627),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1675),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1586),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1626),
.Y(n_1706)
);

INVx4_ASAP7_75t_L g1707 ( 
.A(n_1695),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1574),
.B(n_1488),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1586),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1683),
.A2(n_1503),
.B1(n_1466),
.B2(n_1498),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1579),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1678),
.Y(n_1712)
);

INVx4_ASAP7_75t_L g1713 ( 
.A(n_1695),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1579),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1574),
.B(n_1488),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1683),
.A2(n_1516),
.B1(n_1503),
.B2(n_1455),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1571),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1676),
.B(n_1500),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1585),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1681),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1604),
.B(n_1497),
.Y(n_1722)
);

AO22x2_ASAP7_75t_L g1723 ( 
.A1(n_1565),
.A2(n_1504),
.B1(n_1541),
.B2(n_1477),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1682),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1585),
.Y(n_1725)
);

OAI21xp33_ASAP7_75t_SL g1726 ( 
.A1(n_1668),
.A2(n_1516),
.B(n_1520),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1578),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1692),
.B(n_1527),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1627),
.B(n_1458),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1597),
.B(n_1603),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1604),
.B(n_1497),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1594),
.A2(n_1504),
.B1(n_1490),
.B2(n_1477),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1615),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1684),
.A2(n_1455),
.B1(n_1474),
.B2(n_1441),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1652),
.B(n_1529),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1594),
.B(n_1510),
.Y(n_1736)
);

INVx4_ASAP7_75t_L g1737 ( 
.A(n_1586),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1686),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1577),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1584),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1587),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1588),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1593),
.Y(n_1743)
);

BUFx10_ASAP7_75t_L g1744 ( 
.A(n_1622),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1596),
.Y(n_1745)
);

BUFx10_ASAP7_75t_L g1746 ( 
.A(n_1622),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1671),
.B(n_1547),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1651),
.B(n_1488),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1599),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1572),
.A2(n_1474),
.B1(n_1441),
.B2(n_1432),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1602),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1652),
.B(n_1687),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1626),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1642),
.Y(n_1754)
);

BUFx10_ASAP7_75t_L g1755 ( 
.A(n_1624),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1589),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1610),
.Y(n_1757)
);

NAND3xp33_ASAP7_75t_L g1758 ( 
.A(n_1563),
.B(n_1505),
.C(n_1485),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1691),
.B(n_1529),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1592),
.B(n_1510),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1642),
.Y(n_1761)
);

NAND2xp33_ASAP7_75t_L g1762 ( 
.A(n_1665),
.B(n_1488),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1624),
.B(n_1507),
.Y(n_1763)
);

NAND2xp33_ASAP7_75t_L g1764 ( 
.A(n_1665),
.B(n_1478),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1611),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1677),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1578),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1680),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1612),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1591),
.Y(n_1770)
);

INVx5_ASAP7_75t_L g1771 ( 
.A(n_1623),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1615),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1563),
.B(n_1505),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1564),
.B(n_1498),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_1641),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1616),
.Y(n_1776)
);

INVx5_ASAP7_75t_L g1777 ( 
.A(n_1623),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1616),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1613),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1614),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1680),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_L g1782 ( 
.A(n_1621),
.B(n_1478),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1659),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1617),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1619),
.Y(n_1785)
);

INVx5_ASAP7_75t_L g1786 ( 
.A(n_1623),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1617),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1651),
.B(n_1628),
.Y(n_1788)
);

INVx4_ASAP7_75t_SL g1789 ( 
.A(n_1630),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1620),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1573),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1625),
.Y(n_1792)
);

AO22x2_ASAP7_75t_L g1793 ( 
.A1(n_1645),
.A2(n_1490),
.B1(n_1553),
.B2(n_1388),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1564),
.B(n_1498),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1698),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_SL g1796 ( 
.A(n_1592),
.B(n_1520),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1630),
.B(n_1498),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1698),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1567),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1570),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1643),
.Y(n_1801)
);

AND2x6_ASAP7_75t_L g1802 ( 
.A(n_1645),
.B(n_1493),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1628),
.B(n_1522),
.Y(n_1803)
);

NAND2xp33_ASAP7_75t_L g1804 ( 
.A(n_1631),
.B(n_1478),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1664),
.B(n_1383),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1689),
.B(n_1332),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1608),
.A2(n_1432),
.B1(n_1478),
.B2(n_1540),
.Y(n_1807)
);

NOR3xp33_ASAP7_75t_SL g1808 ( 
.A(n_1664),
.B(n_787),
.C(n_786),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1580),
.Y(n_1809)
);

AND3x2_ASAP7_75t_L g1810 ( 
.A(n_1590),
.B(n_1470),
.C(n_1550),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1643),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1618),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1608),
.A2(n_1549),
.B1(n_1540),
.B2(n_1288),
.Y(n_1813)
);

BUFx4f_ASAP7_75t_L g1814 ( 
.A(n_1689),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1618),
.B(n_1487),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1580),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1648),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1575),
.B(n_1496),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1648),
.Y(n_1819)
);

CKINVDCx12_ASAP7_75t_R g1820 ( 
.A(n_1590),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1629),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1629),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_L g1823 ( 
.A(n_1632),
.B(n_794),
.C(n_833),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1685),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1655),
.Y(n_1825)
);

INVxp33_ASAP7_75t_L g1826 ( 
.A(n_1638),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1638),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1685),
.B(n_1338),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1655),
.A2(n_1549),
.B1(n_1540),
.B2(n_1293),
.Y(n_1829)
);

INVx4_ASAP7_75t_L g1830 ( 
.A(n_1625),
.Y(n_1830)
);

INVx5_ASAP7_75t_L g1831 ( 
.A(n_1625),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1657),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1568),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1636),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1634),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1644),
.Y(n_1836)
);

BUFx10_ASAP7_75t_L g1837 ( 
.A(n_1576),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1657),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_L g1839 ( 
.A(n_1646),
.B(n_1531),
.C(n_1536),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1669),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1634),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1694),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1669),
.Y(n_1843)
);

OR2x6_ASAP7_75t_L g1844 ( 
.A(n_1696),
.B(n_1534),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1569),
.Y(n_1845)
);

OAI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1600),
.A2(n_1229),
.B1(n_1347),
.B2(n_1342),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1637),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1673),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1566),
.Y(n_1849)
);

OAI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1647),
.A2(n_887),
.B1(n_924),
.B2(n_872),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1688),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1649),
.A2(n_1549),
.B1(n_1540),
.B2(n_988),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_L g1853 ( 
.A(n_1634),
.B(n_867),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1697),
.B(n_1484),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1650),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1578),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1653),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1583),
.Y(n_1858)
);

NAND2xp33_ASAP7_75t_L g1859 ( 
.A(n_1773),
.B(n_1639),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1770),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1702),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1727),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1821),
.B(n_1566),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1701),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1730),
.B(n_1359),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1775),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1814),
.B(n_1662),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1822),
.B(n_1654),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1747),
.B(n_1359),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1814),
.B(n_1639),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1699),
.B(n_1639),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1805),
.B(n_1662),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1827),
.B(n_1656),
.Y(n_1873)
);

O2A1O1Ixp33_ASAP7_75t_L g1874 ( 
.A1(n_1766),
.A2(n_1049),
.B(n_1145),
.C(n_983),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1801),
.B(n_1811),
.Y(n_1875)
);

NOR2xp67_ASAP7_75t_L g1876 ( 
.A(n_1758),
.B(n_1640),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1700),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1729),
.B(n_1417),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1732),
.A2(n_1417),
.B1(n_1388),
.B2(n_1658),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1756),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1704),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1773),
.B(n_1660),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1712),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1710),
.A2(n_1662),
.B1(n_787),
.B2(n_788),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1718),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1717),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1732),
.A2(n_1663),
.B1(n_1667),
.B2(n_1661),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1826),
.B(n_1721),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1736),
.B(n_1487),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1724),
.B(n_1670),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1720),
.Y(n_1891)
);

BUFx5_ASAP7_75t_L g1892 ( 
.A(n_1847),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1738),
.B(n_1633),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1708),
.B(n_1487),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1725),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_L g1896 ( 
.A(n_1727),
.Y(n_1896)
);

OAI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1710),
.A2(n_1184),
.B1(n_1179),
.B2(n_788),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1708),
.B(n_1583),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1726),
.A2(n_1674),
.B1(n_1549),
.B2(n_1640),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1739),
.Y(n_1900)
);

BUFx8_ASAP7_75t_L g1901 ( 
.A(n_1711),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1796),
.A2(n_1674),
.B1(n_1635),
.B2(n_1484),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1716),
.B(n_1583),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1733),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1737),
.B(n_1513),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1813),
.A2(n_1740),
.B1(n_1742),
.B2(n_1741),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1722),
.B(n_1595),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1743),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1783),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1745),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1703),
.B(n_1513),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1715),
.B(n_1595),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1715),
.B(n_1595),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1737),
.B(n_1385),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1749),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1772),
.Y(n_1916)
);

BUFx5_ASAP7_75t_L g1917 ( 
.A(n_1851),
.Y(n_1917)
);

INVx3_ASAP7_75t_L g1918 ( 
.A(n_1727),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1751),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1823),
.B(n_790),
.C(n_786),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1781),
.B(n_1598),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1722),
.B(n_1598),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1731),
.B(n_1598),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1776),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1731),
.B(n_1601),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1735),
.B(n_1601),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1735),
.B(n_1601),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1781),
.B(n_1763),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1763),
.B(n_1609),
.Y(n_1929)
);

INVx1_ASAP7_75t_SL g1930 ( 
.A(n_1806),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1753),
.B(n_1609),
.Y(n_1931)
);

BUFx12f_ASAP7_75t_SL g1932 ( 
.A(n_1707),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1757),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1778),
.Y(n_1934)
);

NOR3xp33_ASAP7_75t_L g1935 ( 
.A(n_1788),
.B(n_892),
.C(n_888),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1753),
.B(n_1754),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1765),
.B(n_1609),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1769),
.B(n_1779),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1784),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1780),
.B(n_1531),
.Y(n_1940)
);

NOR2x1p5_ASAP7_75t_L g1941 ( 
.A(n_1714),
.B(n_1470),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1785),
.B(n_1531),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1760),
.B(n_1605),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1790),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1754),
.B(n_1531),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1787),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1761),
.B(n_1606),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1761),
.B(n_1607),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1795),
.Y(n_1949)
);

INVx3_ASAP7_75t_L g1950 ( 
.A(n_1767),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1768),
.B(n_1536),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1723),
.A2(n_1088),
.B1(n_1231),
.B2(n_1075),
.Y(n_1952)
);

NAND2xp33_ASAP7_75t_L g1953 ( 
.A(n_1774),
.B(n_1690),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1798),
.Y(n_1954)
);

NOR3xp33_ASAP7_75t_L g1955 ( 
.A(n_1728),
.B(n_900),
.C(n_899),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1803),
.B(n_1436),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1768),
.B(n_1582),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1767),
.Y(n_1958)
);

AO221x1_ASAP7_75t_L g1959 ( 
.A1(n_1723),
.A2(n_1191),
.B1(n_1004),
.B2(n_906),
.C(n_895),
.Y(n_1959)
);

OAI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1726),
.A2(n_795),
.B1(n_796),
.B2(n_793),
.C(n_790),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1759),
.B(n_1582),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1759),
.B(n_1581),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1812),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1705),
.B(n_1295),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1829),
.A2(n_1088),
.B1(n_1231),
.B2(n_1075),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1706),
.B(n_1849),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1791),
.B(n_1581),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1744),
.B(n_1690),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1799),
.Y(n_1969)
);

INVx2_ASAP7_75t_SL g1970 ( 
.A(n_1744),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1746),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1809),
.B(n_1816),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1800),
.B(n_793),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1767),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1746),
.B(n_1690),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1755),
.B(n_1088),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1709),
.B(n_1299),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1817),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1802),
.A2(n_1231),
.B1(n_1122),
.B2(n_1156),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1819),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1755),
.B(n_1693),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1797),
.B(n_795),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1858),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1825),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1797),
.B(n_796),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1858),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1846),
.B(n_797),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1719),
.B(n_797),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1834),
.B(n_798),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1832),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1789),
.B(n_1693),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1789),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1838),
.Y(n_1993)
);

NAND2xp33_ASAP7_75t_L g1994 ( 
.A(n_1774),
.B(n_1693),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1840),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1858),
.Y(n_1996)
);

BUFx8_ASAP7_75t_L g1997 ( 
.A(n_1824),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1818),
.B(n_798),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1771),
.B(n_799),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1771),
.B(n_799),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1802),
.A2(n_885),
.B1(n_886),
.B2(n_884),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1833),
.B(n_1289),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1836),
.B(n_801),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1843),
.Y(n_2004)
);

INVxp67_ASAP7_75t_L g2005 ( 
.A(n_1802),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1848),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_SL g2007 ( 
.A(n_1707),
.B(n_1289),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1802),
.Y(n_2008)
);

INVxp67_ASAP7_75t_L g2009 ( 
.A(n_1854),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1713),
.B(n_1748),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1845),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1771),
.B(n_801),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1792),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1794),
.B(n_1855),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1794),
.B(n_805),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1857),
.B(n_805),
.Y(n_2016)
);

OAI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1713),
.A2(n_1758),
.B1(n_1850),
.B2(n_1842),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1828),
.B(n_806),
.Y(n_2018)
);

INVxp67_ASAP7_75t_L g2019 ( 
.A(n_1844),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1837),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1835),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1837),
.B(n_1295),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1750),
.A2(n_1752),
.B1(n_1841),
.B2(n_1835),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1777),
.B(n_806),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1752),
.B(n_808),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1792),
.B(n_808),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1841),
.B(n_1298),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1866),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1865),
.A2(n_1793),
.B1(n_1844),
.B2(n_1852),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1875),
.B(n_1762),
.Y(n_2030)
);

HB1xp67_ASAP7_75t_L g2031 ( 
.A(n_1861),
.Y(n_2031)
);

NOR3xp33_ASAP7_75t_SL g2032 ( 
.A(n_1880),
.B(n_811),
.C(n_810),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1998),
.B(n_1808),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1901),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1930),
.A2(n_1764),
.B1(n_1793),
.B2(n_1807),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_2009),
.B(n_1830),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1992),
.B(n_1777),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_2011),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1860),
.B(n_1777),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1877),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1888),
.B(n_1830),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1938),
.B(n_1786),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1881),
.Y(n_2043)
);

INVxp67_ASAP7_75t_SL g2044 ( 
.A(n_1966),
.Y(n_2044)
);

NAND2xp33_ASAP7_75t_L g2045 ( 
.A(n_1892),
.B(n_1786),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1909),
.B(n_1786),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1963),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1990),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1901),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1896),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1864),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1878),
.B(n_1844),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_2007),
.B(n_1831),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1885),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1911),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1883),
.Y(n_2056)
);

BUFx6f_ASAP7_75t_L g2057 ( 
.A(n_1896),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1886),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1891),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1869),
.B(n_1831),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1896),
.Y(n_2061)
);

BUFx2_ASAP7_75t_L g2062 ( 
.A(n_1997),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1906),
.B(n_1831),
.Y(n_2063)
);

CKINVDCx20_ASAP7_75t_R g2064 ( 
.A(n_1932),
.Y(n_2064)
);

AND2x6_ASAP7_75t_L g2065 ( 
.A(n_2013),
.B(n_1815),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_2017),
.B(n_1956),
.Y(n_2066)
);

AOI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1987),
.A2(n_1804),
.B1(n_1782),
.B2(n_1856),
.Y(n_2067)
);

CKINVDCx20_ASAP7_75t_R g2068 ( 
.A(n_1997),
.Y(n_2068)
);

INVx6_ASAP7_75t_L g2069 ( 
.A(n_1941),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1900),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1962),
.A2(n_1815),
.B(n_1839),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1897),
.B(n_1839),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_1905),
.Y(n_2073)
);

BUFx4f_ASAP7_75t_L g2074 ( 
.A(n_1970),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1895),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1958),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1908),
.B(n_1734),
.Y(n_2077)
);

OR2x6_ASAP7_75t_L g2078 ( 
.A(n_1971),
.B(n_1810),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1958),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1910),
.B(n_1915),
.Y(n_2080)
);

BUFx10_ASAP7_75t_L g2081 ( 
.A(n_2022),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1919),
.B(n_810),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1933),
.Y(n_2083)
);

AND2x2_ASAP7_75t_SL g2084 ( 
.A(n_1952),
.B(n_1820),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1879),
.A2(n_1965),
.B1(n_1960),
.B2(n_1959),
.Y(n_2085)
);

OR2x6_ASAP7_75t_L g2086 ( 
.A(n_2019),
.B(n_1078),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_1914),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_2005),
.B(n_811),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1904),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1916),
.Y(n_2090)
);

BUFx2_ASAP7_75t_L g2091 ( 
.A(n_1976),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1944),
.B(n_812),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1924),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_R g2094 ( 
.A(n_2020),
.B(n_1853),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1887),
.B(n_812),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_2010),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1972),
.Y(n_2097)
);

INVx2_ASAP7_75t_SL g2098 ( 
.A(n_1999),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1969),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2025),
.B(n_815),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1988),
.A2(n_891),
.B1(n_893),
.B2(n_890),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1978),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2027),
.B(n_815),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1934),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_2008),
.B(n_819),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1882),
.B(n_819),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1980),
.Y(n_2107)
);

NOR2x2_ASAP7_75t_L g2108 ( 
.A(n_2001),
.B(n_1122),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_1958),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1863),
.B(n_820),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1868),
.B(n_820),
.Y(n_2111)
);

NAND2x1p5_ASAP7_75t_L g2112 ( 
.A(n_1928),
.B(n_1465),
.Y(n_2112)
);

A2O1A1Ixp33_ASAP7_75t_L g2113 ( 
.A1(n_1876),
.A2(n_1159),
.B(n_1163),
.C(n_1156),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1902),
.B(n_821),
.Y(n_2114)
);

BUFx4f_ASAP7_75t_L g2115 ( 
.A(n_1974),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_2013),
.B(n_821),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1984),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1873),
.B(n_822),
.Y(n_2118)
);

BUFx3_ASAP7_75t_L g2119 ( 
.A(n_1974),
.Y(n_2119)
);

NOR2x1p5_ASAP7_75t_L g2120 ( 
.A(n_2018),
.B(n_1291),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2002),
.A2(n_1977),
.B1(n_1964),
.B2(n_1884),
.Y(n_2121)
);

NAND2x2_ASAP7_75t_L g2122 ( 
.A(n_1989),
.B(n_822),
.Y(n_2122)
);

NOR2xp67_ASAP7_75t_L g2123 ( 
.A(n_2026),
.B(n_824),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1943),
.B(n_824),
.Y(n_2124)
);

BUFx3_ASAP7_75t_L g2125 ( 
.A(n_1974),
.Y(n_2125)
);

AOI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_1929),
.A2(n_1898),
.B1(n_1913),
.B2(n_1912),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_2000),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1979),
.B(n_826),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_1935),
.A2(n_896),
.B1(n_903),
.B2(n_894),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_1983),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1993),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_1973),
.B(n_826),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_2012),
.Y(n_2133)
);

OR2x6_ASAP7_75t_L g2134 ( 
.A(n_1991),
.B(n_1159),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1995),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2014),
.B(n_828),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1982),
.B(n_828),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1983),
.B(n_829),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1983),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1985),
.B(n_2015),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1890),
.B(n_829),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1862),
.B(n_901),
.Y(n_2142)
);

INVxp67_ASAP7_75t_L g2143 ( 
.A(n_2003),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_2024),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_2006),
.A2(n_832),
.B1(n_834),
.B2(n_831),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2016),
.B(n_831),
.Y(n_2146)
);

AOI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_2004),
.A2(n_834),
.B1(n_835),
.B2(n_832),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1874),
.B(n_835),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1862),
.B(n_1287),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1986),
.B(n_836),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1893),
.B(n_836),
.Y(n_2151)
);

NOR3xp33_ASAP7_75t_SL g2152 ( 
.A(n_1920),
.B(n_840),
.C(n_839),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1937),
.B(n_839),
.Y(n_2153)
);

BUFx8_ASAP7_75t_SL g2154 ( 
.A(n_1986),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1939),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1955),
.B(n_840),
.Y(n_2156)
);

INVx2_ASAP7_75t_SL g2157 ( 
.A(n_1986),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1946),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1949),
.B(n_841),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1954),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_1918),
.B(n_841),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_1918),
.Y(n_2162)
);

AOI22xp33_ASAP7_75t_L g2163 ( 
.A1(n_1917),
.A2(n_846),
.B1(n_850),
.B2(n_843),
.Y(n_2163)
);

INVx3_ASAP7_75t_L g2164 ( 
.A(n_1950),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1951),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1907),
.B(n_843),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2021),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_SL g2168 ( 
.A(n_1917),
.B(n_1950),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_SL g2169 ( 
.A(n_1876),
.B(n_846),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1917),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1917),
.B(n_850),
.Y(n_2171)
);

AOI22xp5_ASAP7_75t_L g2172 ( 
.A1(n_1867),
.A2(n_905),
.B1(n_910),
.B2(n_904),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1917),
.Y(n_2173)
);

BUFx4f_ASAP7_75t_L g2174 ( 
.A(n_1996),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1996),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1870),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1921),
.Y(n_2177)
);

NAND2xp33_ASAP7_75t_SL g2178 ( 
.A(n_2033),
.B(n_1936),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2096),
.B(n_1872),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_2121),
.B(n_2023),
.Y(n_2180)
);

NAND2xp33_ASAP7_75t_SL g2181 ( 
.A(n_2064),
.B(n_852),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_2169),
.B(n_1922),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_2036),
.B(n_1923),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2044),
.B(n_2066),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2055),
.B(n_852),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_2030),
.B(n_1925),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_2073),
.B(n_1926),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2081),
.B(n_2115),
.Y(n_2188)
);

NAND2xp33_ASAP7_75t_SL g2189 ( 
.A(n_2152),
.B(n_854),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_2081),
.B(n_1927),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_2115),
.B(n_1871),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2165),
.B(n_1968),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_2042),
.B(n_1899),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_2060),
.B(n_1899),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_2072),
.B(n_1961),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2052),
.B(n_2097),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_SL g2197 ( 
.A(n_2176),
.B(n_1892),
.Y(n_2197)
);

NAND2xp33_ASAP7_75t_SL g2198 ( 
.A(n_2103),
.B(n_854),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2159),
.B(n_858),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_SL g2200 ( 
.A(n_2176),
.B(n_2041),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_2176),
.B(n_2074),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2143),
.B(n_1975),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_2074),
.B(n_1892),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_2175),
.B(n_1892),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_2091),
.B(n_1892),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_2050),
.B(n_1947),
.Y(n_2206)
);

NAND2xp33_ASAP7_75t_SL g2207 ( 
.A(n_2068),
.B(n_858),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2031),
.B(n_1981),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_2050),
.B(n_1948),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_2162),
.B(n_2037),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_2037),
.B(n_1894),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_2050),
.B(n_1957),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_2057),
.B(n_1889),
.Y(n_2213)
);

NAND2xp33_ASAP7_75t_SL g2214 ( 
.A(n_2032),
.B(n_860),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2080),
.B(n_860),
.Y(n_2215)
);

NAND2xp33_ASAP7_75t_SL g2216 ( 
.A(n_2140),
.B(n_861),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_2057),
.B(n_1931),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_2057),
.B(n_1945),
.Y(n_2218)
);

NAND2xp33_ASAP7_75t_SL g2219 ( 
.A(n_2087),
.B(n_2094),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_2061),
.B(n_1940),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_2061),
.B(n_1942),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2132),
.B(n_861),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_2061),
.B(n_1903),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_2076),
.B(n_1967),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_2076),
.B(n_863),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_2076),
.B(n_863),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2136),
.B(n_864),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2040),
.B(n_864),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2148),
.B(n_1062),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_SL g2230 ( 
.A(n_2139),
.B(n_2085),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2043),
.B(n_1062),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2056),
.B(n_1065),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2058),
.B(n_1065),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_2139),
.B(n_1298),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2070),
.B(n_2083),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_2139),
.B(n_1299),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_2067),
.B(n_1221),
.Y(n_2237)
);

NAND2xp33_ASAP7_75t_SL g2238 ( 
.A(n_2062),
.B(n_1221),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_2164),
.B(n_1224),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_2164),
.B(n_1224),
.Y(n_2240)
);

NAND2xp33_ASAP7_75t_SL g2241 ( 
.A(n_2100),
.B(n_1226),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2084),
.B(n_1226),
.Y(n_2242)
);

NAND2xp33_ASAP7_75t_SL g2243 ( 
.A(n_2137),
.B(n_1227),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2099),
.B(n_1227),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2174),
.B(n_1228),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_2079),
.B(n_1228),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2079),
.B(n_1230),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2124),
.B(n_1230),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_2130),
.B(n_1234),
.Y(n_2249)
);

NAND2xp33_ASAP7_75t_SL g2250 ( 
.A(n_2146),
.B(n_1234),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_2130),
.B(n_1237),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_2157),
.B(n_1237),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_2063),
.B(n_1238),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_2035),
.B(n_1238),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2126),
.B(n_1240),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2177),
.B(n_1240),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2177),
.B(n_1243),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2106),
.B(n_1243),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2177),
.B(n_1285),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2053),
.B(n_1285),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_2142),
.B(n_1286),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2142),
.B(n_1286),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2149),
.B(n_1290),
.Y(n_2263)
);

NAND2xp33_ASAP7_75t_L g2264 ( 
.A(n_2065),
.B(n_1244),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2149),
.B(n_1290),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2111),
.B(n_2118),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2119),
.B(n_1291),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2141),
.B(n_1244),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2125),
.B(n_1245),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_2123),
.B(n_2098),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2120),
.B(n_1245),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2038),
.B(n_2095),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2127),
.B(n_1246),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2133),
.B(n_1246),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2029),
.B(n_1247),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_2144),
.B(n_1247),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2161),
.B(n_2086),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2109),
.B(n_1251),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2114),
.B(n_1251),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2151),
.B(n_2166),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2028),
.B(n_1253),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_2170),
.B(n_1253),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_2134),
.B(n_1468),
.Y(n_2283)
);

NAND2xp33_ASAP7_75t_SL g2284 ( 
.A(n_2163),
.B(n_1254),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_2173),
.B(n_1254),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2086),
.B(n_2101),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2039),
.B(n_1260),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2082),
.B(n_1260),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2046),
.B(n_1261),
.Y(n_2289)
);

NAND2xp33_ASAP7_75t_SL g2290 ( 
.A(n_2092),
.B(n_1261),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2167),
.B(n_1262),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2088),
.B(n_1262),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2145),
.B(n_1266),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2105),
.B(n_1266),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2077),
.B(n_1268),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2153),
.B(n_1268),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2171),
.B(n_2112),
.Y(n_2297)
);

NAND2xp33_ASAP7_75t_SL g2298 ( 
.A(n_2110),
.B(n_1269),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2102),
.B(n_1281),
.Y(n_2299)
);

NAND2xp33_ASAP7_75t_SL g2300 ( 
.A(n_2116),
.B(n_1269),
.Y(n_2300)
);

NAND2xp33_ASAP7_75t_SL g2301 ( 
.A(n_2138),
.B(n_1271),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2147),
.B(n_1271),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2107),
.B(n_1272),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2117),
.B(n_1283),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_2131),
.B(n_1283),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2135),
.B(n_1272),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_SL g2307 ( 
.A(n_2150),
.B(n_1274),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2168),
.B(n_1274),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2156),
.B(n_1275),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2129),
.B(n_1275),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_2113),
.B(n_1276),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2047),
.B(n_1276),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2048),
.B(n_1277),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2051),
.B(n_1277),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2155),
.B(n_1279),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2134),
.B(n_1468),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_2054),
.B(n_2090),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_2059),
.B(n_1279),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2158),
.B(n_2160),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2075),
.B(n_2089),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_2093),
.B(n_1280),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2071),
.B(n_1859),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2104),
.B(n_1280),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2128),
.B(n_867),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2172),
.B(n_1281),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2049),
.B(n_1284),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2045),
.B(n_867),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_2065),
.B(n_867),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2154),
.B(n_1284),
.Y(n_2329)
);

AOI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2180),
.A2(n_2078),
.B1(n_2034),
.B2(n_911),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2319),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2229),
.B(n_2078),
.Y(n_2332)
);

NAND2x1_ASAP7_75t_L g2333 ( 
.A(n_2184),
.B(n_2065),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2266),
.B(n_908),
.Y(n_2334)
);

HB1xp67_ASAP7_75t_L g2335 ( 
.A(n_2235),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_2210),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_2219),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2280),
.B(n_923),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2272),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2196),
.B(n_927),
.Y(n_2340)
);

BUFx6f_ASAP7_75t_L g2341 ( 
.A(n_2210),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2317),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2255),
.A2(n_2122),
.B1(n_2069),
.B2(n_933),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2199),
.B(n_931),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2195),
.B(n_2108),
.Y(n_2345)
);

AND3x1_ASAP7_75t_SL g2346 ( 
.A(n_2207),
.B(n_1294),
.C(n_1278),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2187),
.B(n_912),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2254),
.A2(n_2065),
.B1(n_1233),
.B2(n_1282),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2277),
.B(n_2286),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_2181),
.Y(n_2350)
);

CKINVDCx8_ASAP7_75t_R g2351 ( 
.A(n_2211),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2320),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2192),
.Y(n_2353)
);

NAND2x1_ASAP7_75t_L g2354 ( 
.A(n_2211),
.B(n_2069),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2185),
.B(n_1296),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2208),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2200),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2242),
.B(n_934),
.Y(n_2358)
);

AND3x1_ASAP7_75t_SL g2359 ( 
.A(n_2238),
.B(n_940),
.C(n_935),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2223),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2215),
.B(n_942),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2201),
.B(n_950),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2186),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2179),
.B(n_954),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_2329),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2190),
.B(n_913),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2271),
.B(n_955),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2206),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2202),
.B(n_958),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2275),
.B(n_959),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2270),
.Y(n_2371)
);

AND2x2_ASAP7_75t_SL g2372 ( 
.A(n_2264),
.B(n_2293),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2283),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2302),
.B(n_2222),
.Y(n_2374)
);

BUFx8_ASAP7_75t_L g2375 ( 
.A(n_2283),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2183),
.B(n_960),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2261),
.B(n_1259),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2228),
.B(n_965),
.Y(n_2378)
);

INVxp67_ASAP7_75t_L g2379 ( 
.A(n_2273),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2209),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2224),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2231),
.B(n_970),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2262),
.B(n_1270),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2205),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2194),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2232),
.B(n_977),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2188),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2212),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2193),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2316),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2316),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2263),
.B(n_979),
.Y(n_2392)
);

AOI21xp5_ASAP7_75t_L g2393 ( 
.A1(n_2322),
.A2(n_1994),
.B(n_1953),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2284),
.A2(n_916),
.B1(n_918),
.B2(n_915),
.Y(n_2394)
);

NAND2x1p5_ASAP7_75t_L g2395 ( 
.A(n_2203),
.B(n_984),
.Y(n_2395)
);

AOI22xp33_ASAP7_75t_L g2396 ( 
.A1(n_2216),
.A2(n_1233),
.B1(n_1282),
.B2(n_1163),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2233),
.B(n_986),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2182),
.B(n_919),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_R g2399 ( 
.A(n_2290),
.B(n_780),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_2323),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2265),
.B(n_1256),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2244),
.B(n_992),
.Y(n_2402)
);

AND3x1_ASAP7_75t_SL g2403 ( 
.A(n_2214),
.B(n_1265),
.C(n_1258),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2303),
.B(n_997),
.Y(n_2404)
);

INVx3_ASAP7_75t_L g2405 ( 
.A(n_2315),
.Y(n_2405)
);

NAND2x1p5_ASAP7_75t_L g2406 ( 
.A(n_2191),
.B(n_999),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2218),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2306),
.B(n_1000),
.Y(n_2408)
);

OAI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2292),
.A2(n_1003),
.B1(n_1009),
.B2(n_1002),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2230),
.A2(n_1020),
.B1(n_1021),
.B2(n_1017),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2326),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2281),
.Y(n_2412)
);

OAI22xp5_ASAP7_75t_SL g2413 ( 
.A1(n_2248),
.A2(n_1032),
.B1(n_1033),
.B2(n_1029),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2295),
.B(n_1034),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2178),
.B(n_1035),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2227),
.B(n_1041),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2217),
.Y(n_2417)
);

BUFx8_ASAP7_75t_L g2418 ( 
.A(n_2245),
.Y(n_2418)
);

INVx3_ASAP7_75t_L g2419 ( 
.A(n_2197),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2258),
.B(n_1046),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2288),
.B(n_1054),
.Y(n_2421)
);

BUFx4f_ASAP7_75t_SL g2422 ( 
.A(n_2267),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2268),
.B(n_2253),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2220),
.Y(n_2424)
);

INVxp67_ASAP7_75t_SL g2425 ( 
.A(n_2327),
.Y(n_2425)
);

AND3x1_ASAP7_75t_SL g2426 ( 
.A(n_2198),
.B(n_1064),
.C(n_1055),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2204),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2299),
.B(n_1071),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2256),
.B(n_1080),
.Y(n_2429)
);

INVx1_ASAP7_75t_SL g2430 ( 
.A(n_2269),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2324),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2221),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2304),
.B(n_1094),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_L g2434 ( 
.A(n_2213),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2294),
.B(n_920),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2257),
.B(n_1097),
.Y(n_2436)
);

BUFx2_ASAP7_75t_L g2437 ( 
.A(n_2301),
.Y(n_2437)
);

OAI22xp5_ASAP7_75t_SL g2438 ( 
.A1(n_2250),
.A2(n_1110),
.B1(n_1116),
.B2(n_1101),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2324),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2259),
.B(n_1118),
.Y(n_2440)
);

BUFx6f_ASAP7_75t_L g2441 ( 
.A(n_2328),
.Y(n_2441)
);

BUFx2_ASAP7_75t_L g2442 ( 
.A(n_2307),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_2328),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2327),
.Y(n_2444)
);

NAND2x1p5_ASAP7_75t_L g2445 ( 
.A(n_2297),
.B(n_1132),
.Y(n_2445)
);

INVx1_ASAP7_75t_SL g2446 ( 
.A(n_2274),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2322),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2276),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2312),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2305),
.B(n_1133),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2313),
.Y(n_2451)
);

OAI22xp5_ASAP7_75t_SL g2452 ( 
.A1(n_2241),
.A2(n_1257),
.B1(n_1255),
.B2(n_1138),
.Y(n_2452)
);

BUFx6f_ASAP7_75t_L g2453 ( 
.A(n_2260),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_2189),
.Y(n_2454)
);

BUFx2_ASAP7_75t_L g2455 ( 
.A(n_2300),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2237),
.B(n_921),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_2298),
.B(n_922),
.Y(n_2457)
);

INVx1_ASAP7_75t_SL g2458 ( 
.A(n_2278),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2243),
.B(n_2225),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2291),
.B(n_1135),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2314),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2296),
.B(n_2226),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2318),
.Y(n_2463)
);

AOI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2310),
.A2(n_926),
.B1(n_928),
.B2(n_925),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2309),
.B(n_1223),
.Y(n_2465)
);

BUFx6f_ASAP7_75t_L g2466 ( 
.A(n_2287),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2234),
.B(n_1140),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2321),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2282),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2285),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2236),
.B(n_1142),
.Y(n_2471)
);

INVx2_ASAP7_75t_SL g2472 ( 
.A(n_2336),
.Y(n_2472)
);

BUFx10_ASAP7_75t_L g2473 ( 
.A(n_2350),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2405),
.B(n_2345),
.Y(n_2474)
);

INVx8_ASAP7_75t_L g2475 ( 
.A(n_2336),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2335),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2331),
.Y(n_2477)
);

OR2x2_ASAP7_75t_L g2478 ( 
.A(n_2356),
.B(n_2252),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2336),
.B(n_2246),
.Y(n_2479)
);

OR2x2_ASAP7_75t_L g2480 ( 
.A(n_2349),
.B(n_2247),
.Y(n_2480)
);

OAI21x1_ASAP7_75t_L g2481 ( 
.A1(n_2393),
.A2(n_2311),
.B(n_2308),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2353),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_2341),
.Y(n_2483)
);

INVx4_ASAP7_75t_L g2484 ( 
.A(n_2387),
.Y(n_2484)
);

AOI21x1_ASAP7_75t_L g2485 ( 
.A1(n_2333),
.A2(n_2251),
.B(n_2249),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2363),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_L g2487 ( 
.A1(n_2431),
.A2(n_2240),
.B(n_2239),
.Y(n_2487)
);

OAI21x1_ASAP7_75t_L g2488 ( 
.A1(n_2439),
.A2(n_2289),
.B(n_2279),
.Y(n_2488)
);

AOI21x1_ASAP7_75t_L g2489 ( 
.A1(n_2415),
.A2(n_2325),
.B(n_1146),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2342),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2339),
.Y(n_2491)
);

OAI21x1_ASAP7_75t_L g2492 ( 
.A1(n_2447),
.A2(n_1148),
.B(n_1144),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2365),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2360),
.Y(n_2494)
);

INVx1_ASAP7_75t_SL g2495 ( 
.A(n_2385),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2381),
.Y(n_2496)
);

AOI22x1_ASAP7_75t_L g2497 ( 
.A1(n_2337),
.A2(n_932),
.B1(n_936),
.B2(n_930),
.Y(n_2497)
);

OAI21x1_ASAP7_75t_L g2498 ( 
.A1(n_2389),
.A2(n_1151),
.B(n_1149),
.Y(n_2498)
);

NAND2x1p5_ASAP7_75t_L g2499 ( 
.A(n_2441),
.B(n_867),
.Y(n_2499)
);

INVxp67_ASAP7_75t_SL g2500 ( 
.A(n_2443),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2352),
.Y(n_2501)
);

BUFx3_ASAP7_75t_L g2502 ( 
.A(n_2354),
.Y(n_2502)
);

OR2x2_ASAP7_75t_L g2503 ( 
.A(n_2340),
.B(n_1152),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_SL g2504 ( 
.A(n_2372),
.B(n_1157),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2341),
.B(n_895),
.Y(n_2505)
);

BUFx3_ASAP7_75t_L g2506 ( 
.A(n_2375),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2341),
.B(n_895),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2357),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_SL g2509 ( 
.A(n_2351),
.B(n_1158),
.Y(n_2509)
);

BUFx3_ASAP7_75t_L g2510 ( 
.A(n_2375),
.Y(n_2510)
);

OAI21x1_ASAP7_75t_L g2511 ( 
.A1(n_2419),
.A2(n_1168),
.B(n_1162),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2384),
.B(n_2368),
.Y(n_2512)
);

AO21x2_ASAP7_75t_L g2513 ( 
.A1(n_2425),
.A2(n_1235),
.B(n_1225),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2417),
.Y(n_2514)
);

OAI21x1_ASAP7_75t_L g2515 ( 
.A1(n_2419),
.A2(n_1181),
.B(n_1177),
.Y(n_2515)
);

INVx1_ASAP7_75t_SL g2516 ( 
.A(n_2444),
.Y(n_2516)
);

INVx6_ASAP7_75t_L g2517 ( 
.A(n_2418),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2407),
.Y(n_2518)
);

NAND2x1p5_ASAP7_75t_L g2519 ( 
.A(n_2441),
.B(n_895),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2424),
.Y(n_2520)
);

OA21x2_ASAP7_75t_L g2521 ( 
.A1(n_2380),
.A2(n_1195),
.B(n_1183),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2388),
.Y(n_2522)
);

AO21x2_ASAP7_75t_L g2523 ( 
.A1(n_2432),
.A2(n_1252),
.B(n_1250),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2434),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2427),
.Y(n_2525)
);

OAI21xp5_ASAP7_75t_L g2526 ( 
.A1(n_2394),
.A2(n_1202),
.B(n_1198),
.Y(n_2526)
);

BUFx3_ASAP7_75t_L g2527 ( 
.A(n_2418),
.Y(n_2527)
);

AOI22x1_ASAP7_75t_L g2528 ( 
.A1(n_2454),
.A2(n_938),
.B1(n_941),
.B2(n_937),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2434),
.Y(n_2529)
);

OAI21xp5_ASAP7_75t_L g2530 ( 
.A1(n_2394),
.A2(n_1209),
.B(n_1205),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2434),
.Y(n_2531)
);

OAI21x1_ASAP7_75t_L g2532 ( 
.A1(n_2427),
.A2(n_1210),
.B(n_1216),
.Y(n_2532)
);

AO21x2_ASAP7_75t_L g2533 ( 
.A1(n_2376),
.A2(n_1241),
.B(n_1236),
.Y(n_2533)
);

AND2x4_ASAP7_75t_L g2534 ( 
.A(n_2373),
.B(n_895),
.Y(n_2534)
);

NAND2xp33_ASAP7_75t_L g2535 ( 
.A(n_2399),
.B(n_906),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2374),
.B(n_1248),
.Y(n_2536)
);

INVx3_ASAP7_75t_SL g2537 ( 
.A(n_2412),
.Y(n_2537)
);

OA21x2_ASAP7_75t_L g2538 ( 
.A1(n_2390),
.A2(n_945),
.B(n_944),
.Y(n_2538)
);

AO21x2_ASAP7_75t_L g2539 ( 
.A1(n_2370),
.A2(n_1199),
.B(n_1439),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2441),
.Y(n_2540)
);

BUFx4_ASAP7_75t_SL g2541 ( 
.A(n_2411),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2400),
.Y(n_2542)
);

AOI21xp5_ASAP7_75t_L g2543 ( 
.A1(n_2444),
.A2(n_1004),
.B(n_906),
.Y(n_2543)
);

AOI22x1_ASAP7_75t_L g2544 ( 
.A1(n_2455),
.A2(n_947),
.B1(n_949),
.B2(n_948),
.Y(n_2544)
);

OAI21x1_ASAP7_75t_SL g2545 ( 
.A1(n_2330),
.A2(n_1),
.B(n_3),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2400),
.Y(n_2546)
);

BUFx3_ASAP7_75t_L g2547 ( 
.A(n_2391),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2405),
.Y(n_2548)
);

NAND2x1p5_ASAP7_75t_L g2549 ( 
.A(n_2444),
.B(n_906),
.Y(n_2549)
);

OAI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2334),
.A2(n_952),
.B(n_951),
.Y(n_2550)
);

BUFx3_ASAP7_75t_L g2551 ( 
.A(n_2453),
.Y(n_2551)
);

AOI21x1_ASAP7_75t_L g2552 ( 
.A1(n_2369),
.A2(n_1443),
.B(n_1442),
.Y(n_2552)
);

BUFx2_ASAP7_75t_L g2553 ( 
.A(n_2371),
.Y(n_2553)
);

INVx2_ASAP7_75t_SL g2554 ( 
.A(n_2453),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2422),
.Y(n_2555)
);

OAI21x1_ASAP7_75t_SL g2556 ( 
.A1(n_2330),
.A2(n_1),
.B(n_4),
.Y(n_2556)
);

AO21x2_ASAP7_75t_L g2557 ( 
.A1(n_2398),
.A2(n_1443),
.B(n_1442),
.Y(n_2557)
);

OAI21x1_ASAP7_75t_L g2558 ( 
.A1(n_2395),
.A2(n_1443),
.B(n_1442),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2451),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2469),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_2332),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2453),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2461),
.Y(n_2563)
);

AOI22x1_ASAP7_75t_L g2564 ( 
.A1(n_2437),
.A2(n_953),
.B1(n_957),
.B2(n_956),
.Y(n_2564)
);

INVx4_ASAP7_75t_L g2565 ( 
.A(n_2466),
.Y(n_2565)
);

OAI21x1_ASAP7_75t_L g2566 ( 
.A1(n_2470),
.A2(n_1451),
.B(n_781),
.Y(n_2566)
);

OR2x2_ASAP7_75t_L g2567 ( 
.A(n_2364),
.B(n_2344),
.Y(n_2567)
);

INVx2_ASAP7_75t_SL g2568 ( 
.A(n_2466),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2468),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2449),
.Y(n_2570)
);

BUFx3_ASAP7_75t_L g2571 ( 
.A(n_2466),
.Y(n_2571)
);

NAND2x1p5_ASAP7_75t_L g2572 ( 
.A(n_2362),
.B(n_2442),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2355),
.B(n_2367),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2512),
.Y(n_2574)
);

BUFx3_ASAP7_75t_L g2575 ( 
.A(n_2555),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2512),
.Y(n_2576)
);

INVx4_ASAP7_75t_L g2577 ( 
.A(n_2517),
.Y(n_2577)
);

BUFx2_ASAP7_75t_L g2578 ( 
.A(n_2553),
.Y(n_2578)
);

BUFx6f_ASAP7_75t_L g2579 ( 
.A(n_2562),
.Y(n_2579)
);

BUFx12f_ASAP7_75t_L g2580 ( 
.A(n_2493),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2504),
.A2(n_2413),
.B1(n_2452),
.B2(n_2404),
.Y(n_2581)
);

INVx1_ASAP7_75t_SL g2582 ( 
.A(n_2495),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2490),
.Y(n_2583)
);

BUFx12f_ASAP7_75t_L g2584 ( 
.A(n_2493),
.Y(n_2584)
);

BUFx2_ASAP7_75t_L g2585 ( 
.A(n_2548),
.Y(n_2585)
);

CKINVDCx11_ASAP7_75t_R g2586 ( 
.A(n_2537),
.Y(n_2586)
);

AOI22xp33_ASAP7_75t_L g2587 ( 
.A1(n_2504),
.A2(n_2452),
.B1(n_2421),
.B2(n_2377),
.Y(n_2587)
);

BUFx2_ASAP7_75t_SL g2588 ( 
.A(n_2527),
.Y(n_2588)
);

BUFx3_ASAP7_75t_L g2589 ( 
.A(n_2506),
.Y(n_2589)
);

AOI22xp33_ASAP7_75t_L g2590 ( 
.A1(n_2573),
.A2(n_2383),
.B1(n_2401),
.B2(n_2392),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2561),
.B(n_2430),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2486),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2560),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2561),
.B(n_2446),
.Y(n_2594)
);

CKINVDCx11_ASAP7_75t_R g2595 ( 
.A(n_2537),
.Y(n_2595)
);

OAI22xp33_ASAP7_75t_L g2596 ( 
.A1(n_2509),
.A2(n_2445),
.B1(n_2458),
.B2(n_2406),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2514),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2501),
.Y(n_2598)
);

OAI22xp33_ASAP7_75t_SL g2599 ( 
.A1(n_2509),
.A2(n_2338),
.B1(n_2361),
.B2(n_2459),
.Y(n_2599)
);

BUFx12f_ASAP7_75t_L g2600 ( 
.A(n_2517),
.Y(n_2600)
);

OAI21xp5_ASAP7_75t_L g2601 ( 
.A1(n_2535),
.A2(n_2410),
.B(n_2396),
.Y(n_2601)
);

BUFx3_ASAP7_75t_L g2602 ( 
.A(n_2510),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2535),
.A2(n_2463),
.B1(n_2433),
.B2(n_2428),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2525),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2562),
.Y(n_2605)
);

OAI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2526),
.A2(n_2464),
.B1(n_2423),
.B2(n_2420),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2476),
.B(n_2379),
.Y(n_2607)
);

INVx6_ASAP7_75t_L g2608 ( 
.A(n_2473),
.Y(n_2608)
);

OAI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2572),
.A2(n_2448),
.B1(n_2464),
.B2(n_2462),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2526),
.A2(n_2438),
.B1(n_2348),
.B2(n_2416),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2538),
.A2(n_2465),
.B1(n_2362),
.B2(n_2343),
.Y(n_2611)
);

CKINVDCx6p67_ASAP7_75t_R g2612 ( 
.A(n_2473),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2495),
.B(n_2542),
.Y(n_2613)
);

CKINVDCx11_ASAP7_75t_R g2614 ( 
.A(n_2484),
.Y(n_2614)
);

INVx6_ASAP7_75t_L g2615 ( 
.A(n_2562),
.Y(n_2615)
);

INVx3_ASAP7_75t_L g2616 ( 
.A(n_2525),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2571),
.Y(n_2617)
);

INVx1_ASAP7_75t_SL g2618 ( 
.A(n_2551),
.Y(n_2618)
);

INVxp67_ASAP7_75t_SL g2619 ( 
.A(n_2500),
.Y(n_2619)
);

INVx2_ASAP7_75t_SL g2620 ( 
.A(n_2551),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2520),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2494),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2482),
.B(n_2378),
.Y(n_2623)
);

BUFx6f_ASAP7_75t_L g2624 ( 
.A(n_2531),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_L g2625 ( 
.A1(n_2538),
.A2(n_2414),
.B1(n_2386),
.B2(n_2397),
.Y(n_2625)
);

BUFx8_ASAP7_75t_SL g2626 ( 
.A(n_2531),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_SL g2627 ( 
.A1(n_2533),
.A2(n_2435),
.B1(n_2409),
.B2(n_2402),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2546),
.B(n_2382),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2496),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2539),
.A2(n_2408),
.B1(n_2358),
.B2(n_2456),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2539),
.A2(n_2440),
.B1(n_2429),
.B2(n_2436),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2518),
.Y(n_2632)
);

INVx8_ASAP7_75t_L g2633 ( 
.A(n_2475),
.Y(n_2633)
);

OAI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2572),
.A2(n_2471),
.B1(n_2467),
.B2(n_2450),
.Y(n_2634)
);

CKINVDCx11_ASAP7_75t_R g2635 ( 
.A(n_2484),
.Y(n_2635)
);

CKINVDCx6p67_ASAP7_75t_R g2636 ( 
.A(n_2541),
.Y(n_2636)
);

INVx4_ASAP7_75t_L g2637 ( 
.A(n_2517),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2522),
.Y(n_2638)
);

OAI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2567),
.A2(n_2460),
.B1(n_2359),
.B2(n_2347),
.Y(n_2639)
);

INVx5_ASAP7_75t_L g2640 ( 
.A(n_2531),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2508),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2491),
.Y(n_2642)
);

AOI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2474),
.A2(n_2426),
.B1(n_2346),
.B2(n_2403),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2559),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2563),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2569),
.Y(n_2646)
);

AOI22xp33_ASAP7_75t_SL g2647 ( 
.A1(n_2533),
.A2(n_1214),
.B1(n_961),
.B2(n_963),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2502),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2477),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2570),
.A2(n_2366),
.B1(n_2457),
.B2(n_1004),
.Y(n_2650)
);

BUFx10_ASAP7_75t_L g2651 ( 
.A(n_2479),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2582),
.Y(n_2652)
);

AOI21xp5_ASAP7_75t_L g2653 ( 
.A1(n_2606),
.A2(n_2543),
.B(n_2500),
.Y(n_2653)
);

OA21x2_ASAP7_75t_L g2654 ( 
.A1(n_2619),
.A2(n_2576),
.B(n_2574),
.Y(n_2654)
);

AOI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2606),
.A2(n_2543),
.B(n_2474),
.Y(n_2655)
);

AOI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2619),
.A2(n_2530),
.B(n_2557),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2648),
.B(n_2565),
.Y(n_2657)
);

AOI21xp5_ASAP7_75t_L g2658 ( 
.A1(n_2609),
.A2(n_2530),
.B(n_2557),
.Y(n_2658)
);

OAI21x1_ASAP7_75t_L g2659 ( 
.A1(n_2623),
.A2(n_2552),
.B(n_2566),
.Y(n_2659)
);

INVx1_ASAP7_75t_SL g2660 ( 
.A(n_2582),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2586),
.Y(n_2661)
);

OAI21x1_ASAP7_75t_L g2662 ( 
.A1(n_2623),
.A2(n_2540),
.B(n_2631),
.Y(n_2662)
);

AOI22xp33_ASAP7_75t_L g2663 ( 
.A1(n_2627),
.A2(n_2513),
.B1(n_2523),
.B2(n_2521),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2578),
.B(n_2536),
.Y(n_2664)
);

NAND2x1_ASAP7_75t_L g2665 ( 
.A(n_2604),
.B(n_2565),
.Y(n_2665)
);

OAI21x1_ASAP7_75t_L g2666 ( 
.A1(n_2604),
.A2(n_2540),
.B(n_2521),
.Y(n_2666)
);

AOI21xp5_ASAP7_75t_L g2667 ( 
.A1(n_2639),
.A2(n_2599),
.B(n_2610),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2613),
.B(n_2478),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2608),
.B(n_2503),
.Y(n_2669)
);

AO21x2_ASAP7_75t_L g2670 ( 
.A1(n_2634),
.A2(n_2529),
.B(n_2524),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2592),
.Y(n_2671)
);

A2O1A1Ixp33_ASAP7_75t_L g2672 ( 
.A1(n_2627),
.A2(n_2550),
.B(n_2480),
.C(n_2479),
.Y(n_2672)
);

OA21x2_ASAP7_75t_L g2673 ( 
.A1(n_2622),
.A2(n_2487),
.B(n_2488),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2598),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2610),
.A2(n_2513),
.B1(n_2523),
.B2(n_2547),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2628),
.B(n_2568),
.Y(n_2676)
);

OAI21xp33_ASAP7_75t_L g2677 ( 
.A1(n_2599),
.A2(n_2550),
.B(n_1191),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2629),
.B(n_2554),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2632),
.Y(n_2679)
);

HB1xp67_ASAP7_75t_L g2680 ( 
.A(n_2585),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2581),
.A2(n_2547),
.B1(n_2556),
.B2(n_2545),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2641),
.Y(n_2682)
);

CKINVDCx20_ASAP7_75t_R g2683 ( 
.A(n_2595),
.Y(n_2683)
);

BUFx2_ASAP7_75t_L g2684 ( 
.A(n_2626),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2638),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2644),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2643),
.A2(n_2485),
.B1(n_2564),
.B2(n_2544),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2645),
.B(n_2516),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2607),
.Y(n_2689)
);

AOI21xp5_ASAP7_75t_L g2690 ( 
.A1(n_2601),
.A2(n_2558),
.B(n_2481),
.Y(n_2690)
);

AO31x2_ASAP7_75t_L g2691 ( 
.A1(n_2583),
.A2(n_2516),
.A3(n_2534),
.B(n_2549),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2646),
.Y(n_2692)
);

CKINVDCx16_ASAP7_75t_R g2693 ( 
.A(n_2580),
.Y(n_2693)
);

OAI21x1_ASAP7_75t_L g2694 ( 
.A1(n_2616),
.A2(n_2499),
.B(n_2519),
.Y(n_2694)
);

AOI21xp5_ASAP7_75t_L g2695 ( 
.A1(n_2601),
.A2(n_2492),
.B(n_2499),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2642),
.B(n_2618),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2649),
.Y(n_2697)
);

AO21x2_ASAP7_75t_L g2698 ( 
.A1(n_2596),
.A2(n_2534),
.B(n_2489),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_SL g2699 ( 
.A1(n_2594),
.A2(n_2591),
.B1(n_2648),
.B2(n_2651),
.Y(n_2699)
);

A2O1A1Ixp33_ASAP7_75t_L g2700 ( 
.A1(n_2647),
.A2(n_2498),
.B(n_2532),
.C(n_2515),
.Y(n_2700)
);

CKINVDCx14_ASAP7_75t_R g2701 ( 
.A(n_2636),
.Y(n_2701)
);

AOI221xp5_ASAP7_75t_L g2702 ( 
.A1(n_2625),
.A2(n_964),
.B1(n_967),
.B2(n_966),
.C(n_962),
.Y(n_2702)
);

OR2x6_ASAP7_75t_L g2703 ( 
.A(n_2620),
.B(n_2475),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2593),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2618),
.B(n_2505),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2616),
.B(n_2472),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2643),
.A2(n_2519),
.B1(n_2549),
.B2(n_2483),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2597),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2617),
.B(n_2648),
.Y(n_2709)
);

A2O1A1Ixp33_ASAP7_75t_L g2710 ( 
.A1(n_2647),
.A2(n_2511),
.B(n_2507),
.C(n_2505),
.Y(n_2710)
);

AOI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2640),
.A2(n_2475),
.B(n_2507),
.Y(n_2711)
);

AOI21xp5_ASAP7_75t_L g2712 ( 
.A1(n_2640),
.A2(n_2497),
.B(n_2528),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2587),
.A2(n_1004),
.B1(n_1061),
.B2(n_906),
.Y(n_2713)
);

OAI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2630),
.A2(n_969),
.B(n_968),
.Y(n_2714)
);

AOI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2640),
.A2(n_1061),
.B(n_1004),
.Y(n_2715)
);

AO31x2_ASAP7_75t_L g2716 ( 
.A1(n_2621),
.A2(n_1161),
.A3(n_1191),
.B(n_1061),
.Y(n_2716)
);

AOI221xp5_ASAP7_75t_L g2717 ( 
.A1(n_2611),
.A2(n_973),
.B1(n_975),
.B2(n_972),
.C(n_971),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2651),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2579),
.B(n_1061),
.Y(n_2719)
);

AO21x2_ASAP7_75t_L g2720 ( 
.A1(n_2603),
.A2(n_2541),
.B(n_1161),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_SL g2721 ( 
.A1(n_2577),
.A2(n_1161),
.B1(n_1191),
.B2(n_1061),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2579),
.B(n_2605),
.Y(n_2722)
);

AOI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_2633),
.A2(n_1191),
.B(n_1161),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2671),
.Y(n_2724)
);

HB1xp67_ASAP7_75t_L g2725 ( 
.A(n_2654),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_2677),
.A2(n_2590),
.B1(n_2650),
.B2(n_2608),
.Y(n_2726)
);

OAI211xp5_ASAP7_75t_L g2727 ( 
.A1(n_2667),
.A2(n_2614),
.B(n_2635),
.C(n_2577),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2689),
.B(n_2637),
.Y(n_2728)
);

OAI211xp5_ASAP7_75t_L g2729 ( 
.A1(n_2677),
.A2(n_2637),
.B(n_2602),
.C(n_2589),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2673),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2680),
.B(n_2588),
.Y(n_2731)
);

A2O1A1Ixp33_ASAP7_75t_L g2732 ( 
.A1(n_2672),
.A2(n_2575),
.B(n_978),
.C(n_980),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_L g2733 ( 
.A1(n_2675),
.A2(n_2615),
.B1(n_2605),
.B2(n_2579),
.Y(n_2733)
);

AOI22xp33_ASAP7_75t_L g2734 ( 
.A1(n_2663),
.A2(n_2615),
.B1(n_2624),
.B2(n_2605),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2673),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2660),
.B(n_2612),
.Y(n_2736)
);

AOI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2720),
.A2(n_2624),
.B1(n_2600),
.B2(n_1264),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2655),
.A2(n_2633),
.B1(n_2624),
.B2(n_2584),
.Y(n_2738)
);

OAI22xp33_ASAP7_75t_L g2739 ( 
.A1(n_2653),
.A2(n_2633),
.B1(n_1264),
.B2(n_1161),
.Y(n_2739)
);

AOI22xp33_ASAP7_75t_L g2740 ( 
.A1(n_2720),
.A2(n_1264),
.B1(n_1220),
.B2(n_981),
.Y(n_2740)
);

INVxp67_ASAP7_75t_SL g2741 ( 
.A(n_2654),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2674),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2698),
.A2(n_1264),
.B1(n_1300),
.B2(n_982),
.Y(n_2743)
);

AND2x6_ASAP7_75t_L g2744 ( 
.A(n_2660),
.B(n_1264),
.Y(n_2744)
);

OAI211xp5_ASAP7_75t_SL g2745 ( 
.A1(n_2664),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_2745)
);

AOI22xp33_ASAP7_75t_L g2746 ( 
.A1(n_2698),
.A2(n_1213),
.B1(n_1200),
.B2(n_985),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_SL g2747 ( 
.A1(n_2670),
.A2(n_1005),
.B1(n_1024),
.B2(n_976),
.Y(n_2747)
);

AOI221xp5_ASAP7_75t_L g2748 ( 
.A1(n_2702),
.A2(n_990),
.B1(n_993),
.B2(n_989),
.C(n_987),
.Y(n_2748)
);

OAI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2681),
.A2(n_998),
.B1(n_1001),
.B2(n_995),
.Y(n_2749)
);

OAI21xp33_ASAP7_75t_L g2750 ( 
.A1(n_2696),
.A2(n_1013),
.B(n_1008),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2714),
.A2(n_1015),
.B1(n_1018),
.B2(n_1014),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_2717),
.A2(n_1023),
.B1(n_1026),
.B2(n_1022),
.Y(n_2752)
);

AOI22xp33_ASAP7_75t_L g2753 ( 
.A1(n_2658),
.A2(n_2670),
.B1(n_2687),
.B2(n_2713),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_L g2754 ( 
.A(n_2693),
.B(n_6),
.Y(n_2754)
);

OAI21xp5_ASAP7_75t_SL g2755 ( 
.A1(n_2701),
.A2(n_7),
.B(n_9),
.Y(n_2755)
);

BUFx2_ASAP7_75t_L g2756 ( 
.A(n_2652),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2706),
.B(n_9),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2668),
.B(n_1028),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2718),
.B(n_10),
.Y(n_2759)
);

INVxp67_ASAP7_75t_L g2760 ( 
.A(n_2669),
.Y(n_2760)
);

OAI22xp33_ASAP7_75t_L g2761 ( 
.A1(n_2656),
.A2(n_1031),
.B1(n_1036),
.B2(n_1030),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2684),
.Y(n_2762)
);

AOI22xp33_ASAP7_75t_L g2763 ( 
.A1(n_2695),
.A2(n_1039),
.B1(n_1040),
.B2(n_1038),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2690),
.A2(n_1043),
.B(n_1042),
.Y(n_2764)
);

AOI22xp5_ASAP7_75t_L g2765 ( 
.A1(n_2707),
.A2(n_1045),
.B1(n_1047),
.B2(n_1044),
.Y(n_2765)
);

AOI221xp5_ASAP7_75t_L g2766 ( 
.A1(n_2697),
.A2(n_1053),
.B1(n_1056),
.B2(n_1051),
.C(n_1048),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2724),
.Y(n_2767)
);

HB1xp67_ASAP7_75t_L g2768 ( 
.A(n_2756),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2730),
.Y(n_2769)
);

INVx3_ASAP7_75t_L g2770 ( 
.A(n_2735),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2728),
.B(n_2709),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2725),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2725),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2741),
.B(n_2662),
.Y(n_2774)
);

INVx3_ASAP7_75t_L g2775 ( 
.A(n_2762),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2741),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_2736),
.B(n_2703),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2742),
.Y(n_2778)
);

AND2x4_ASAP7_75t_L g2779 ( 
.A(n_2731),
.B(n_2703),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2760),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2757),
.B(n_2703),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2755),
.B(n_2661),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2744),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2761),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2744),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2744),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2759),
.B(n_2679),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2744),
.Y(n_2788)
);

BUFx2_ASAP7_75t_L g2789 ( 
.A(n_2738),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2744),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2727),
.B(n_2685),
.Y(n_2791)
);

NAND4xp25_ASAP7_75t_L g2792 ( 
.A(n_2753),
.B(n_2692),
.C(n_2678),
.D(n_2723),
.Y(n_2792)
);

AND2x4_ASAP7_75t_L g2793 ( 
.A(n_2734),
.B(n_2666),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2754),
.B(n_2699),
.Y(n_2794)
);

BUFx2_ASAP7_75t_L g2795 ( 
.A(n_2758),
.Y(n_2795)
);

BUFx6f_ASAP7_75t_L g2796 ( 
.A(n_2747),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2750),
.B(n_2683),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2761),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2733),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2729),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2746),
.A2(n_2682),
.B1(n_2686),
.B2(n_2704),
.Y(n_2801)
);

INVx1_ASAP7_75t_SL g2802 ( 
.A(n_2765),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2789),
.B(n_2665),
.Y(n_2803)
);

O2A1O1Ixp33_ASAP7_75t_L g2804 ( 
.A1(n_2784),
.A2(n_2732),
.B(n_2745),
.C(n_2739),
.Y(n_2804)
);

AOI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2789),
.A2(n_2739),
.B(n_2764),
.Y(n_2805)
);

AO21x2_ASAP7_75t_L g2806 ( 
.A1(n_2776),
.A2(n_2749),
.B(n_2719),
.Y(n_2806)
);

AOI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2800),
.A2(n_2743),
.B(n_2763),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2773),
.Y(n_2808)
);

CKINVDCx6p67_ASAP7_75t_R g2809 ( 
.A(n_2796),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2780),
.B(n_2763),
.Y(n_2810)
);

HB1xp67_ASAP7_75t_L g2811 ( 
.A(n_2768),
.Y(n_2811)
);

OA21x2_ASAP7_75t_L g2812 ( 
.A1(n_2776),
.A2(n_2740),
.B(n_2737),
.Y(n_2812)
);

AO21x2_ASAP7_75t_L g2813 ( 
.A1(n_2772),
.A2(n_2715),
.B(n_2659),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2767),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2800),
.A2(n_2657),
.B(n_2726),
.Y(n_2815)
);

AO31x2_ASAP7_75t_L g2816 ( 
.A1(n_2773),
.A2(n_2710),
.A3(n_2700),
.B(n_2708),
.Y(n_2816)
);

A2O1A1Ixp33_ASAP7_75t_L g2817 ( 
.A1(n_2784),
.A2(n_2751),
.B(n_2712),
.C(n_2766),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_L g2818 ( 
.A1(n_2799),
.A2(n_2751),
.B1(n_2676),
.B2(n_2752),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2777),
.B(n_2722),
.Y(n_2819)
);

OR2x2_ASAP7_75t_L g2820 ( 
.A(n_2780),
.B(n_2688),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2769),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2769),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2767),
.Y(n_2823)
);

HB1xp67_ASAP7_75t_L g2824 ( 
.A(n_2795),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2769),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_2795),
.Y(n_2826)
);

INVx4_ASAP7_75t_L g2827 ( 
.A(n_2775),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2777),
.B(n_2705),
.Y(n_2828)
);

BUFx2_ASAP7_75t_L g2829 ( 
.A(n_2777),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2770),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2772),
.Y(n_2831)
);

OAI21xp33_ASAP7_75t_L g2832 ( 
.A1(n_2792),
.A2(n_2798),
.B(n_2774),
.Y(n_2832)
);

O2A1O1Ixp5_ASAP7_75t_L g2833 ( 
.A1(n_2793),
.A2(n_2711),
.B(n_2721),
.C(n_2752),
.Y(n_2833)
);

AOI22xp33_ASAP7_75t_SL g2834 ( 
.A1(n_2794),
.A2(n_2694),
.B1(n_1059),
.B2(n_1060),
.Y(n_2834)
);

AO21x2_ASAP7_75t_L g2835 ( 
.A1(n_2774),
.A2(n_2716),
.B(n_2748),
.Y(n_2835)
);

INVx3_ASAP7_75t_L g2836 ( 
.A(n_2774),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2798),
.B(n_2716),
.Y(n_2837)
);

OAI21x1_ASAP7_75t_L g2838 ( 
.A1(n_2770),
.A2(n_2716),
.B(n_2691),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2787),
.Y(n_2839)
);

HB1xp67_ASAP7_75t_L g2840 ( 
.A(n_2775),
.Y(n_2840)
);

INVxp67_ASAP7_75t_SL g2841 ( 
.A(n_2775),
.Y(n_2841)
);

OR2x2_ASAP7_75t_L g2842 ( 
.A(n_2824),
.B(n_2770),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2826),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2814),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2826),
.Y(n_2845)
);

BUFx2_ASAP7_75t_L g2846 ( 
.A(n_2829),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2803),
.B(n_2777),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2814),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2803),
.B(n_2779),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2806),
.Y(n_2850)
);

NOR2xp33_ASAP7_75t_L g2851 ( 
.A(n_2810),
.B(n_2782),
.Y(n_2851)
);

NAND4xp25_ASAP7_75t_L g2852 ( 
.A(n_2832),
.B(n_2797),
.C(n_2791),
.D(n_2794),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2829),
.B(n_2779),
.Y(n_2853)
);

BUFx2_ASAP7_75t_L g2854 ( 
.A(n_2841),
.Y(n_2854)
);

OAI211xp5_ASAP7_75t_SL g2855 ( 
.A1(n_2807),
.A2(n_2802),
.B(n_2799),
.C(n_2783),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2831),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2831),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2819),
.B(n_2779),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2823),
.Y(n_2859)
);

INVx2_ASAP7_75t_SL g2860 ( 
.A(n_2836),
.Y(n_2860)
);

INVx3_ASAP7_75t_L g2861 ( 
.A(n_2836),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2839),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2806),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2819),
.B(n_2779),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2839),
.B(n_2791),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2811),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2827),
.B(n_2781),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2808),
.Y(n_2868)
);

AO21x2_ASAP7_75t_L g2869 ( 
.A1(n_2805),
.A2(n_2774),
.B(n_2783),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2806),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_2840),
.Y(n_2871)
);

OR2x2_ASAP7_75t_L g2872 ( 
.A(n_2808),
.B(n_2787),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2838),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2815),
.B(n_2785),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2827),
.B(n_2781),
.Y(n_2875)
);

OA332x1_ASAP7_75t_L g2876 ( 
.A1(n_2827),
.A2(n_2771),
.A3(n_2796),
.B1(n_2793),
.B2(n_16),
.B3(n_12),
.C1(n_15),
.C2(n_14),
.Y(n_2876)
);

AOI33xp33_ASAP7_75t_L g2877 ( 
.A1(n_2818),
.A2(n_2793),
.A3(n_2801),
.B1(n_2786),
.B2(n_2785),
.B3(n_2790),
.Y(n_2877)
);

INVxp67_ASAP7_75t_SL g2878 ( 
.A(n_2854),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2844),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2847),
.B(n_2820),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2847),
.B(n_2820),
.Y(n_2881)
);

OR2x2_ASAP7_75t_L g2882 ( 
.A(n_2872),
.B(n_2837),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2849),
.B(n_2853),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_SL g2884 ( 
.A(n_2851),
.B(n_2833),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2846),
.B(n_2817),
.Y(n_2885)
);

OR2x2_ASAP7_75t_L g2886 ( 
.A(n_2872),
.B(n_2828),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2846),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2849),
.B(n_2771),
.Y(n_2888)
);

OR2x2_ASAP7_75t_L g2889 ( 
.A(n_2866),
.B(n_2828),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2844),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2859),
.B(n_2835),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2856),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2853),
.Y(n_2893)
);

INVx4_ASAP7_75t_L g2894 ( 
.A(n_2843),
.Y(n_2894)
);

NAND2x1p5_ASAP7_75t_L g2895 ( 
.A(n_2854),
.B(n_2843),
.Y(n_2895)
);

AND2x2_ASAP7_75t_SL g2896 ( 
.A(n_2877),
.B(n_2812),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2845),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2867),
.B(n_2836),
.Y(n_2898)
);

AND2x4_ASAP7_75t_L g2899 ( 
.A(n_2845),
.B(n_2830),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2852),
.B(n_2821),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2856),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2857),
.Y(n_2902)
);

INVx3_ASAP7_75t_L g2903 ( 
.A(n_2861),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2867),
.B(n_2821),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2875),
.B(n_2822),
.Y(n_2905)
);

AND2x4_ASAP7_75t_L g2906 ( 
.A(n_2875),
.B(n_2822),
.Y(n_2906)
);

O2A1O1Ixp33_ASAP7_75t_L g2907 ( 
.A1(n_2855),
.A2(n_2804),
.B(n_2835),
.C(n_2812),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2860),
.B(n_2825),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2861),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2857),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2848),
.Y(n_2911)
);

AND2x4_ASAP7_75t_SL g2912 ( 
.A(n_2858),
.B(n_2809),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2858),
.B(n_2825),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2862),
.B(n_2835),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2868),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2868),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2860),
.B(n_2830),
.Y(n_2917)
);

AND2x4_ASAP7_75t_L g2918 ( 
.A(n_2864),
.B(n_2786),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2861),
.Y(n_2919)
);

OR2x2_ASAP7_75t_L g2920 ( 
.A(n_2865),
.B(n_2812),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2864),
.B(n_2788),
.Y(n_2921)
);

OR2x2_ASAP7_75t_L g2922 ( 
.A(n_2865),
.B(n_2813),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2871),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2842),
.Y(n_2924)
);

INVxp67_ASAP7_75t_L g2925 ( 
.A(n_2897),
.Y(n_2925)
);

INVxp67_ASAP7_75t_SL g2926 ( 
.A(n_2885),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2878),
.B(n_2869),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2878),
.B(n_2896),
.Y(n_2928)
);

NOR3xp33_ASAP7_75t_L g2929 ( 
.A(n_2884),
.B(n_2874),
.C(n_2834),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2879),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2893),
.B(n_2869),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_L g2932 ( 
.A(n_2894),
.B(n_2869),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2885),
.Y(n_2933)
);

OR2x2_ASAP7_75t_L g2934 ( 
.A(n_2886),
.B(n_2842),
.Y(n_2934)
);

NAND4xp75_ASAP7_75t_SL g2935 ( 
.A(n_2883),
.B(n_2876),
.C(n_2809),
.D(n_2813),
.Y(n_2935)
);

INVxp67_ASAP7_75t_SL g2936 ( 
.A(n_2895),
.Y(n_2936)
);

AND2x2_ASAP7_75t_L g2937 ( 
.A(n_2888),
.B(n_2788),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2895),
.Y(n_2938)
);

OAI31xp33_ASAP7_75t_L g2939 ( 
.A1(n_2884),
.A2(n_2876),
.A3(n_2863),
.B(n_2870),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2896),
.B(n_2850),
.Y(n_2940)
);

NAND4xp75_ASAP7_75t_L g2941 ( 
.A(n_2891),
.B(n_2863),
.C(n_2870),
.D(n_2850),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2880),
.B(n_2873),
.Y(n_2942)
);

INVxp67_ASAP7_75t_SL g2943 ( 
.A(n_2903),
.Y(n_2943)
);

BUFx2_ASAP7_75t_L g2944 ( 
.A(n_2894),
.Y(n_2944)
);

NAND4xp75_ASAP7_75t_L g2945 ( 
.A(n_2891),
.B(n_2873),
.C(n_2790),
.D(n_2796),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2890),
.Y(n_2946)
);

XOR2x1_ASAP7_75t_L g2947 ( 
.A(n_2887),
.B(n_2796),
.Y(n_2947)
);

BUFx2_ASAP7_75t_L g2948 ( 
.A(n_2899),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2881),
.B(n_2813),
.Y(n_2949)
);

NOR4xp75_ASAP7_75t_L g2950 ( 
.A(n_2908),
.B(n_2796),
.C(n_2816),
.D(n_12),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2920),
.B(n_2816),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2892),
.Y(n_2952)
);

XNOR2xp5_ASAP7_75t_L g2953 ( 
.A(n_2912),
.B(n_2838),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_2912),
.Y(n_2954)
);

NAND3xp33_ASAP7_75t_SL g2955 ( 
.A(n_2907),
.B(n_2922),
.C(n_2900),
.Y(n_2955)
);

HB1xp67_ASAP7_75t_L g2956 ( 
.A(n_2919),
.Y(n_2956)
);

XNOR2xp5_ASAP7_75t_L g2957 ( 
.A(n_2918),
.B(n_2778),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2924),
.B(n_2816),
.Y(n_2958)
);

NAND4xp75_ASAP7_75t_L g2959 ( 
.A(n_2908),
.B(n_2816),
.C(n_2778),
.D(n_13),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2899),
.B(n_2816),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2901),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2902),
.Y(n_2962)
);

BUFx2_ASAP7_75t_L g2963 ( 
.A(n_2898),
.Y(n_2963)
);

INVxp67_ASAP7_75t_SL g2964 ( 
.A(n_2903),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2910),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2913),
.B(n_10),
.Y(n_2966)
);

INVx4_ASAP7_75t_L g2967 ( 
.A(n_2909),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2915),
.Y(n_2968)
);

XNOR2x2_ASAP7_75t_L g2969 ( 
.A(n_2923),
.B(n_11),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2916),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2904),
.B(n_14),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2911),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2882),
.Y(n_2973)
);

NOR3xp33_ASAP7_75t_SL g2974 ( 
.A(n_2917),
.B(n_1197),
.C(n_1196),
.Y(n_2974)
);

INVx3_ASAP7_75t_L g2975 ( 
.A(n_2909),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2889),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2905),
.B(n_16),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2921),
.Y(n_2978)
);

NAND4xp75_ASAP7_75t_SL g2979 ( 
.A(n_2917),
.B(n_19),
.C(n_17),
.D(n_18),
.Y(n_2979)
);

XNOR2x2_ASAP7_75t_L g2980 ( 
.A(n_2914),
.B(n_2907),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2914),
.Y(n_2981)
);

INVx2_ASAP7_75t_SL g2982 ( 
.A(n_2918),
.Y(n_2982)
);

NAND4xp75_ASAP7_75t_SL g2983 ( 
.A(n_2906),
.B(n_21),
.C(n_17),
.D(n_20),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2906),
.Y(n_2984)
);

NAND4xp75_ASAP7_75t_L g2985 ( 
.A(n_2896),
.B(n_22),
.C(n_20),
.D(n_21),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2883),
.B(n_22),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2894),
.B(n_1057),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2878),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2878),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2883),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2883),
.Y(n_2991)
);

AOI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2955),
.A2(n_1068),
.B1(n_1070),
.B2(n_1067),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2928),
.Y(n_2993)
);

BUFx2_ASAP7_75t_L g2994 ( 
.A(n_2948),
.Y(n_2994)
);

NOR5xp2_ASAP7_75t_L g2995 ( 
.A(n_2925),
.B(n_26),
.C(n_23),
.D(n_25),
.E(n_28),
.Y(n_2995)
);

INVx3_ASAP7_75t_SL g2996 ( 
.A(n_2986),
.Y(n_2996)
);

HB1xp67_ASAP7_75t_L g2997 ( 
.A(n_2963),
.Y(n_2997)
);

INVxp67_ASAP7_75t_SL g2998 ( 
.A(n_2928),
.Y(n_2998)
);

NAND2x1p5_ASAP7_75t_L g2999 ( 
.A(n_2971),
.B(n_2977),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2954),
.B(n_1072),
.Y(n_3000)
);

AOI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2929),
.A2(n_1076),
.B1(n_1077),
.B2(n_1074),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2988),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2954),
.B(n_1081),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_2990),
.B(n_1083),
.Y(n_3004)
);

AND2x4_ASAP7_75t_L g3005 ( 
.A(n_2982),
.B(n_26),
.Y(n_3005)
);

OAI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2926),
.A2(n_1087),
.B1(n_1089),
.B2(n_1086),
.Y(n_3006)
);

AOI221xp5_ASAP7_75t_L g3007 ( 
.A1(n_2940),
.A2(n_1093),
.B1(n_1095),
.B2(n_1092),
.C(n_1091),
.Y(n_3007)
);

OR2x6_ASAP7_75t_L g3008 ( 
.A(n_2985),
.B(n_28),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2966),
.B(n_1098),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2989),
.Y(n_3010)
);

OR2x2_ASAP7_75t_L g3011 ( 
.A(n_2934),
.B(n_29),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2947),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2940),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2980),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2944),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2927),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2991),
.B(n_1100),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2927),
.Y(n_3018)
);

AND2x2_ASAP7_75t_L g3019 ( 
.A(n_2936),
.B(n_1103),
.Y(n_3019)
);

AOI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2959),
.A2(n_1106),
.B1(n_1107),
.B2(n_1104),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2975),
.Y(n_3021)
);

OR2x2_ASAP7_75t_L g3022 ( 
.A(n_2976),
.B(n_29),
.Y(n_3022)
);

OR2x2_ASAP7_75t_L g3023 ( 
.A(n_2973),
.B(n_2978),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2937),
.B(n_1108),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2956),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2939),
.B(n_1109),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2984),
.B(n_30),
.Y(n_3027)
);

OR2x2_ASAP7_75t_L g3028 ( 
.A(n_2942),
.B(n_30),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2933),
.A2(n_1113),
.B1(n_1119),
.B2(n_1111),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2938),
.B(n_1120),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2930),
.Y(n_3031)
);

AOI32xp33_ASAP7_75t_L g3032 ( 
.A1(n_2932),
.A2(n_1124),
.A3(n_1125),
.B1(n_1123),
.B2(n_1121),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2946),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2931),
.B(n_32),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2952),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2975),
.Y(n_3036)
);

BUFx2_ASAP7_75t_L g3037 ( 
.A(n_2943),
.Y(n_3037)
);

NOR2x1_ASAP7_75t_L g3038 ( 
.A(n_2967),
.B(n_32),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2939),
.B(n_1127),
.Y(n_3039)
);

BUFx2_ASAP7_75t_L g3040 ( 
.A(n_2964),
.Y(n_3040)
);

OR2x2_ASAP7_75t_L g3041 ( 
.A(n_2969),
.B(n_33),
.Y(n_3041)
);

INVxp67_ASAP7_75t_SL g3042 ( 
.A(n_2987),
.Y(n_3042)
);

NOR2xp67_ASAP7_75t_SL g3043 ( 
.A(n_2945),
.B(n_1129),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2957),
.B(n_1130),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2961),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2962),
.Y(n_3046)
);

OR2x2_ASAP7_75t_L g3047 ( 
.A(n_2949),
.B(n_33),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2974),
.B(n_1131),
.Y(n_3048)
);

AOI211xp5_ASAP7_75t_L g3049 ( 
.A1(n_2953),
.A2(n_1136),
.B(n_1137),
.C(n_1134),
.Y(n_3049)
);

INVx1_ASAP7_75t_SL g3050 ( 
.A(n_2983),
.Y(n_3050)
);

NAND3xp33_ASAP7_75t_SL g3051 ( 
.A(n_2950),
.B(n_1141),
.C(n_1139),
.Y(n_3051)
);

NAND2x1_ASAP7_75t_L g3052 ( 
.A(n_2967),
.B(n_34),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2941),
.Y(n_3053)
);

NAND2x1p5_ASAP7_75t_L g3054 ( 
.A(n_2972),
.B(n_38),
.Y(n_3054)
);

NAND2x1p5_ASAP7_75t_L g3055 ( 
.A(n_2968),
.B(n_39),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2970),
.B(n_1143),
.Y(n_3056)
);

AOI211xp5_ASAP7_75t_L g3057 ( 
.A1(n_2958),
.A2(n_1150),
.B(n_1154),
.C(n_1147),
.Y(n_3057)
);

OAI21xp5_ASAP7_75t_L g3058 ( 
.A1(n_2951),
.A2(n_1164),
.B(n_1160),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2965),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2981),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_L g3061 ( 
.A(n_2960),
.B(n_1165),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2935),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2979),
.Y(n_3063)
);

INVxp67_ASAP7_75t_L g3064 ( 
.A(n_2950),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_2928),
.B(n_36),
.Y(n_3065)
);

OR2x2_ASAP7_75t_L g3066 ( 
.A(n_2928),
.B(n_39),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2986),
.B(n_1166),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2948),
.Y(n_3068)
);

OAI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_2928),
.A2(n_1170),
.B1(n_1171),
.B2(n_1167),
.Y(n_3069)
);

BUFx2_ASAP7_75t_L g3070 ( 
.A(n_2948),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2948),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2939),
.B(n_1172),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2986),
.B(n_1173),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2986),
.B(n_1174),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2948),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2986),
.B(n_1176),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2948),
.Y(n_3077)
);

OAI221xp5_ASAP7_75t_SL g3078 ( 
.A1(n_2928),
.A2(n_1182),
.B1(n_1185),
.B2(n_1180),
.C(n_1178),
.Y(n_3078)
);

INVxp67_ASAP7_75t_L g3079 ( 
.A(n_2948),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2948),
.Y(n_3080)
);

CKINVDCx16_ASAP7_75t_R g3081 ( 
.A(n_2986),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2928),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2986),
.B(n_1189),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2928),
.Y(n_3084)
);

OAI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_3014),
.A2(n_1192),
.B1(n_1193),
.B2(n_1190),
.Y(n_3085)
);

OAI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_2992),
.A2(n_1203),
.B(n_1201),
.Y(n_3086)
);

OAI21xp33_ASAP7_75t_SL g3087 ( 
.A1(n_2998),
.A2(n_40),
.B(n_41),
.Y(n_3087)
);

OAI22xp33_ASAP7_75t_L g3088 ( 
.A1(n_3053),
.A2(n_1206),
.B1(n_1208),
.B2(n_1204),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2996),
.B(n_1211),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2997),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2994),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_3070),
.Y(n_3092)
);

XNOR2x1_ASAP7_75t_L g3093 ( 
.A(n_3041),
.B(n_1212),
.Y(n_3093)
);

OR2x2_ASAP7_75t_L g3094 ( 
.A(n_3071),
.B(n_3077),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_L g3095 ( 
.A(n_3081),
.B(n_1217),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_3005),
.B(n_1218),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_3072),
.A2(n_1219),
.B(n_40),
.Y(n_3097)
);

INVxp67_ASAP7_75t_L g3098 ( 
.A(n_3038),
.Y(n_3098)
);

OAI21xp33_ASAP7_75t_L g3099 ( 
.A1(n_3062),
.A2(n_42),
.B(n_43),
.Y(n_3099)
);

NAND3xp33_ASAP7_75t_L g3100 ( 
.A(n_3043),
.B(n_44),
.C(n_47),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_3037),
.Y(n_3101)
);

XNOR2x1_ASAP7_75t_L g3102 ( 
.A(n_2999),
.B(n_48),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3040),
.Y(n_3103)
);

INVx1_ASAP7_75t_SL g3104 ( 
.A(n_3024),
.Y(n_3104)
);

AOI31xp33_ASAP7_75t_L g3105 ( 
.A1(n_3079),
.A2(n_771),
.A3(n_772),
.B(n_770),
.Y(n_3105)
);

OAI221xp5_ASAP7_75t_SL g3106 ( 
.A1(n_2993),
.A2(n_50),
.B1(n_44),
.B2(n_48),
.C(n_51),
.Y(n_3106)
);

OAI31xp33_ASAP7_75t_L g3107 ( 
.A1(n_2993),
.A2(n_53),
.A3(n_51),
.B(n_52),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_3064),
.A2(n_2691),
.B1(n_1451),
.B2(n_54),
.Y(n_3108)
);

INVx1_ASAP7_75t_SL g3109 ( 
.A(n_3050),
.Y(n_3109)
);

XOR2x2_ASAP7_75t_L g3110 ( 
.A(n_3051),
.B(n_3052),
.Y(n_3110)
);

AOI22xp5_ASAP7_75t_L g3111 ( 
.A1(n_3082),
.A2(n_2691),
.B1(n_1451),
.B2(n_55),
.Y(n_3111)
);

OAI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_3026),
.A2(n_52),
.B(n_53),
.Y(n_3112)
);

OAI21xp5_ASAP7_75t_SL g3113 ( 
.A1(n_3082),
.A2(n_55),
.B(n_56),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_3084),
.A2(n_3013),
.B1(n_3039),
.B2(n_3018),
.Y(n_3114)
);

XNOR2xp5_ASAP7_75t_L g3115 ( 
.A(n_3001),
.B(n_58),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3011),
.Y(n_3116)
);

NAND3xp33_ASAP7_75t_L g3117 ( 
.A(n_3084),
.B(n_58),
.C(n_59),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_3008),
.A2(n_59),
.B(n_60),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_3068),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_3054),
.Y(n_3120)
);

AOI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_3008),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_3121)
);

OAI22xp33_ASAP7_75t_L g3122 ( 
.A1(n_3065),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_3122)
);

OAI221xp5_ASAP7_75t_L g3123 ( 
.A1(n_3066),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_3012),
.A2(n_65),
.B(n_66),
.Y(n_3124)
);

OAI21xp33_ASAP7_75t_L g3125 ( 
.A1(n_3075),
.A2(n_67),
.B(n_68),
.Y(n_3125)
);

AOI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_3061),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_3055),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_3005),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_3080),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_3022),
.Y(n_3130)
);

OAI22xp33_ASAP7_75t_L g3131 ( 
.A1(n_3028),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_3131)
);

OAI21xp5_ASAP7_75t_L g3132 ( 
.A1(n_3025),
.A2(n_75),
.B(n_76),
.Y(n_3132)
);

OAI22xp33_ASAP7_75t_L g3133 ( 
.A1(n_3027),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_3133)
);

OAI21xp33_ASAP7_75t_L g3134 ( 
.A1(n_3042),
.A2(n_77),
.B(n_78),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3023),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_3019),
.B(n_80),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3034),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3047),
.Y(n_3138)
);

NAND3xp33_ASAP7_75t_L g3139 ( 
.A(n_3057),
.B(n_81),
.C(n_82),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3004),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3017),
.Y(n_3141)
);

AOI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_3063),
.A2(n_84),
.B1(n_81),
.B2(n_82),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3015),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3002),
.Y(n_3144)
);

NAND3xp33_ASAP7_75t_L g3145 ( 
.A(n_3049),
.B(n_84),
.C(n_85),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3010),
.Y(n_3146)
);

OAI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_3021),
.A2(n_3036),
.B1(n_3029),
.B2(n_3078),
.Y(n_3147)
);

OAI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_3044),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_3148)
);

XOR2x2_ASAP7_75t_L g3149 ( 
.A(n_3020),
.B(n_87),
.Y(n_3149)
);

OAI21xp33_ASAP7_75t_L g3150 ( 
.A1(n_3032),
.A2(n_86),
.B(n_88),
.Y(n_3150)
);

AOI21xp33_ASAP7_75t_L g3151 ( 
.A1(n_3069),
.A2(n_88),
.B(n_89),
.Y(n_3151)
);

INVxp67_ASAP7_75t_L g3152 ( 
.A(n_3003),
.Y(n_3152)
);

XNOR2x2_ASAP7_75t_L g3153 ( 
.A(n_3006),
.B(n_89),
.Y(n_3153)
);

OAI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_3000),
.A2(n_90),
.B(n_91),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_3030),
.Y(n_3155)
);

NAND3xp33_ASAP7_75t_L g3156 ( 
.A(n_3058),
.B(n_90),
.C(n_91),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_3009),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3157)
);

OAI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_3007),
.A2(n_92),
.B(n_94),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_3067),
.B(n_3073),
.Y(n_3159)
);

AOI21xp33_ASAP7_75t_SL g3160 ( 
.A1(n_3074),
.A2(n_96),
.B(n_97),
.Y(n_3160)
);

AOI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_3076),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_3083),
.A2(n_98),
.B(n_100),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_L g3163 ( 
.A(n_3056),
.B(n_3048),
.Y(n_3163)
);

O2A1O1Ixp5_ASAP7_75t_L g3164 ( 
.A1(n_3016),
.A2(n_113),
.B(n_122),
.C(n_101),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_3031),
.Y(n_3165)
);

INVx1_ASAP7_75t_SL g3166 ( 
.A(n_3033),
.Y(n_3166)
);

HB1xp67_ASAP7_75t_L g3167 ( 
.A(n_3060),
.Y(n_3167)
);

OAI22xp5_ASAP7_75t_L g3168 ( 
.A1(n_3035),
.A2(n_107),
.B1(n_101),
.B2(n_104),
.Y(n_3168)
);

NAND3xp33_ASAP7_75t_L g3169 ( 
.A(n_3045),
.B(n_104),
.C(n_107),
.Y(n_3169)
);

XOR2x2_ASAP7_75t_L g3170 ( 
.A(n_3046),
.B(n_109),
.Y(n_3170)
);

AOI211xp5_ASAP7_75t_L g3171 ( 
.A1(n_3059),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2995),
.Y(n_3172)
);

AOI21xp5_ASAP7_75t_L g3173 ( 
.A1(n_3014),
.A2(n_108),
.B(n_110),
.Y(n_3173)
);

AOI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_3014),
.A2(n_114),
.B1(n_111),
.B2(n_112),
.Y(n_3174)
);

O2A1O1Ixp33_ASAP7_75t_SL g3175 ( 
.A1(n_3052),
.A2(n_114),
.B(n_111),
.C(n_112),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_3014),
.A2(n_118),
.B1(n_115),
.B2(n_116),
.Y(n_3176)
);

NOR3xp33_ASAP7_75t_L g3177 ( 
.A(n_3014),
.B(n_116),
.C(n_119),
.Y(n_3177)
);

AND2x4_ASAP7_75t_SL g3178 ( 
.A(n_2997),
.B(n_119),
.Y(n_3178)
);

AND2x4_ASAP7_75t_L g3179 ( 
.A(n_3071),
.B(n_120),
.Y(n_3179)
);

INVxp67_ASAP7_75t_L g3180 ( 
.A(n_2997),
.Y(n_3180)
);

OAI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_3014),
.A2(n_120),
.B(n_121),
.Y(n_3181)
);

OAI21xp33_ASAP7_75t_L g3182 ( 
.A1(n_3014),
.A2(n_121),
.B(n_122),
.Y(n_3182)
);

OAI21xp33_ASAP7_75t_L g3183 ( 
.A1(n_3014),
.A2(n_125),
.B(n_126),
.Y(n_3183)
);

OR2x2_ASAP7_75t_L g3184 ( 
.A(n_2997),
.B(n_126),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_3014),
.A2(n_127),
.B(n_128),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_3081),
.B(n_127),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_3014),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_SL g3188 ( 
.A(n_3081),
.B(n_129),
.Y(n_3188)
);

NAND4xp25_ASAP7_75t_SL g3189 ( 
.A(n_2992),
.B(n_132),
.C(n_130),
.D(n_131),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2999),
.Y(n_3190)
);

OAI21xp33_ASAP7_75t_L g3191 ( 
.A1(n_3014),
.A2(n_133),
.B(n_135),
.Y(n_3191)
);

OAI22xp5_ASAP7_75t_L g3192 ( 
.A1(n_3014),
.A2(n_139),
.B1(n_135),
.B2(n_137),
.Y(n_3192)
);

AOI22xp33_ASAP7_75t_SL g3193 ( 
.A1(n_3014),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_3193)
);

AOI22xp5_ASAP7_75t_L g3194 ( 
.A1(n_3014),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2999),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2997),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_3081),
.B(n_143),
.Y(n_3197)
);

OAI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_3014),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_3198)
);

CKINVDCx5p33_ASAP7_75t_R g3199 ( 
.A(n_3081),
.Y(n_3199)
);

AOI21xp33_ASAP7_75t_L g3200 ( 
.A1(n_3014),
.A2(n_144),
.B(n_146),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2997),
.Y(n_3201)
);

OAI21xp33_ASAP7_75t_L g3202 ( 
.A1(n_3014),
.A2(n_146),
.B(n_147),
.Y(n_3202)
);

NOR3xp33_ASAP7_75t_L g3203 ( 
.A(n_3014),
.B(n_148),
.C(n_149),
.Y(n_3203)
);

AOI22xp5_ASAP7_75t_L g3204 ( 
.A1(n_3014),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_3204)
);

OAI22xp33_ASAP7_75t_SL g3205 ( 
.A1(n_3014),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_3205)
);

AOI21xp33_ASAP7_75t_SL g3206 ( 
.A1(n_3081),
.A2(n_153),
.B(n_154),
.Y(n_3206)
);

NOR3xp33_ASAP7_75t_L g3207 ( 
.A(n_3014),
.B(n_153),
.C(n_154),
.Y(n_3207)
);

OAI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_3014),
.A2(n_155),
.B(n_156),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2997),
.Y(n_3209)
);

OAI21xp5_ASAP7_75t_SL g3210 ( 
.A1(n_3014),
.A2(n_156),
.B(n_157),
.Y(n_3210)
);

OAI211xp5_ASAP7_75t_L g3211 ( 
.A1(n_2992),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_3211)
);

OAI22xp33_ASAP7_75t_L g3212 ( 
.A1(n_3014),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_3212)
);

BUFx3_ASAP7_75t_L g3213 ( 
.A(n_2996),
.Y(n_3213)
);

AOI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_3014),
.A2(n_164),
.B1(n_161),
.B2(n_163),
.Y(n_3214)
);

OAI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_3014),
.A2(n_164),
.B(n_165),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2997),
.Y(n_3216)
);

AOI22xp5_ASAP7_75t_L g3217 ( 
.A1(n_3014),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_3217)
);

OAI22xp33_ASAP7_75t_L g3218 ( 
.A1(n_3014),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2999),
.Y(n_3219)
);

OAI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_3014),
.A2(n_170),
.B(n_171),
.Y(n_3220)
);

OAI21xp33_ASAP7_75t_L g3221 ( 
.A1(n_3014),
.A2(n_170),
.B(n_172),
.Y(n_3221)
);

INVxp67_ASAP7_75t_SL g3222 ( 
.A(n_3014),
.Y(n_3222)
);

AOI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_3014),
.A2(n_173),
.B(n_174),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2997),
.Y(n_3224)
);

NAND3xp33_ASAP7_75t_L g3225 ( 
.A(n_3014),
.B(n_173),
.C(n_174),
.Y(n_3225)
);

AOI22xp5_ASAP7_75t_L g3226 ( 
.A1(n_3014),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2997),
.Y(n_3227)
);

OAI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3014),
.A2(n_179),
.B1(n_175),
.B2(n_178),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_SL g3229 ( 
.A1(n_3014),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_3229)
);

AOI21xp33_ASAP7_75t_SL g3230 ( 
.A1(n_3081),
.A2(n_181),
.B(n_182),
.Y(n_3230)
);

AOI22xp5_ASAP7_75t_L g3231 ( 
.A1(n_3014),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_3231)
);

AOI211xp5_ASAP7_75t_SL g3232 ( 
.A1(n_3014),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_3232)
);

O2A1O1Ixp33_ASAP7_75t_L g3233 ( 
.A1(n_3014),
.A2(n_189),
.B(n_185),
.C(n_188),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_3014),
.A2(n_190),
.B(n_191),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2997),
.Y(n_3235)
);

INVx1_ASAP7_75t_SL g3236 ( 
.A(n_2996),
.Y(n_3236)
);

AOI21xp5_ASAP7_75t_L g3237 ( 
.A1(n_3014),
.A2(n_190),
.B(n_191),
.Y(n_3237)
);

OAI211xp5_ASAP7_75t_SL g3238 ( 
.A1(n_2992),
.A2(n_194),
.B(n_192),
.C(n_193),
.Y(n_3238)
);

INVxp67_ASAP7_75t_L g3239 ( 
.A(n_2997),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2997),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3199),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3102),
.Y(n_3242)
);

NOR4xp25_ASAP7_75t_L g3243 ( 
.A(n_3222),
.B(n_195),
.C(n_192),
.D(n_193),
.Y(n_3243)
);

AOI22xp33_ASAP7_75t_L g3244 ( 
.A1(n_3109),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_3244)
);

AOI22xp33_ASAP7_75t_SL g3245 ( 
.A1(n_3153),
.A2(n_3104),
.B1(n_3087),
.B2(n_3085),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_3213),
.B(n_3236),
.Y(n_3246)
);

AOI222xp33_ASAP7_75t_L g3247 ( 
.A1(n_3087),
.A2(n_198),
.B1(n_201),
.B2(n_196),
.C1(n_197),
.C2(n_199),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3186),
.Y(n_3248)
);

OAI22xp5_ASAP7_75t_L g3249 ( 
.A1(n_3094),
.A2(n_202),
.B1(n_199),
.B2(n_201),
.Y(n_3249)
);

AOI221xp5_ASAP7_75t_L g3250 ( 
.A1(n_3098),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.C(n_206),
.Y(n_3250)
);

AOI22xp5_ASAP7_75t_SL g3251 ( 
.A1(n_3205),
.A2(n_206),
.B1(n_203),
.B2(n_204),
.Y(n_3251)
);

OAI332xp33_ASAP7_75t_L g3252 ( 
.A1(n_3166),
.A2(n_214),
.A3(n_213),
.B1(n_209),
.B2(n_215),
.B3(n_207),
.C1(n_208),
.C2(n_210),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3232),
.B(n_207),
.Y(n_3253)
);

OAI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3173),
.A2(n_210),
.B(n_216),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3197),
.Y(n_3255)
);

INVxp67_ASAP7_75t_L g3256 ( 
.A(n_3095),
.Y(n_3256)
);

AOI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_3177),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3184),
.Y(n_3258)
);

NOR2x1_ASAP7_75t_SL g3259 ( 
.A(n_3188),
.B(n_217),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_3110),
.Y(n_3260)
);

AOI221xp5_ASAP7_75t_SL g3261 ( 
.A1(n_3180),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.C(n_222),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3179),
.Y(n_3262)
);

NAND3xp33_ASAP7_75t_L g3263 ( 
.A(n_3203),
.B(n_222),
.C(n_223),
.Y(n_3263)
);

AOI22xp5_ASAP7_75t_L g3264 ( 
.A1(n_3163),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_3264)
);

OAI21xp5_ASAP7_75t_SL g3265 ( 
.A1(n_3239),
.A2(n_226),
.B(n_227),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3179),
.B(n_226),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3206),
.B(n_227),
.Y(n_3267)
);

OAI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_3185),
.A2(n_228),
.B(n_229),
.Y(n_3268)
);

OAI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_3135),
.A2(n_231),
.B1(n_228),
.B2(n_230),
.Y(n_3269)
);

AOI321xp33_ASAP7_75t_L g3270 ( 
.A1(n_3114),
.A2(n_233),
.A3(n_235),
.B1(n_236),
.B2(n_231),
.C(n_234),
.Y(n_3270)
);

NAND3xp33_ASAP7_75t_L g3271 ( 
.A(n_3207),
.B(n_230),
.C(n_233),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_3230),
.B(n_235),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3175),
.A2(n_236),
.B(n_237),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3091),
.B(n_238),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3178),
.B(n_239),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3128),
.B(n_3105),
.Y(n_3276)
);

NAND2xp33_ASAP7_75t_L g3277 ( 
.A(n_3092),
.B(n_240),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_3089),
.B(n_3118),
.Y(n_3278)
);

OAI22xp5_ASAP7_75t_L g3279 ( 
.A1(n_3190),
.A2(n_244),
.B1(n_241),
.B2(n_242),
.Y(n_3279)
);

AND3x1_ASAP7_75t_L g3280 ( 
.A(n_3195),
.B(n_242),
.C(n_245),
.Y(n_3280)
);

AOI221xp5_ASAP7_75t_L g3281 ( 
.A1(n_3223),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.C(n_248),
.Y(n_3281)
);

A2O1A1Ixp33_ASAP7_75t_L g3282 ( 
.A1(n_3234),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_3237),
.A2(n_251),
.B(n_252),
.Y(n_3283)
);

AOI22xp5_ASAP7_75t_L g3284 ( 
.A1(n_3159),
.A2(n_255),
.B1(n_252),
.B2(n_253),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_3219),
.Y(n_3285)
);

OAI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_3174),
.A2(n_259),
.B1(n_256),
.B2(n_257),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3167),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3143),
.B(n_259),
.Y(n_3288)
);

INVxp67_ASAP7_75t_L g3289 ( 
.A(n_3096),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_3120),
.Y(n_3290)
);

AND2x4_ASAP7_75t_SL g3291 ( 
.A(n_3127),
.B(n_260),
.Y(n_3291)
);

AOI22xp5_ASAP7_75t_L g3292 ( 
.A1(n_3116),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_3292)
);

OR2x2_ASAP7_75t_L g3293 ( 
.A(n_3101),
.B(n_262),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_3090),
.B(n_3196),
.Y(n_3294)
);

AOI221xp5_ASAP7_75t_L g3295 ( 
.A1(n_3200),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_267),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_3201),
.B(n_263),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3233),
.A2(n_265),
.B(n_267),
.Y(n_3297)
);

INVx1_ASAP7_75t_SL g3298 ( 
.A(n_3170),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3193),
.B(n_269),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3155),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3138),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3137),
.Y(n_3302)
);

OAI22xp5_ASAP7_75t_L g3303 ( 
.A1(n_3229),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_3130),
.A2(n_275),
.B1(n_270),
.B2(n_273),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_R g3305 ( 
.A1(n_3147),
.A2(n_273),
.B(n_275),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3093),
.B(n_276),
.Y(n_3306)
);

INVxp67_ASAP7_75t_L g3307 ( 
.A(n_3136),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3209),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3149),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3113),
.B(n_276),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3216),
.Y(n_3311)
);

AOI21xp33_ASAP7_75t_L g3312 ( 
.A1(n_3088),
.A2(n_277),
.B(n_278),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3224),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3227),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3140),
.Y(n_3315)
);

AOI21xp33_ASAP7_75t_SL g3316 ( 
.A1(n_3172),
.A2(n_277),
.B(n_278),
.Y(n_3316)
);

OR2x2_ASAP7_75t_L g3317 ( 
.A(n_3103),
.B(n_279),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_3235),
.B(n_279),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_SL g3319 ( 
.A1(n_3225),
.A2(n_3181),
.B1(n_3215),
.B2(n_3208),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3240),
.Y(n_3320)
);

OAI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3176),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3321)
);

AOI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3141),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3210),
.B(n_285),
.Y(n_3323)
);

AND3x1_ASAP7_75t_L g3324 ( 
.A(n_3182),
.B(n_3191),
.C(n_3183),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_3212),
.B(n_285),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3164),
.Y(n_3326)
);

OR2x2_ASAP7_75t_L g3327 ( 
.A(n_3119),
.B(n_286),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3129),
.Y(n_3328)
);

AOI222xp33_ASAP7_75t_L g3329 ( 
.A1(n_3220),
.A2(n_288),
.B1(n_290),
.B2(n_286),
.C1(n_287),
.C2(n_289),
.Y(n_3329)
);

OAI31xp33_ASAP7_75t_L g3330 ( 
.A1(n_3192),
.A2(n_291),
.A3(n_289),
.B(n_290),
.Y(n_3330)
);

NAND2xp33_ASAP7_75t_L g3331 ( 
.A(n_3125),
.B(n_3165),
.Y(n_3331)
);

AOI32xp33_ASAP7_75t_L g3332 ( 
.A1(n_3218),
.A2(n_294),
.A3(n_292),
.B1(n_293),
.B2(n_295),
.Y(n_3332)
);

OAI21xp33_ASAP7_75t_L g3333 ( 
.A1(n_3152),
.A2(n_292),
.B(n_293),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_L g3334 ( 
.A1(n_3202),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_3334)
);

NAND3xp33_ASAP7_75t_L g3335 ( 
.A(n_3187),
.B(n_296),
.C(n_297),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3121),
.B(n_298),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3117),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3198),
.Y(n_3338)
);

AOI221xp5_ASAP7_75t_L g3339 ( 
.A1(n_3221),
.A2(n_304),
.B1(n_300),
.B2(n_303),
.C(n_305),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_3132),
.B(n_300),
.Y(n_3340)
);

OAI21xp33_ASAP7_75t_L g3341 ( 
.A1(n_3194),
.A2(n_303),
.B(n_304),
.Y(n_3341)
);

AOI22xp33_ASAP7_75t_L g3342 ( 
.A1(n_3124),
.A2(n_3238),
.B1(n_3112),
.B2(n_3162),
.Y(n_3342)
);

OR2x2_ASAP7_75t_L g3343 ( 
.A(n_3144),
.B(n_777),
.Y(n_3343)
);

INVxp67_ASAP7_75t_SL g3344 ( 
.A(n_3171),
.Y(n_3344)
);

AOI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_3204),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_3345)
);

NAND2x1_ASAP7_75t_L g3346 ( 
.A(n_3146),
.B(n_307),
.Y(n_3346)
);

OAI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_3214),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3133),
.B(n_309),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_3217),
.A2(n_3226),
.B1(n_3231),
.B2(n_3228),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3115),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3169),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3154),
.B(n_311),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3168),
.Y(n_3353)
);

AOI21xp5_ASAP7_75t_L g3354 ( 
.A1(n_3097),
.A2(n_311),
.B(n_312),
.Y(n_3354)
);

INVxp67_ASAP7_75t_L g3355 ( 
.A(n_3189),
.Y(n_3355)
);

AOI21xp33_ASAP7_75t_L g3356 ( 
.A1(n_3150),
.A2(n_312),
.B(n_313),
.Y(n_3356)
);

INVx1_ASAP7_75t_SL g3357 ( 
.A(n_3142),
.Y(n_3357)
);

OAI21xp33_ASAP7_75t_L g3358 ( 
.A1(n_3099),
.A2(n_313),
.B(n_314),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3145),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3157),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3161),
.Y(n_3361)
);

AOI211xp5_ASAP7_75t_L g3362 ( 
.A1(n_3106),
.A2(n_317),
.B(n_314),
.C(n_316),
.Y(n_3362)
);

INVxp67_ASAP7_75t_L g3363 ( 
.A(n_3100),
.Y(n_3363)
);

AOI22xp33_ASAP7_75t_L g3364 ( 
.A1(n_3108),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_3158),
.A2(n_322),
.B1(n_319),
.B2(n_321),
.Y(n_3365)
);

OAI221xp5_ASAP7_75t_L g3366 ( 
.A1(n_3111),
.A2(n_323),
.B1(n_319),
.B2(n_322),
.C(n_324),
.Y(n_3366)
);

AOI211xp5_ASAP7_75t_L g3367 ( 
.A1(n_3151),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_3367)
);

INVxp67_ASAP7_75t_L g3368 ( 
.A(n_3280),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3266),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3243),
.B(n_3122),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3288),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3253),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3251),
.B(n_3131),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3242),
.B(n_3107),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3247),
.B(n_3134),
.Y(n_3375)
);

AOI31xp33_ASAP7_75t_L g3376 ( 
.A1(n_3241),
.A2(n_3246),
.A3(n_3285),
.B(n_3287),
.Y(n_3376)
);

OAI21xp33_ASAP7_75t_L g3377 ( 
.A1(n_3290),
.A2(n_3126),
.B(n_3139),
.Y(n_3377)
);

NOR2xp67_ASAP7_75t_L g3378 ( 
.A(n_3326),
.B(n_3156),
.Y(n_3378)
);

AOI221xp5_ASAP7_75t_L g3379 ( 
.A1(n_3324),
.A2(n_3160),
.B1(n_3148),
.B2(n_3123),
.C(n_3211),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3298),
.B(n_3086),
.Y(n_3380)
);

AOI22xp5_ASAP7_75t_L g3381 ( 
.A1(n_3248),
.A2(n_328),
.B1(n_325),
.B2(n_327),
.Y(n_3381)
);

NAND3xp33_ASAP7_75t_L g3382 ( 
.A(n_3245),
.B(n_328),
.C(n_329),
.Y(n_3382)
);

AOI221xp5_ASAP7_75t_SL g3383 ( 
.A1(n_3331),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_3383)
);

INVx3_ASAP7_75t_L g3384 ( 
.A(n_3346),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_3259),
.Y(n_3385)
);

HB1xp67_ASAP7_75t_L g3386 ( 
.A(n_3276),
.Y(n_3386)
);

AOI322xp5_ASAP7_75t_L g3387 ( 
.A1(n_3342),
.A2(n_337),
.A3(n_336),
.B1(n_334),
.B2(n_332),
.C1(n_333),
.C2(n_335),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3262),
.Y(n_3388)
);

AOI21xp33_ASAP7_75t_L g3389 ( 
.A1(n_3307),
.A2(n_334),
.B(n_335),
.Y(n_3389)
);

INVxp67_ASAP7_75t_L g3390 ( 
.A(n_3275),
.Y(n_3390)
);

AND2x4_ASAP7_75t_L g3391 ( 
.A(n_3315),
.B(n_336),
.Y(n_3391)
);

AOI21xp33_ASAP7_75t_SL g3392 ( 
.A1(n_3274),
.A2(n_338),
.B(n_339),
.Y(n_3392)
);

AOI22xp5_ASAP7_75t_L g3393 ( 
.A1(n_3255),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_3393)
);

OAI21xp33_ASAP7_75t_L g3394 ( 
.A1(n_3294),
.A2(n_340),
.B(n_341),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3327),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_3265),
.B(n_341),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3273),
.B(n_342),
.Y(n_3397)
);

OR2x2_ASAP7_75t_L g3398 ( 
.A(n_3293),
.B(n_342),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3261),
.B(n_343),
.Y(n_3399)
);

AOI32xp33_ASAP7_75t_L g3400 ( 
.A1(n_3351),
.A2(n_347),
.A3(n_345),
.B1(n_346),
.B2(n_349),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3291),
.B(n_3258),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3343),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3296),
.B(n_3318),
.Y(n_3403)
);

OAI21xp5_ASAP7_75t_SL g3404 ( 
.A1(n_3301),
.A2(n_345),
.B(n_346),
.Y(n_3404)
);

INVxp67_ASAP7_75t_SL g3405 ( 
.A(n_3277),
.Y(n_3405)
);

AOI21xp33_ASAP7_75t_L g3406 ( 
.A1(n_3278),
.A2(n_347),
.B(n_349),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3317),
.Y(n_3407)
);

AOI221xp5_ASAP7_75t_L g3408 ( 
.A1(n_3316),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.C(n_353),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_SL g3409 ( 
.A(n_3270),
.B(n_351),
.Y(n_3409)
);

NAND3xp33_ASAP7_75t_L g3410 ( 
.A(n_3362),
.B(n_354),
.C(n_355),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3306),
.Y(n_3411)
);

INVxp67_ASAP7_75t_L g3412 ( 
.A(n_3267),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3272),
.Y(n_3413)
);

AO22x1_ASAP7_75t_L g3414 ( 
.A1(n_3344),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_3414)
);

AND2x2_ASAP7_75t_L g3415 ( 
.A(n_3302),
.B(n_356),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3252),
.B(n_357),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3310),
.Y(n_3417)
);

OAI221xp5_ASAP7_75t_SL g3418 ( 
.A1(n_3260),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.C(n_362),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3308),
.B(n_360),
.Y(n_3419)
);

NOR2xp33_ASAP7_75t_L g3420 ( 
.A(n_3355),
.B(n_362),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3323),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3299),
.Y(n_3422)
);

OAI22xp33_ASAP7_75t_L g3423 ( 
.A1(n_3349),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3300),
.Y(n_3424)
);

AOI31xp33_ASAP7_75t_L g3425 ( 
.A1(n_3311),
.A2(n_366),
.A3(n_363),
.B(n_364),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_3309),
.A2(n_371),
.B1(n_367),
.B2(n_369),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_3313),
.B(n_367),
.Y(n_3427)
);

O2A1O1Ixp33_ASAP7_75t_L g3428 ( 
.A1(n_3282),
.A2(n_374),
.B(n_369),
.C(n_372),
.Y(n_3428)
);

INVxp67_ASAP7_75t_L g3429 ( 
.A(n_3352),
.Y(n_3429)
);

AOI32xp33_ASAP7_75t_L g3430 ( 
.A1(n_3337),
.A2(n_377),
.A3(n_375),
.B1(n_376),
.B2(n_378),
.Y(n_3430)
);

O2A1O1Ixp33_ASAP7_75t_L g3431 ( 
.A1(n_3363),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_3431)
);

NOR3xp33_ASAP7_75t_SL g3432 ( 
.A(n_3314),
.B(n_3320),
.C(n_3328),
.Y(n_3432)
);

AOI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3256),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_SL g3434 ( 
.A1(n_3303),
.A2(n_382),
.B(n_383),
.Y(n_3434)
);

OAI33xp33_ASAP7_75t_L g3435 ( 
.A1(n_3353),
.A2(n_3338),
.A3(n_3289),
.B1(n_3360),
.B2(n_3361),
.B3(n_3325),
.Y(n_3435)
);

NOR2xp33_ASAP7_75t_L g3436 ( 
.A(n_3333),
.B(n_383),
.Y(n_3436)
);

OAI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3244),
.A2(n_389),
.B1(n_385),
.B2(n_388),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3257),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3319),
.B(n_385),
.Y(n_3439)
);

OAI22xp5_ASAP7_75t_L g3440 ( 
.A1(n_3334),
.A2(n_393),
.B1(n_388),
.B2(n_391),
.Y(n_3440)
);

INVxp67_ASAP7_75t_L g3441 ( 
.A(n_3340),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3257),
.Y(n_3442)
);

OAI21xp33_ASAP7_75t_L g3443 ( 
.A1(n_3349),
.A2(n_391),
.B(n_393),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3348),
.Y(n_3444)
);

OAI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_3305),
.A2(n_397),
.B1(n_394),
.B2(n_395),
.Y(n_3445)
);

AOI221xp5_ASAP7_75t_L g3446 ( 
.A1(n_3354),
.A2(n_400),
.B1(n_395),
.B2(n_398),
.C(n_401),
.Y(n_3446)
);

AOI211xp5_ASAP7_75t_L g3447 ( 
.A1(n_3279),
.A2(n_403),
.B(n_401),
.C(n_402),
.Y(n_3447)
);

OAI211xp5_ASAP7_75t_SL g3448 ( 
.A1(n_3329),
.A2(n_405),
.B(n_403),
.C(n_404),
.Y(n_3448)
);

OAI31xp33_ASAP7_75t_L g3449 ( 
.A1(n_3357),
.A2(n_407),
.A3(n_405),
.B(n_406),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3336),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3283),
.B(n_408),
.Y(n_3451)
);

AO21x1_ASAP7_75t_L g3452 ( 
.A1(n_3249),
.A2(n_409),
.B(n_410),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3359),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3263),
.Y(n_3454)
);

AOI221xp5_ASAP7_75t_L g3455 ( 
.A1(n_3254),
.A2(n_3268),
.B1(n_3297),
.B2(n_3341),
.C(n_3366),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3271),
.Y(n_3456)
);

AOI21xp33_ASAP7_75t_L g3457 ( 
.A1(n_3350),
.A2(n_412),
.B(n_413),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3284),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3332),
.B(n_412),
.Y(n_3459)
);

INVx1_ASAP7_75t_SL g3460 ( 
.A(n_3345),
.Y(n_3460)
);

XNOR2xp5_ASAP7_75t_L g3461 ( 
.A(n_3367),
.B(n_414),
.Y(n_3461)
);

OAI221xp5_ASAP7_75t_SL g3462 ( 
.A1(n_3358),
.A2(n_777),
.B1(n_417),
.B2(n_415),
.C(n_416),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3269),
.Y(n_3463)
);

OAI221xp5_ASAP7_75t_L g3464 ( 
.A1(n_3345),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.C(n_420),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3281),
.B(n_419),
.Y(n_3465)
);

AOI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_3347),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3330),
.B(n_421),
.Y(n_3467)
);

OAI221xp5_ASAP7_75t_L g3468 ( 
.A1(n_3364),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.C(n_428),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3292),
.B(n_425),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3365),
.B(n_426),
.Y(n_3470)
);

INVxp67_ASAP7_75t_L g3471 ( 
.A(n_3335),
.Y(n_3471)
);

OR2x2_ASAP7_75t_L g3472 ( 
.A(n_3304),
.B(n_427),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3264),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3286),
.B(n_3321),
.Y(n_3474)
);

OAI31xp33_ASAP7_75t_L g3475 ( 
.A1(n_3356),
.A2(n_431),
.A3(n_429),
.B(n_430),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_3312),
.A2(n_429),
.B(n_430),
.Y(n_3476)
);

HB1xp67_ASAP7_75t_L g3477 ( 
.A(n_3339),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3322),
.Y(n_3478)
);

OAI22xp33_ASAP7_75t_L g3479 ( 
.A1(n_3295),
.A2(n_776),
.B1(n_433),
.B2(n_431),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3250),
.Y(n_3480)
);

OR2x2_ASAP7_75t_L g3481 ( 
.A(n_3326),
.B(n_432),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3243),
.B(n_433),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3266),
.Y(n_3483)
);

AOI222xp33_ASAP7_75t_L g3484 ( 
.A1(n_3326),
.A2(n_436),
.B1(n_438),
.B2(n_434),
.C1(n_435),
.C2(n_437),
.Y(n_3484)
);

AOI21xp33_ASAP7_75t_L g3485 ( 
.A1(n_3326),
.A2(n_434),
.B(n_435),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3266),
.Y(n_3486)
);

AOI21xp33_ASAP7_75t_L g3487 ( 
.A1(n_3326),
.A2(n_437),
.B(n_438),
.Y(n_3487)
);

AOI22xp5_ASAP7_75t_L g3488 ( 
.A1(n_3298),
.A2(n_443),
.B1(n_439),
.B2(n_440),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3326),
.B(n_440),
.Y(n_3489)
);

AOI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3298),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_3490)
);

AOI21xp5_ASAP7_75t_L g3491 ( 
.A1(n_3277),
.A2(n_444),
.B(n_445),
.Y(n_3491)
);

OAI21xp33_ASAP7_75t_L g3492 ( 
.A1(n_3285),
.A2(n_446),
.B(n_447),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3248),
.A2(n_449),
.B1(n_446),
.B2(n_447),
.Y(n_3493)
);

NOR3xp33_ASAP7_75t_SL g3494 ( 
.A(n_3241),
.B(n_774),
.C(n_449),
.Y(n_3494)
);

INVxp67_ASAP7_75t_SL g3495 ( 
.A(n_3259),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3243),
.B(n_450),
.Y(n_3496)
);

OAI221xp5_ASAP7_75t_L g3497 ( 
.A1(n_3243),
.A2(n_453),
.B1(n_450),
.B2(n_451),
.C(n_454),
.Y(n_3497)
);

OAI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_3326),
.A2(n_455),
.B1(n_451),
.B2(n_454),
.Y(n_3498)
);

OR2x2_ASAP7_75t_L g3499 ( 
.A(n_3326),
.B(n_455),
.Y(n_3499)
);

AOI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3298),
.A2(n_459),
.B1(n_456),
.B2(n_458),
.Y(n_3500)
);

AOI21xp33_ASAP7_75t_L g3501 ( 
.A1(n_3326),
.A2(n_456),
.B(n_458),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3280),
.Y(n_3502)
);

OAI32xp33_ASAP7_75t_L g3503 ( 
.A1(n_3326),
.A2(n_773),
.A3(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_3503)
);

OAI22xp33_ASAP7_75t_SL g3504 ( 
.A1(n_3298),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3266),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3266),
.Y(n_3506)
);

OR2x2_ASAP7_75t_L g3507 ( 
.A(n_3326),
.B(n_463),
.Y(n_3507)
);

AOI32xp33_ASAP7_75t_L g3508 ( 
.A1(n_3326),
.A2(n_465),
.A3(n_463),
.B1(n_464),
.B2(n_467),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3246),
.B(n_465),
.Y(n_3509)
);

INVxp67_ASAP7_75t_SL g3510 ( 
.A(n_3259),
.Y(n_3510)
);

OAI221xp5_ASAP7_75t_L g3511 ( 
.A1(n_3243),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.C(n_471),
.Y(n_3511)
);

AOI222xp33_ASAP7_75t_L g3512 ( 
.A1(n_3326),
.A2(n_468),
.B1(n_470),
.B2(n_472),
.C1(n_474),
.C2(n_475),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3243),
.B(n_474),
.Y(n_3513)
);

AOI221xp5_ASAP7_75t_L g3514 ( 
.A1(n_3243),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.C(n_479),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3298),
.B(n_478),
.Y(n_3515)
);

OAI21xp5_ASAP7_75t_SL g3516 ( 
.A1(n_3326),
.A2(n_480),
.B(n_481),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3266),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3246),
.B(n_480),
.Y(n_3518)
);

AOI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3298),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_3519)
);

OAI321xp33_ASAP7_75t_L g3520 ( 
.A1(n_3241),
.A2(n_483),
.A3(n_485),
.B1(n_486),
.B2(n_487),
.C(n_489),
.Y(n_3520)
);

AOI222xp33_ASAP7_75t_L g3521 ( 
.A1(n_3326),
.A2(n_485),
.B1(n_489),
.B2(n_490),
.C1(n_491),
.C2(n_493),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3266),
.Y(n_3522)
);

OR2x2_ASAP7_75t_L g3523 ( 
.A(n_3326),
.B(n_494),
.Y(n_3523)
);

AOI21xp33_ASAP7_75t_L g3524 ( 
.A1(n_3326),
.A2(n_495),
.B(n_496),
.Y(n_3524)
);

NOR2xp67_ASAP7_75t_SL g3525 ( 
.A(n_3241),
.B(n_495),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3277),
.A2(n_497),
.B(n_499),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_SL g3527 ( 
.A(n_3384),
.B(n_499),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3414),
.B(n_3403),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3376),
.A2(n_500),
.B(n_501),
.Y(n_3529)
);

O2A1O1Ixp5_ASAP7_75t_L g3530 ( 
.A1(n_3384),
.A2(n_502),
.B(n_500),
.C(n_501),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3509),
.B(n_502),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3504),
.B(n_503),
.Y(n_3532)
);

AOI211xp5_ASAP7_75t_L g3533 ( 
.A1(n_3485),
.A2(n_3487),
.B(n_3524),
.C(n_3501),
.Y(n_3533)
);

NAND2x1_ASAP7_75t_L g3534 ( 
.A(n_3518),
.B(n_503),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3391),
.Y(n_3535)
);

NOR2xp67_ASAP7_75t_L g3536 ( 
.A(n_3386),
.B(n_504),
.Y(n_3536)
);

OAI221xp5_ASAP7_75t_L g3537 ( 
.A1(n_3495),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.C(n_507),
.Y(n_3537)
);

AOI211xp5_ASAP7_75t_L g3538 ( 
.A1(n_3516),
.A2(n_773),
.B(n_509),
.C(n_506),
.Y(n_3538)
);

NOR2xp33_ASAP7_75t_L g3539 ( 
.A(n_3435),
.B(n_508),
.Y(n_3539)
);

NOR3xp33_ASAP7_75t_L g3540 ( 
.A(n_3382),
.B(n_772),
.C(n_508),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3509),
.B(n_509),
.Y(n_3541)
);

AND2x4_ASAP7_75t_L g3542 ( 
.A(n_3510),
.B(n_510),
.Y(n_3542)
);

OAI21xp33_ASAP7_75t_SL g3543 ( 
.A1(n_3378),
.A2(n_510),
.B(n_511),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3425),
.B(n_511),
.Y(n_3544)
);

OAI21xp33_ASAP7_75t_L g3545 ( 
.A1(n_3405),
.A2(n_512),
.B(n_513),
.Y(n_3545)
);

NOR2xp33_ASAP7_75t_L g3546 ( 
.A(n_3385),
.B(n_513),
.Y(n_3546)
);

AOI21xp33_ASAP7_75t_L g3547 ( 
.A1(n_3368),
.A2(n_514),
.B(n_515),
.Y(n_3547)
);

HB1xp67_ASAP7_75t_L g3548 ( 
.A(n_3391),
.Y(n_3548)
);

AOI211xp5_ASAP7_75t_L g3549 ( 
.A1(n_3481),
.A2(n_771),
.B(n_517),
.C(n_515),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3398),
.Y(n_3550)
);

NAND3xp33_ASAP7_75t_L g3551 ( 
.A(n_3449),
.B(n_516),
.C(n_517),
.Y(n_3551)
);

INVxp67_ASAP7_75t_SL g3552 ( 
.A(n_3482),
.Y(n_3552)
);

NOR3xp33_ASAP7_75t_SL g3553 ( 
.A(n_3401),
.B(n_516),
.C(n_518),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3497),
.B(n_520),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3494),
.B(n_521),
.Y(n_3555)
);

AOI211x1_ASAP7_75t_L g3556 ( 
.A1(n_3377),
.A2(n_523),
.B(n_521),
.C(n_522),
.Y(n_3556)
);

AOI221xp5_ASAP7_75t_L g3557 ( 
.A1(n_3372),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.C(n_525),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3511),
.B(n_525),
.Y(n_3558)
);

NOR3xp33_ASAP7_75t_L g3559 ( 
.A(n_3515),
.B(n_526),
.C(n_527),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3383),
.B(n_527),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3525),
.B(n_528),
.Y(n_3561)
);

NOR2x1_ASAP7_75t_L g3562 ( 
.A(n_3489),
.B(n_529),
.Y(n_3562)
);

OAI22xp33_ASAP7_75t_L g3563 ( 
.A1(n_3496),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3513),
.Y(n_3564)
);

NOR3x1_ASAP7_75t_L g3565 ( 
.A(n_3404),
.B(n_530),
.C(n_531),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3415),
.B(n_532),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_SL g3567 ( 
.A(n_3514),
.B(n_532),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_3416),
.A2(n_770),
.B(n_534),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3461),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3409),
.A2(n_534),
.B(n_535),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3503),
.A2(n_3399),
.B(n_3397),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3371),
.B(n_536),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3419),
.B(n_537),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_3439),
.A2(n_767),
.B(n_537),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3427),
.Y(n_3575)
);

NAND3xp33_ASAP7_75t_L g3576 ( 
.A(n_3432),
.B(n_540),
.C(n_541),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3407),
.B(n_541),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3502),
.Y(n_3578)
);

NOR2xp33_ASAP7_75t_L g3579 ( 
.A(n_3418),
.B(n_542),
.Y(n_3579)
);

OAI21xp33_ASAP7_75t_L g3580 ( 
.A1(n_3453),
.A2(n_543),
.B(n_544),
.Y(n_3580)
);

CKINVDCx5p33_ASAP7_75t_R g3581 ( 
.A(n_3420),
.Y(n_3581)
);

INVx2_ASAP7_75t_SL g3582 ( 
.A(n_3499),
.Y(n_3582)
);

INVx1_ASAP7_75t_SL g3583 ( 
.A(n_3507),
.Y(n_3583)
);

OR2x2_ASAP7_75t_L g3584 ( 
.A(n_3523),
.B(n_767),
.Y(n_3584)
);

AOI211xp5_ASAP7_75t_L g3585 ( 
.A1(n_3498),
.A2(n_545),
.B(n_543),
.C(n_544),
.Y(n_3585)
);

NOR2xp33_ASAP7_75t_SL g3586 ( 
.A(n_3462),
.B(n_545),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_SL g3587 ( 
.A(n_3484),
.B(n_546),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3392),
.B(n_547),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_SL g3589 ( 
.A(n_3512),
.B(n_548),
.Y(n_3589)
);

NOR3xp33_ASAP7_75t_SL g3590 ( 
.A(n_3424),
.B(n_548),
.C(n_549),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_L g3591 ( 
.A(n_3491),
.B(n_550),
.Y(n_3591)
);

NOR3x1_ASAP7_75t_L g3592 ( 
.A(n_3410),
.B(n_551),
.C(n_552),
.Y(n_3592)
);

NOR3x1_ASAP7_75t_L g3593 ( 
.A(n_3370),
.B(n_3375),
.C(n_3454),
.Y(n_3593)
);

AOI221xp5_ASAP7_75t_SL g3594 ( 
.A1(n_3471),
.A2(n_551),
.B1(n_553),
.B2(n_554),
.C(n_555),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3451),
.Y(n_3595)
);

OAI21xp33_ASAP7_75t_L g3596 ( 
.A1(n_3458),
.A2(n_554),
.B(n_555),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3526),
.A2(n_766),
.B(n_556),
.Y(n_3597)
);

NOR3x1_ASAP7_75t_L g3598 ( 
.A(n_3456),
.B(n_556),
.C(n_557),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_SL g3599 ( 
.A(n_3521),
.B(n_559),
.Y(n_3599)
);

AOI221xp5_ASAP7_75t_L g3600 ( 
.A1(n_3417),
.A2(n_559),
.B1(n_560),
.B2(n_561),
.C(n_562),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3395),
.B(n_560),
.Y(n_3601)
);

NOR2xp33_ASAP7_75t_L g3602 ( 
.A(n_3448),
.B(n_562),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_3408),
.B(n_564),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3431),
.A2(n_564),
.B(n_565),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3452),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3402),
.B(n_565),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3388),
.Y(n_3607)
);

NAND3xp33_ASAP7_75t_L g3608 ( 
.A(n_3508),
.B(n_3475),
.C(n_3443),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3441),
.B(n_566),
.Y(n_3609)
);

NAND3xp33_ASAP7_75t_L g3610 ( 
.A(n_3429),
.B(n_566),
.C(n_567),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3380),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3396),
.B(n_3488),
.Y(n_3612)
);

NOR4xp75_ASAP7_75t_L g3613 ( 
.A(n_3374),
.B(n_570),
.C(n_568),
.D(n_569),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3434),
.A2(n_765),
.B(n_568),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3445),
.B(n_569),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3373),
.Y(n_3616)
);

NAND3xp33_ASAP7_75t_L g3617 ( 
.A(n_3430),
.B(n_572),
.C(n_573),
.Y(n_3617)
);

NOR3x1_ASAP7_75t_L g3618 ( 
.A(n_3459),
.B(n_572),
.C(n_573),
.Y(n_3618)
);

NOR2xp33_ASAP7_75t_L g3619 ( 
.A(n_3492),
.B(n_574),
.Y(n_3619)
);

NAND3xp33_ASAP7_75t_SL g3620 ( 
.A(n_3460),
.B(n_574),
.C(n_575),
.Y(n_3620)
);

OAI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3528),
.A2(n_3422),
.B1(n_3500),
.B2(n_3490),
.Y(n_3621)
);

OAI211xp5_ASAP7_75t_L g3622 ( 
.A1(n_3529),
.A2(n_3394),
.B(n_3400),
.C(n_3480),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3556),
.B(n_3387),
.Y(n_3623)
);

OAI21xp33_ASAP7_75t_L g3624 ( 
.A1(n_3586),
.A2(n_3463),
.B(n_3444),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3553),
.B(n_3379),
.Y(n_3625)
);

OAI32xp33_ASAP7_75t_L g3626 ( 
.A1(n_3539),
.A2(n_3607),
.A3(n_3605),
.B1(n_3543),
.B2(n_3616),
.Y(n_3626)
);

A2O1A1Ixp33_ASAP7_75t_L g3627 ( 
.A1(n_3568),
.A2(n_3428),
.B(n_3421),
.C(n_3390),
.Y(n_3627)
);

AOI311xp33_ASAP7_75t_L g3628 ( 
.A1(n_3564),
.A2(n_3413),
.A3(n_3450),
.B(n_3369),
.C(n_3517),
.Y(n_3628)
);

AOI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_3552),
.A2(n_3412),
.B1(n_3469),
.B2(n_3411),
.Y(n_3629)
);

OAI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3560),
.A2(n_3519),
.B1(n_3472),
.B2(n_3465),
.Y(n_3630)
);

AOI221xp5_ASAP7_75t_L g3631 ( 
.A1(n_3571),
.A2(n_3522),
.B1(n_3483),
.B2(n_3506),
.C(n_3505),
.Y(n_3631)
);

NAND3xp33_ASAP7_75t_L g3632 ( 
.A(n_3590),
.B(n_3486),
.C(n_3406),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3542),
.B(n_3447),
.Y(n_3633)
);

OAI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3578),
.A2(n_3478),
.B1(n_3442),
.B2(n_3438),
.Y(n_3634)
);

NAND2x1_ASAP7_75t_L g3635 ( 
.A(n_3542),
.B(n_3473),
.Y(n_3635)
);

O2A1O1Ixp33_ASAP7_75t_L g3636 ( 
.A1(n_3527),
.A2(n_3477),
.B(n_3423),
.C(n_3467),
.Y(n_3636)
);

AOI211xp5_ASAP7_75t_L g3637 ( 
.A1(n_3576),
.A2(n_3479),
.B(n_3455),
.C(n_3457),
.Y(n_3637)
);

AOI221x1_ASAP7_75t_L g3638 ( 
.A1(n_3546),
.A2(n_3389),
.B1(n_3476),
.B2(n_3474),
.C(n_3437),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3555),
.A2(n_3436),
.B(n_3520),
.Y(n_3639)
);

OAI22xp5_ASAP7_75t_L g3640 ( 
.A1(n_3610),
.A2(n_3426),
.B1(n_3393),
.B2(n_3381),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3565),
.B(n_3470),
.Y(n_3641)
);

OAI211xp5_ASAP7_75t_SL g3642 ( 
.A1(n_3611),
.A2(n_3446),
.B(n_3493),
.C(n_3433),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_SL g3643 ( 
.A(n_3594),
.B(n_3466),
.Y(n_3643)
);

NAND4xp25_ASAP7_75t_L g3644 ( 
.A(n_3593),
.B(n_3468),
.C(n_3440),
.D(n_3464),
.Y(n_3644)
);

OAI22xp5_ASAP7_75t_L g3645 ( 
.A1(n_3538),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_3645)
);

NOR3xp33_ASAP7_75t_L g3646 ( 
.A(n_3620),
.B(n_576),
.C(n_577),
.Y(n_3646)
);

NAND2xp33_ASAP7_75t_L g3647 ( 
.A(n_3540),
.B(n_578),
.Y(n_3647)
);

AOI221xp5_ASAP7_75t_L g3648 ( 
.A1(n_3563),
.A2(n_578),
.B1(n_579),
.B2(n_580),
.C(n_581),
.Y(n_3648)
);

AOI221xp5_ASAP7_75t_L g3649 ( 
.A1(n_3583),
.A2(n_579),
.B1(n_580),
.B2(n_583),
.C(n_584),
.Y(n_3649)
);

NAND3xp33_ASAP7_75t_SL g3650 ( 
.A(n_3581),
.B(n_585),
.C(n_586),
.Y(n_3650)
);

A2O1A1Ixp33_ASAP7_75t_L g3651 ( 
.A1(n_3570),
.A2(n_588),
.B(n_585),
.C(n_587),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3544),
.B(n_3614),
.Y(n_3652)
);

OAI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3537),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3536),
.B(n_765),
.Y(n_3654)
);

OAI211xp5_ASAP7_75t_SL g3655 ( 
.A1(n_3569),
.A2(n_591),
.B(n_589),
.C(n_590),
.Y(n_3655)
);

AOI21xp33_ASAP7_75t_SL g3656 ( 
.A1(n_3532),
.A2(n_591),
.B(n_592),
.Y(n_3656)
);

OAI211xp5_ASAP7_75t_L g3657 ( 
.A1(n_3545),
.A2(n_592),
.B(n_594),
.C(n_595),
.Y(n_3657)
);

AOI221xp5_ASAP7_75t_L g3658 ( 
.A1(n_3595),
.A2(n_595),
.B1(n_596),
.B2(n_597),
.C(n_598),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3580),
.A2(n_596),
.B(n_598),
.Y(n_3659)
);

AOI221x1_ASAP7_75t_L g3660 ( 
.A1(n_3547),
.A2(n_599),
.B1(n_600),
.B2(n_604),
.C(n_605),
.Y(n_3660)
);

AND2x2_ASAP7_75t_L g3661 ( 
.A(n_3612),
.B(n_599),
.Y(n_3661)
);

AOI221xp5_ASAP7_75t_L g3662 ( 
.A1(n_3582),
.A2(n_600),
.B1(n_604),
.B2(n_606),
.C(n_607),
.Y(n_3662)
);

NAND3xp33_ASAP7_75t_L g3663 ( 
.A(n_3549),
.B(n_606),
.C(n_607),
.Y(n_3663)
);

AOI221xp5_ASAP7_75t_L g3664 ( 
.A1(n_3587),
.A2(n_608),
.B1(n_609),
.B2(n_611),
.C(n_612),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3598),
.B(n_764),
.Y(n_3665)
);

A2O1A1Ixp33_ASAP7_75t_L g3666 ( 
.A1(n_3530),
.A2(n_608),
.B(n_609),
.C(n_613),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_SL g3667 ( 
.A(n_3596),
.B(n_614),
.Y(n_3667)
);

AOI221xp5_ASAP7_75t_L g3668 ( 
.A1(n_3589),
.A2(n_614),
.B1(n_615),
.B2(n_616),
.C(n_618),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3548),
.Y(n_3669)
);

INVxp67_ASAP7_75t_L g3670 ( 
.A(n_3562),
.Y(n_3670)
);

NAND5xp2_ASAP7_75t_SL g3671 ( 
.A(n_3574),
.B(n_615),
.C(n_620),
.D(n_621),
.E(n_622),
.Y(n_3671)
);

OAI31xp33_ASAP7_75t_L g3672 ( 
.A1(n_3575),
.A2(n_3551),
.A3(n_3535),
.B(n_3599),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3561),
.A2(n_620),
.B(n_621),
.Y(n_3673)
);

AOI211x1_ASAP7_75t_L g3674 ( 
.A1(n_3608),
.A2(n_622),
.B(n_623),
.C(n_626),
.Y(n_3674)
);

OAI21xp33_ASAP7_75t_L g3675 ( 
.A1(n_3579),
.A2(n_626),
.B(n_627),
.Y(n_3675)
);

A2O1A1Ixp33_ASAP7_75t_L g3676 ( 
.A1(n_3554),
.A2(n_3558),
.B(n_3597),
.C(n_3619),
.Y(n_3676)
);

OAI211xp5_ASAP7_75t_SL g3677 ( 
.A1(n_3533),
.A2(n_628),
.B(n_629),
.C(n_630),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_3550),
.Y(n_3678)
);

OAI22xp33_ASAP7_75t_L g3679 ( 
.A1(n_3577),
.A2(n_764),
.B1(n_629),
.B2(n_631),
.Y(n_3679)
);

OAI221xp5_ASAP7_75t_L g3680 ( 
.A1(n_3572),
.A2(n_628),
.B1(n_632),
.B2(n_634),
.C(n_635),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3534),
.B(n_632),
.Y(n_3681)
);

AOI221x1_ASAP7_75t_L g3682 ( 
.A1(n_3559),
.A2(n_634),
.B1(n_636),
.B2(n_637),
.C(n_638),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3602),
.B(n_763),
.Y(n_3683)
);

A2O1A1Ixp33_ASAP7_75t_SL g3684 ( 
.A1(n_3669),
.A2(n_3609),
.B(n_3601),
.C(n_3606),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3635),
.Y(n_3685)
);

AOI221xp5_ASAP7_75t_L g3686 ( 
.A1(n_3626),
.A2(n_3567),
.B1(n_3603),
.B2(n_3617),
.C(n_3604),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3661),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3654),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3674),
.Y(n_3689)
);

INVxp67_ASAP7_75t_L g3690 ( 
.A(n_3641),
.Y(n_3690)
);

OA22x2_ASAP7_75t_L g3691 ( 
.A1(n_3629),
.A2(n_3615),
.B1(n_3591),
.B2(n_3573),
.Y(n_3691)
);

AOI221xp5_ASAP7_75t_L g3692 ( 
.A1(n_3621),
.A2(n_3566),
.B1(n_3588),
.B2(n_3584),
.C(n_3585),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3665),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3670),
.Y(n_3694)
);

OAI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3678),
.A2(n_3541),
.B1(n_3531),
.B2(n_3557),
.Y(n_3695)
);

AO22x2_ASAP7_75t_L g3696 ( 
.A1(n_3632),
.A2(n_3618),
.B1(n_3613),
.B2(n_3592),
.Y(n_3696)
);

AO22x1_ASAP7_75t_SL g3697 ( 
.A1(n_3628),
.A2(n_3600),
.B1(n_638),
.B2(n_639),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3681),
.Y(n_3698)
);

AOI22xp5_ASAP7_75t_L g3699 ( 
.A1(n_3630),
.A2(n_637),
.B1(n_640),
.B2(n_641),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3625),
.Y(n_3700)
);

AOI22xp33_ASAP7_75t_L g3701 ( 
.A1(n_3646),
.A2(n_640),
.B1(n_641),
.B2(n_642),
.Y(n_3701)
);

HB1xp67_ASAP7_75t_L g3702 ( 
.A(n_3671),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3623),
.Y(n_3703)
);

OAI22x1_ASAP7_75t_L g3704 ( 
.A1(n_3663),
.A2(n_642),
.B1(n_644),
.B2(n_645),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3652),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3633),
.Y(n_3706)
);

INVxp67_ASAP7_75t_L g3707 ( 
.A(n_3667),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3660),
.Y(n_3708)
);

AOI221xp5_ASAP7_75t_L g3709 ( 
.A1(n_3656),
.A2(n_644),
.B1(n_646),
.B2(n_647),
.C(n_648),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3682),
.Y(n_3710)
);

INVx2_ASAP7_75t_SL g3711 ( 
.A(n_3643),
.Y(n_3711)
);

INVxp67_ASAP7_75t_L g3712 ( 
.A(n_3650),
.Y(n_3712)
);

AOI31xp33_ASAP7_75t_L g3713 ( 
.A1(n_3631),
.A2(n_648),
.A3(n_649),
.B(n_650),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3634),
.Y(n_3714)
);

OAI22xp5_ASAP7_75t_L g3715 ( 
.A1(n_3680),
.A2(n_649),
.B1(n_651),
.B2(n_652),
.Y(n_3715)
);

OAI22xp5_ASAP7_75t_L g3716 ( 
.A1(n_3666),
.A2(n_651),
.B1(n_652),
.B2(n_653),
.Y(n_3716)
);

O2A1O1Ixp33_ASAP7_75t_SL g3717 ( 
.A1(n_3651),
.A2(n_653),
.B(n_654),
.C(n_655),
.Y(n_3717)
);

INVxp67_ASAP7_75t_SL g3718 ( 
.A(n_3636),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3683),
.Y(n_3719)
);

AO22x2_ASAP7_75t_L g3720 ( 
.A1(n_3638),
.A2(n_654),
.B1(n_656),
.B2(n_657),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3677),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3711),
.B(n_3673),
.Y(n_3722)
);

AOI211xp5_ASAP7_75t_L g3723 ( 
.A1(n_3690),
.A2(n_3622),
.B(n_3675),
.C(n_3644),
.Y(n_3723)
);

AOI21xp33_ASAP7_75t_L g3724 ( 
.A1(n_3708),
.A2(n_3672),
.B(n_3647),
.Y(n_3724)
);

NOR3xp33_ASAP7_75t_L g3725 ( 
.A(n_3685),
.B(n_3624),
.C(n_3642),
.Y(n_3725)
);

NAND3xp33_ASAP7_75t_L g3726 ( 
.A(n_3714),
.B(n_3668),
.C(n_3664),
.Y(n_3726)
);

AOI211xp5_ASAP7_75t_SL g3727 ( 
.A1(n_3713),
.A2(n_3639),
.B(n_3679),
.C(n_3637),
.Y(n_3727)
);

AOI221xp5_ASAP7_75t_L g3728 ( 
.A1(n_3700),
.A2(n_3640),
.B1(n_3676),
.B2(n_3627),
.C(n_3659),
.Y(n_3728)
);

AOI22x1_ASAP7_75t_L g3729 ( 
.A1(n_3694),
.A2(n_3649),
.B1(n_3657),
.B2(n_3662),
.Y(n_3729)
);

AOI222xp33_ASAP7_75t_L g3730 ( 
.A1(n_3710),
.A2(n_3653),
.B1(n_3655),
.B2(n_3645),
.C1(n_3648),
.C2(n_3658),
.Y(n_3730)
);

O2A1O1Ixp33_ASAP7_75t_L g3731 ( 
.A1(n_3684),
.A2(n_656),
.B(n_657),
.C(n_658),
.Y(n_3731)
);

AOI221xp5_ASAP7_75t_L g3732 ( 
.A1(n_3693),
.A2(n_659),
.B1(n_661),
.B2(n_662),
.C(n_663),
.Y(n_3732)
);

A2O1A1Ixp33_ASAP7_75t_L g3733 ( 
.A1(n_3703),
.A2(n_661),
.B(n_662),
.C(n_663),
.Y(n_3733)
);

NOR3xp33_ASAP7_75t_SL g3734 ( 
.A(n_3695),
.B(n_762),
.C(n_664),
.Y(n_3734)
);

NOR3xp33_ASAP7_75t_L g3735 ( 
.A(n_3718),
.B(n_3705),
.C(n_3706),
.Y(n_3735)
);

NAND4xp75_ASAP7_75t_L g3736 ( 
.A(n_3686),
.B(n_664),
.C(n_665),
.D(n_666),
.Y(n_3736)
);

INVx2_ASAP7_75t_SL g3737 ( 
.A(n_3720),
.Y(n_3737)
);

AOI22xp5_ASAP7_75t_L g3738 ( 
.A1(n_3698),
.A2(n_665),
.B1(n_666),
.B2(n_667),
.Y(n_3738)
);

OAI211xp5_ASAP7_75t_L g3739 ( 
.A1(n_3712),
.A2(n_669),
.B(n_670),
.C(n_671),
.Y(n_3739)
);

HB1xp67_ASAP7_75t_L g3740 ( 
.A(n_3702),
.Y(n_3740)
);

AOI221xp5_ASAP7_75t_SL g3741 ( 
.A1(n_3731),
.A2(n_3707),
.B1(n_3692),
.B2(n_3721),
.C(n_3689),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3737),
.Y(n_3742)
);

A2O1A1Ixp33_ASAP7_75t_L g3743 ( 
.A1(n_3740),
.A2(n_3699),
.B(n_3719),
.C(n_3687),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3722),
.Y(n_3744)
);

AOI221xp5_ASAP7_75t_L g3745 ( 
.A1(n_3724),
.A2(n_3720),
.B1(n_3696),
.B2(n_3688),
.C(n_3717),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3736),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_3735),
.B(n_3696),
.Y(n_3747)
);

O2A1O1Ixp33_ASAP7_75t_L g3748 ( 
.A1(n_3725),
.A2(n_3715),
.B(n_3716),
.C(n_3701),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_L g3749 ( 
.A1(n_3729),
.A2(n_3691),
.B1(n_3704),
.B2(n_3709),
.Y(n_3749)
);

AOI322xp5_ASAP7_75t_L g3750 ( 
.A1(n_3728),
.A2(n_3697),
.A3(n_671),
.B1(n_672),
.B2(n_673),
.C1(n_674),
.C2(n_677),
.Y(n_3750)
);

NOR3xp33_ASAP7_75t_L g3751 ( 
.A(n_3723),
.B(n_669),
.C(n_677),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3734),
.B(n_678),
.Y(n_3752)
);

AOI221xp5_ASAP7_75t_L g3753 ( 
.A1(n_3726),
.A2(n_678),
.B1(n_679),
.B2(n_680),
.C(n_681),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3747),
.B(n_3727),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3752),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3742),
.Y(n_3756)
);

OAI21xp5_ASAP7_75t_L g3757 ( 
.A1(n_3750),
.A2(n_3730),
.B(n_3739),
.Y(n_3757)
);

AND2x4_ASAP7_75t_L g3758 ( 
.A(n_3744),
.B(n_3733),
.Y(n_3758)
);

NAND3xp33_ASAP7_75t_SL g3759 ( 
.A(n_3745),
.B(n_3732),
.C(n_3738),
.Y(n_3759)
);

AOI21xp33_ASAP7_75t_L g3760 ( 
.A1(n_3748),
.A2(n_3741),
.B(n_3749),
.Y(n_3760)
);

OAI221xp5_ASAP7_75t_SL g3761 ( 
.A1(n_3743),
.A2(n_762),
.B1(n_680),
.B2(n_681),
.C(n_682),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3746),
.B(n_679),
.Y(n_3762)
);

NOR3xp33_ASAP7_75t_L g3763 ( 
.A(n_3751),
.B(n_682),
.C(n_683),
.Y(n_3763)
);

NAND4xp25_ASAP7_75t_L g3764 ( 
.A(n_3760),
.B(n_3753),
.C(n_684),
.D(n_685),
.Y(n_3764)
);

NOR2xp67_ASAP7_75t_L g3765 ( 
.A(n_3756),
.B(n_3754),
.Y(n_3765)
);

AOI211xp5_ASAP7_75t_SL g3766 ( 
.A1(n_3761),
.A2(n_3759),
.B(n_3758),
.C(n_3762),
.Y(n_3766)
);

AND2x4_ASAP7_75t_L g3767 ( 
.A(n_3755),
.B(n_3757),
.Y(n_3767)
);

XOR2xp5_ASAP7_75t_L g3768 ( 
.A(n_3763),
.B(n_683),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3765),
.Y(n_3769)
);

NAND4xp25_ASAP7_75t_SL g3770 ( 
.A(n_3766),
.B(n_687),
.C(n_689),
.D(n_690),
.Y(n_3770)
);

AND5x1_ASAP7_75t_L g3771 ( 
.A(n_3764),
.B(n_687),
.C(n_689),
.D(n_691),
.E(n_693),
.Y(n_3771)
);

INVxp67_ASAP7_75t_SL g3772 ( 
.A(n_3769),
.Y(n_3772)
);

AOI22xp5_ASAP7_75t_L g3773 ( 
.A1(n_3772),
.A2(n_3767),
.B1(n_3770),
.B2(n_3768),
.Y(n_3773)
);

OAI31xp33_ASAP7_75t_SL g3774 ( 
.A1(n_3773),
.A2(n_3771),
.A3(n_693),
.B(n_695),
.Y(n_3774)
);

AOI211xp5_ASAP7_75t_L g3775 ( 
.A1(n_3774),
.A2(n_691),
.B(n_695),
.C(n_697),
.Y(n_3775)
);

AOI22xp33_ASAP7_75t_L g3776 ( 
.A1(n_3775),
.A2(n_698),
.B1(n_701),
.B2(n_702),
.Y(n_3776)
);

OAI22xp5_ASAP7_75t_SL g3777 ( 
.A1(n_3776),
.A2(n_698),
.B1(n_701),
.B2(n_702),
.Y(n_3777)
);

OR2x6_ASAP7_75t_L g3778 ( 
.A(n_3777),
.B(n_703),
.Y(n_3778)
);

AO21x2_ASAP7_75t_L g3779 ( 
.A1(n_3778),
.A2(n_703),
.B(n_704),
.Y(n_3779)
);

AOI222xp33_ASAP7_75t_L g3780 ( 
.A1(n_3778),
.A2(n_705),
.B1(n_706),
.B2(n_707),
.C1(n_708),
.C2(n_709),
.Y(n_3780)
);

AND2x2_ASAP7_75t_SL g3781 ( 
.A(n_3779),
.B(n_706),
.Y(n_3781)
);

OR2x2_ASAP7_75t_L g3782 ( 
.A(n_3780),
.B(n_710),
.Y(n_3782)
);

OR2x6_ASAP7_75t_L g3783 ( 
.A(n_3782),
.B(n_710),
.Y(n_3783)
);

AOI221xp5_ASAP7_75t_L g3784 ( 
.A1(n_3783),
.A2(n_3781),
.B1(n_712),
.B2(n_713),
.C(n_714),
.Y(n_3784)
);

AOI211xp5_ASAP7_75t_L g3785 ( 
.A1(n_3784),
.A2(n_711),
.B(n_712),
.C(n_715),
.Y(n_3785)
);


endmodule