module fake_netlist_5_917_n_2391 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2391);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2391;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_901;
wire n_553;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_857;
wire n_832;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_2022;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_604;
wire n_368;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_703;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_386;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2044;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_142),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_97),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_145),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_203),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_120),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_53),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_179),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_125),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_115),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_68),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_164),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_20),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_86),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_64),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_202),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_53),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_81),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_32),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_98),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_18),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_129),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_110),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_13),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_55),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_32),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_57),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_209),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_133),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_86),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_117),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_71),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_181),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_4),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_178),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_135),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_27),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_10),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_170),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_85),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_160),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_3),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_182),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_25),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_171),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_226),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_87),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_17),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_162),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_21),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_235),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_42),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_163),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_183),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_138),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_56),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_230),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_70),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_137),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_26),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_28),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_200),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_141),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_81),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_48),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_40),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_113),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_69),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_9),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_66),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_227),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_38),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_77),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_131),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_75),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_94),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_14),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_148),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_150),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_118),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_132),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_82),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_75),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_5),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_144),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_121),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_33),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_221),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_109),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_201),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_77),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_7),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_73),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_136),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_197),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_234),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_52),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_92),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_124),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_76),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_73),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_83),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_175),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_49),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_106),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_69),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_22),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_50),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_172),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_13),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_207),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_99),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_25),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_23),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_232),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_146),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_134),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_88),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_191),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_112),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_128),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_49),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_70),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_156),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_177),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_63),
.Y(n_379)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_154),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_54),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_213),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_123),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_12),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_83),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_102),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_84),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_33),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_42),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_122),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_218),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_108),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_195),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_152),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_52),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_63),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_35),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_62),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_85),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_48),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_119),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_68),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_56),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_30),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_187),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_55),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_8),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_228),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_24),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_237),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_8),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_212),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_22),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_216),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_67),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_130),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_71),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_67),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_149),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_31),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_50),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_76),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_62),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_26),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_19),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_51),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_180),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_6),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_196),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_127),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_103),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_14),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_114),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_15),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_40),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_211),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_9),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_10),
.Y(n_438)
);

BUFx8_ASAP7_75t_SL g439 ( 
.A(n_151),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_111),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_66),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_192),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_193),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_168),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_158),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_204),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_186),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_169),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_157),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_167),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_23),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_29),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_90),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_30),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_60),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_100),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_79),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_147),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_7),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_224),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_236),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_0),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_18),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_36),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_231),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_74),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_43),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_365),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_439),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_365),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_365),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_359),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_404),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_332),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_286),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_351),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_286),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_312),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_246),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_257),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_239),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_351),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_333),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_241),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_312),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_349),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_242),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_309),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_349),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_243),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_244),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_250),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_269),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_360),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_377),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_266),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_417),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_271),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_417),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_359),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_380),
.Y(n_511)
);

INVxp33_ASAP7_75t_SL g512 ( 
.A(n_466),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_380),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_319),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_428),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_416),
.Y(n_519)
);

INVxp33_ASAP7_75t_SL g520 ( 
.A(n_466),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_272),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_282),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_377),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_293),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_434),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_293),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_333),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_293),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_265),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_245),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_245),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_248),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_380),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_248),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_255),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_255),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_333),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_285),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_258),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_258),
.Y(n_541)
);

INVxp33_ASAP7_75t_SL g542 ( 
.A(n_251),
.Y(n_542)
);

BUFx2_ASAP7_75t_SL g543 ( 
.A(n_263),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_270),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_392),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_380),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_270),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_283),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_305),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_283),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_288),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_288),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_299),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_299),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_316),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_316),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_392),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_318),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_342),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_318),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_294),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_329),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_329),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_339),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_336),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_346),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_296),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_339),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_297),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_344),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_344),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_352),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_352),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_246),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_354),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_354),
.Y(n_576)
);

INVxp33_ASAP7_75t_SL g577 ( 
.A(n_254),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_300),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_380),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_336),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_303),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_388),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_388),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_249),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_399),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_307),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_311),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_314),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_323),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_399),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_407),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_407),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_418),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_413),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_418),
.Y(n_595)
);

INVxp33_ASAP7_75t_SL g596 ( 
.A(n_256),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_487),
.B(n_413),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_491),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_489),
.B(n_263),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_493),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_530),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_497),
.B(n_331),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_528),
.B(n_301),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_468),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_500),
.B(n_331),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_574),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_501),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_530),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_468),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_565),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_502),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_488),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_545),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_530),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_478),
.B(n_259),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_470),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_470),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_475),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_475),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_491),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_542),
.B(n_373),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_471),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_530),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_506),
.B(n_373),
.Y(n_625)
);

NOR2x1_ASAP7_75t_L g626 ( 
.A(n_471),
.B(n_240),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_508),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_472),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_584),
.B(n_450),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_472),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_473),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_473),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_474),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_476),
.Y(n_635)
);

AND2x2_ASAP7_75t_SL g636 ( 
.A(n_594),
.B(n_265),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_538),
.B(n_301),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_476),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_531),
.B(n_450),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_477),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_521),
.B(n_240),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_532),
.B(n_252),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_492),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_557),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_527),
.B(n_400),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_479),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_479),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_522),
.B(n_252),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_539),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_565),
.Y(n_651)
);

OA21x2_ASAP7_75t_L g652 ( 
.A1(n_480),
.A2(n_253),
.B(n_249),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_561),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_480),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_527),
.B(n_400),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_482),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_482),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_533),
.B(n_302),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_535),
.B(n_302),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_536),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_512),
.A2(n_409),
.B1(n_423),
.B2(n_274),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_569),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_536),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_524),
.B(n_325),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_492),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_537),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_537),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_495),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_578),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_495),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g671 ( 
.A1(n_520),
.A2(n_503),
.B1(n_516),
.B2(n_498),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_577),
.B(n_247),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_511),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_515),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_581),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_586),
.B(n_315),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_515),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_534),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_540),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_529),
.B(n_315),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_534),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_580),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_540),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_541),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_529),
.B(n_328),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_546),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_579),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_579),
.Y(n_691)
);

AND2x2_ASAP7_75t_SL g692 ( 
.A(n_524),
.B(n_265),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_541),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_483),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_544),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_672),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_629),
.B(n_587),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_672),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_SL g699 ( 
.A(n_664),
.B(n_566),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_601),
.Y(n_700)
);

BUFx10_ASAP7_75t_L g701 ( 
.A(n_674),
.Y(n_701)
);

AND3x2_ASAP7_75t_L g702 ( 
.A(n_622),
.B(n_374),
.C(n_317),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_601),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_619),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_636),
.B(n_588),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_672),
.Y(n_706)
);

NOR2x1p5_ASAP7_75t_L g707 ( 
.A(n_664),
.B(n_469),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_672),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_665),
.Y(n_709)
);

AND3x1_ASAP7_75t_L g710 ( 
.A(n_604),
.B(n_454),
.C(n_425),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_673),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_668),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_619),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_668),
.Y(n_714)
);

AO21x2_ASAP7_75t_L g715 ( 
.A1(n_641),
.A2(n_262),
.B(n_253),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_673),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_668),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_679),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_636),
.B(n_589),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_601),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_598),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_679),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_601),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_636),
.B(n_596),
.Y(n_724)
);

INVx8_ASAP7_75t_L g725 ( 
.A(n_629),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_613),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_604),
.B(n_484),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_616),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_679),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_601),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_599),
.B(n_567),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_619),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_629),
.B(n_649),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_620),
.Y(n_734)
);

BUFx4f_ASAP7_75t_L g735 ( 
.A(n_692),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_680),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_680),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_620),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_692),
.B(n_549),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_601),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_620),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_609),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_680),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_600),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_683),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_683),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_692),
.B(n_549),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_608),
.B(n_490),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_683),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_688),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_688),
.Y(n_751)
);

AO21x2_ASAP7_75t_L g752 ( 
.A1(n_678),
.A2(n_273),
.B(n_262),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_665),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_637),
.B(n_523),
.C(n_505),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_629),
.B(n_481),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_665),
.Y(n_756)
);

BUFx6f_ASAP7_75t_SL g757 ( 
.A(n_598),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_688),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_612),
.B(n_627),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_690),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_650),
.B(n_559),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_690),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_637),
.B(n_265),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_690),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_598),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_605),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_602),
.B(n_543),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_611),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_605),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_677),
.B(n_510),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_621),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_682),
.A2(n_543),
.B1(n_504),
.B2(n_454),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_610),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_610),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_617),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_617),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_606),
.B(n_265),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_618),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_630),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_618),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_625),
.B(n_281),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_630),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_621),
.B(n_306),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_623),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_623),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_265),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_628),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_609),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_651),
.B(n_519),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_635),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_684),
.B(n_554),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_635),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_607),
.A2(n_384),
.B1(n_389),
.B2(n_343),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_609),
.Y(n_796)
);

CKINVDCx6p67_ASAP7_75t_R g797 ( 
.A(n_597),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_614),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_645),
.B(n_291),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_621),
.B(n_305),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_614),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_628),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_638),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_609),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_609),
.Y(n_805)
);

AND3x2_ASAP7_75t_L g806 ( 
.A(n_653),
.B(n_369),
.C(n_328),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_662),
.B(n_558),
.Y(n_807)
);

INVxp33_ASAP7_75t_L g808 ( 
.A(n_661),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_652),
.B(n_275),
.C(n_273),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_638),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_669),
.A2(n_335),
.B1(n_261),
.B2(n_264),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_609),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_639),
.B(n_393),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_631),
.Y(n_814)
);

INVx5_ASAP7_75t_L g815 ( 
.A(n_665),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_638),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_640),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_655),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_631),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_633),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_639),
.A2(n_267),
.B1(n_268),
.B2(n_260),
.Y(n_821)
);

INVxp67_ASAP7_75t_SL g822 ( 
.A(n_665),
.Y(n_822)
);

AND2x6_ASAP7_75t_L g823 ( 
.A(n_639),
.B(n_291),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_682),
.B(n_275),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_640),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_652),
.B(n_278),
.C(n_276),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_633),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_639),
.B(n_665),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_640),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_615),
.Y(n_830)
);

BUFx10_ASAP7_75t_L g831 ( 
.A(n_642),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_655),
.B(n_305),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_656),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_634),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_670),
.B(n_326),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_656),
.Y(n_836)
);

AND2x6_ASAP7_75t_L g837 ( 
.A(n_626),
.B(n_291),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_634),
.Y(n_838)
);

AO21x2_ASAP7_75t_L g839 ( 
.A1(n_647),
.A2(n_278),
.B(n_276),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_671),
.B(n_277),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_647),
.Y(n_841)
);

BUFx10_ASAP7_75t_L g842 ( 
.A(n_642),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_670),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_682),
.A2(n_425),
.B1(n_457),
.B2(n_429),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_648),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_615),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_670),
.B(n_330),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_670),
.B(n_337),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_SL g849 ( 
.A1(n_671),
.A2(n_385),
.B1(n_437),
.B2(n_426),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_656),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_670),
.B(n_338),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_682),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_648),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_657),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_657),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_694),
.Y(n_856)
);

OAI21xp33_ASAP7_75t_SL g857 ( 
.A1(n_660),
.A2(n_457),
.B(n_544),
.Y(n_857)
);

NOR2x1p5_ASAP7_75t_L g858 ( 
.A(n_660),
.B(n_279),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_694),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_733),
.B(n_284),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_R g861 ( 
.A(n_726),
.B(n_699),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_852),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_725),
.B(n_670),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_852),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_711),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_725),
.B(n_676),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_725),
.B(n_676),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_746),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_735),
.A2(n_287),
.B1(n_295),
.B2(n_280),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_725),
.B(n_676),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_725),
.B(n_696),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_828),
.Y(n_872)
);

O2A1O1Ixp5_ASAP7_75t_L g873 ( 
.A1(n_735),
.A2(n_687),
.B(n_658),
.C(n_659),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_735),
.A2(n_658),
.B1(n_659),
.B2(n_642),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_766),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_697),
.B(n_289),
.Y(n_876)
);

INVx8_ASAP7_75t_L g877 ( 
.A(n_757),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_696),
.B(n_676),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_SL g879 ( 
.A(n_809),
.B(n_291),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_698),
.B(n_676),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_698),
.B(n_676),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_706),
.B(n_708),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_818),
.B(n_644),
.Y(n_883)
);

INVx8_ASAP7_75t_L g884 ( 
.A(n_757),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_754),
.B(n_290),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_744),
.B(n_644),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_818),
.B(n_291),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_706),
.B(n_689),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_711),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_708),
.B(n_689),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_801),
.B(n_687),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_842),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_808),
.A2(n_287),
.B1(n_295),
.B2(n_280),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_771),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_801),
.B(n_687),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_746),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_782),
.B(n_727),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_766),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_754),
.B(n_292),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_727),
.B(n_689),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_858),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_739),
.A2(n_429),
.B(n_369),
.C(n_687),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_767),
.B(n_689),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_842),
.B(n_291),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_769),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_749),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_749),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_842),
.B(n_436),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_769),
.B(n_689),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_773),
.B(n_774),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_750),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_793),
.B(n_663),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_705),
.B(n_298),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_716),
.B(n_663),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_774),
.B(n_689),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_750),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_809),
.A2(n_652),
.B1(n_341),
.B2(n_348),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_842),
.B(n_436),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_L g919 ( 
.A(n_807),
.B(n_308),
.C(n_304),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_701),
.B(n_666),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_751),
.Y(n_921)
);

INVx8_ASAP7_75t_L g922 ( 
.A(n_757),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_775),
.B(n_691),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_771),
.Y(n_924)
);

AO22x2_ASAP7_75t_L g925 ( 
.A1(n_747),
.A2(n_341),
.B1(n_348),
.B2(n_340),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_826),
.A2(n_652),
.B1(n_340),
.B2(n_382),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_765),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_831),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_719),
.B(n_310),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_831),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_SL g931 ( 
.A(n_707),
.B(n_313),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_831),
.B(n_436),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_775),
.B(n_691),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_728),
.B(n_436),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_776),
.B(n_691),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_776),
.B(n_691),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_858),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_778),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_701),
.B(n_666),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_724),
.B(n_320),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_751),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_778),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_781),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_781),
.B(n_691),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_755),
.B(n_436),
.Y(n_945)
);

INVx8_ASAP7_75t_L g946 ( 
.A(n_763),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_785),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_785),
.B(n_786),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_786),
.B(n_691),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_768),
.B(n_667),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_L g951 ( 
.A(n_770),
.B(n_322),
.C(n_321),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_789),
.B(n_643),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_826),
.A2(n_361),
.B1(n_383),
.B2(n_382),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_789),
.B(n_643),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_802),
.B(n_643),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_824),
.B(n_436),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_L g957 ( 
.A(n_731),
.B(n_667),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_802),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_814),
.B(n_643),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_814),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_819),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_758),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_819),
.B(n_675),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_791),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_820),
.B(n_675),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_839),
.A2(n_361),
.B1(n_390),
.B2(n_383),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_820),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_827),
.B(n_675),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_827),
.B(n_675),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_824),
.B(n_380),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_834),
.B(n_642),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_834),
.B(n_658),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_838),
.B(n_658),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_838),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_765),
.B(n_324),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_839),
.A2(n_401),
.B1(n_414),
.B2(n_390),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_758),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_841),
.B(n_659),
.Y(n_978)
);

NAND2x1_ASAP7_75t_L g979 ( 
.A(n_723),
.B(n_603),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_701),
.B(n_681),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_841),
.Y(n_981)
);

OR2x6_ASAP7_75t_L g982 ( 
.A(n_798),
.B(n_401),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_835),
.A2(n_615),
.B(n_603),
.Y(n_983)
);

OAI221xp5_ASAP7_75t_L g984 ( 
.A1(n_844),
.A2(n_695),
.B1(n_693),
.B2(n_686),
.C(n_685),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_811),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_845),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_824),
.B(n_380),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_845),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_824),
.B(n_659),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_813),
.B(n_681),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_854),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_SL g992 ( 
.A(n_707),
.B(n_327),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_710),
.A2(n_440),
.B1(n_449),
.B2(n_414),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_854),
.B(n_347),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_853),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_855),
.B(n_350),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_726),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_853),
.B(n_694),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_772),
.B(n_685),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_855),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_784),
.B(n_821),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_821),
.A2(n_449),
.B1(n_453),
.B2(n_440),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_721),
.B(n_334),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_715),
.B(n_752),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_760),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_712),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_712),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_710),
.B(n_355),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_744),
.B(n_686),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_704),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_857),
.A2(n_453),
.B(n_626),
.C(n_693),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_748),
.B(n_345),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_715),
.B(n_694),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_857),
.A2(n_695),
.B(n_548),
.C(n_550),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_715),
.B(n_694),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_752),
.B(n_694),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_752),
.B(n_603),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_714),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_856),
.B(n_357),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_763),
.B(n_603),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_760),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_763),
.B(n_624),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_763),
.B(n_624),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_761),
.B(n_353),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_832),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_714),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_856),
.B(n_363),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_763),
.B(n_624),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_806),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_763),
.B(n_624),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_763),
.B(n_822),
.Y(n_1031)
);

OAI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_797),
.A2(n_795),
.B1(n_356),
.B2(n_362),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_797),
.B(n_800),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_914),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_991),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_1001),
.A2(n_759),
.B1(n_849),
.B2(n_848),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_892),
.B(n_744),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_991),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_997),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_892),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_924),
.B(n_702),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_897),
.B(n_860),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_871),
.A2(n_753),
.B(n_709),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_892),
.B(n_859),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_1010),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1000),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_930),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_894),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_861),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_860),
.B(n_847),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_894),
.B(n_547),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_964),
.B(n_840),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_900),
.B(n_851),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1010),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_912),
.B(n_839),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1006),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_875),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_920),
.B(n_385),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_898),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_957),
.B(n_717),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1007),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_905),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1018),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_872),
.B(n_717),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_966),
.A2(n_823),
.B1(n_837),
.B2(n_777),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_892),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_930),
.B(n_859),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_938),
.Y(n_1068)
);

BUFx4f_ASAP7_75t_L g1069 ( 
.A(n_877),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_930),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_939),
.B(n_385),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_942),
.Y(n_1072)
);

INVx5_ASAP7_75t_L g1073 ( 
.A(n_946),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_966),
.A2(n_823),
.B1(n_837),
.B2(n_799),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_877),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_930),
.B(n_709),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_943),
.B(n_718),
.Y(n_1077)
);

AND2x6_ASAP7_75t_SL g1078 ( 
.A(n_982),
.B(n_547),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_718),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_980),
.B(n_1009),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_874),
.B(n_709),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_958),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_901),
.B(n_937),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_928),
.B(n_753),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_960),
.B(n_722),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_961),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_967),
.B(n_722),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_974),
.B(n_729),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_883),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_868),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_981),
.Y(n_1091)
);

AO22x1_ASAP7_75t_L g1092 ( 
.A1(n_913),
.A2(n_358),
.B1(n_375),
.B2(n_366),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_928),
.B(n_753),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_865),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_986),
.B(n_988),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_976),
.A2(n_823),
.B1(n_837),
.B2(n_788),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_989),
.B(n_756),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_995),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_976),
.A2(n_823),
.B1(n_837),
.B2(n_736),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_877),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_985),
.B(n_756),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_910),
.B(n_729),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1026),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_862),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_953),
.A2(n_823),
.B1(n_837),
.B2(n_737),
.Y(n_1105)
);

NAND2xp33_ASAP7_75t_L g1106 ( 
.A(n_946),
.B(n_823),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_913),
.A2(n_823),
.B1(n_843),
.B2(n_756),
.Y(n_1107)
);

NOR2x2_ASAP7_75t_L g1108 ( 
.A(n_891),
.B(n_385),
.Y(n_1108)
);

AND3x2_ASAP7_75t_SL g1109 ( 
.A(n_1002),
.B(n_869),
.C(n_893),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_864),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1004),
.B(n_843),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_896),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_948),
.B(n_736),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_884),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_953),
.A2(n_837),
.B1(n_743),
.B2(n_745),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_906),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_971),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_972),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_876),
.B(n_737),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_975),
.B(n_950),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_973),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_861),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_884),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_884),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_1033),
.B(n_548),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_907),
.Y(n_1126)
);

NOR2x2_ASAP7_75t_L g1127 ( 
.A(n_891),
.B(n_426),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_911),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_946),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_876),
.B(n_743),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_916),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_978),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_927),
.B(n_843),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_SL g1134 ( 
.A(n_1012),
.B(n_381),
.C(n_379),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_909),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_889),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_922),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_929),
.A2(n_745),
.B1(n_364),
.B2(n_368),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1029),
.B(n_550),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_922),
.B(n_551),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_891),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_921),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_873),
.B(n_700),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_922),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_941),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_915),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_990),
.B(n_762),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1003),
.B(n_762),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_927),
.B(n_723),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_929),
.B(n_940),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_895),
.B(n_551),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_895),
.Y(n_1152)
);

INVx5_ASAP7_75t_L g1153 ( 
.A(n_895),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_979),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_962),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_982),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_923),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_933),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_869),
.A2(n_837),
.B1(n_426),
.B2(n_437),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_977),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1005),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_935),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1003),
.B(n_764),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_936),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_944),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_982),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_949),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_885),
.B(n_764),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_931),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1012),
.A2(n_395),
.B1(n_396),
.B2(n_387),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1021),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_998),
.Y(n_1172)
);

OR2x6_ASAP7_75t_L g1173 ( 
.A(n_1025),
.B(n_552),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_882),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_885),
.B(n_723),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_999),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_952),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_899),
.B(n_730),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_989),
.B(n_552),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_975),
.B(n_899),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_940),
.B(n_730),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_903),
.B(n_730),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_878),
.Y(n_1183)
);

NOR2x1p5_ASAP7_75t_L g1184 ( 
.A(n_919),
.B(n_397),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_SL g1185 ( 
.A(n_1002),
.B(n_402),
.C(n_398),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_880),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1008),
.B(n_742),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_925),
.B(n_742),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_SL g1189 ( 
.A(n_1024),
.B(n_406),
.C(n_403),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_954),
.Y(n_1190)
);

BUFx12f_ASAP7_75t_L g1191 ( 
.A(n_886),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_955),
.Y(n_1192)
);

NAND2xp33_ASAP7_75t_L g1193 ( 
.A(n_917),
.B(n_700),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_863),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_959),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_881),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1008),
.B(n_742),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_879),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_951),
.B(n_553),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_963),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_994),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1024),
.A2(n_1014),
.B(n_993),
.C(n_1011),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1032),
.A2(n_415),
.B1(n_420),
.B2(n_411),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_965),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_888),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_925),
.B(n_796),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_994),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_968),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_925),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_917),
.B(n_796),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_926),
.B(n_796),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_893),
.A2(n_422),
.B1(n_432),
.B2(n_421),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_926),
.A2(n_367),
.B1(n_371),
.B2(n_370),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_970),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_866),
.A2(n_815),
.B(n_703),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_992),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_970),
.B(n_804),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_R g1218 ( 
.A(n_1017),
.B(n_372),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_890),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1013),
.B(n_700),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_987),
.B(n_553),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_996),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_996),
.Y(n_1223)
);

O2A1O1Ixp5_ASAP7_75t_L g1224 ( 
.A1(n_945),
.A2(n_804),
.B(n_846),
.C(n_805),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_L g1225 ( 
.A(n_902),
.B(n_700),
.Y(n_1225)
);

AND2x6_ASAP7_75t_SL g1226 ( 
.A(n_1032),
.B(n_555),
.Y(n_1226)
);

OR2x2_ASAP7_75t_SL g1227 ( 
.A(n_1015),
.B(n_555),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1053),
.A2(n_870),
.B(n_867),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1180),
.B(n_1019),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1215),
.A2(n_983),
.B(n_1016),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1080),
.B(n_1120),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1034),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1042),
.A2(n_987),
.B(n_887),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1056),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1056),
.Y(n_1235)
);

O2A1O1Ixp5_ASAP7_75t_L g1236 ( 
.A1(n_1150),
.A2(n_934),
.B(n_932),
.C(n_945),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1057),
.Y(n_1237)
);

AND2x2_ASAP7_75t_SL g1238 ( 
.A(n_1069),
.B(n_1031),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1193),
.A2(n_908),
.B(n_904),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1047),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1150),
.A2(n_984),
.B1(n_887),
.B2(n_934),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1047),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1176),
.B(n_1089),
.Y(n_1243)
);

AOI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1143),
.A2(n_1111),
.B(n_1044),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1059),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1061),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1062),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1173),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1061),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1063),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_1187),
.A2(n_932),
.B(n_908),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1173),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_SL g1253 ( 
.A1(n_1052),
.A2(n_969),
.B(n_805),
.C(n_830),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1047),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1050),
.A2(n_918),
.B(n_904),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1058),
.B(n_426),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1047),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1176),
.B(n_1019),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1117),
.B(n_918),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1036),
.A2(n_1027),
.B(n_956),
.C(n_1022),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1075),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1039),
.Y(n_1262)
);

XOR2xp5_ASAP7_75t_L g1263 ( 
.A(n_1049),
.B(n_1122),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1118),
.B(n_956),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1212),
.A2(n_1027),
.B(n_1023),
.C(n_1020),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1121),
.B(n_779),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1040),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1040),
.A2(n_1030),
.B(n_1028),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1222),
.A2(n_433),
.B1(n_376),
.B2(n_378),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1040),
.A2(n_815),
.B(n_703),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1202),
.A2(n_804),
.B(n_846),
.C(n_805),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1134),
.A2(n_305),
.B1(n_456),
.B2(n_448),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1132),
.B(n_779),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1212),
.A2(n_1189),
.B(n_1202),
.C(n_1052),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1209),
.A2(n_435),
.B1(n_438),
.B2(n_441),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_SL g1276 ( 
.A(n_1185),
.B(n_452),
.C(n_451),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1124),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1153),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1063),
.Y(n_1279)
);

O2A1O1Ixp5_ASAP7_75t_L g1280 ( 
.A1(n_1143),
.A2(n_850),
.B(n_780),
.C(n_836),
.Y(n_1280)
);

NAND2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1169),
.B(n_386),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1094),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1191),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1111),
.A2(n_783),
.B(n_780),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1040),
.A2(n_815),
.B(n_703),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1066),
.A2(n_815),
.B(n_703),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1048),
.B(n_556),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1153),
.Y(n_1288)
);

AOI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1044),
.A2(n_787),
.B(n_783),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1071),
.B(n_437),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1055),
.B(n_787),
.Y(n_1291)
);

AO22x1_ASAP7_75t_L g1292 ( 
.A1(n_1153),
.A2(n_455),
.B1(n_459),
.B2(n_462),
.Y(n_1292)
);

OR2x6_ASAP7_75t_L g1293 ( 
.A(n_1144),
.B(n_556),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1095),
.A2(n_575),
.B(n_560),
.C(n_562),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1103),
.Y(n_1295)
);

OA22x2_ASAP7_75t_L g1296 ( 
.A1(n_1203),
.A2(n_464),
.B1(n_463),
.B2(n_467),
.Y(n_1296)
);

XOR2xp5_ASAP7_75t_L g1297 ( 
.A(n_1216),
.B(n_391),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1068),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1129),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1223),
.A2(n_405),
.B1(n_394),
.B2(n_408),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1136),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1037),
.A2(n_582),
.B(n_560),
.C(n_562),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1173),
.B(n_1201),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_SL g1304 ( 
.A1(n_1187),
.A2(n_830),
.B(n_846),
.C(n_836),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1207),
.A2(n_410),
.B1(n_412),
.B2(n_465),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1175),
.A2(n_703),
.B(n_700),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_L g1307 ( 
.A(n_1185),
.B(n_427),
.C(n_419),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1151),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_1137),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1066),
.A2(n_815),
.B(n_740),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1153),
.B(n_430),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1051),
.B(n_1139),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1066),
.A2(n_815),
.B(n_740),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1051),
.B(n_437),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1174),
.B(n_792),
.Y(n_1315)
);

O2A1O1Ixp5_ASAP7_75t_L g1316 ( 
.A1(n_1178),
.A2(n_1197),
.B(n_1181),
.C(n_1130),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1101),
.B(n_1048),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1141),
.B(n_563),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1072),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1066),
.B(n_830),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1214),
.A2(n_1179),
.B1(n_1209),
.B2(n_1221),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1125),
.B(n_431),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1129),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1199),
.A2(n_442),
.B1(n_443),
.B2(n_444),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1139),
.B(n_563),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1082),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1178),
.A2(n_445),
.B(n_446),
.C(n_447),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1151),
.B(n_564),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_L g1329 ( 
.A(n_1092),
.B(n_460),
.C(n_458),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1174),
.B(n_792),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1101),
.B(n_461),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1129),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1075),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1100),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1156),
.B(n_720),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1166),
.B(n_720),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1156),
.B(n_720),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1166),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1179),
.B(n_720),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1043),
.A2(n_803),
.B(n_794),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_SL g1341 ( 
.A1(n_1197),
.A2(n_850),
.B(n_833),
.C(n_829),
.Y(n_1341)
);

O2A1O1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1037),
.A2(n_576),
.B(n_564),
.C(n_568),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1214),
.A2(n_833),
.B(n_829),
.C(n_825),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1224),
.A2(n_803),
.B(n_794),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1081),
.A2(n_720),
.B(n_740),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1100),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1138),
.A2(n_575),
.B(n_568),
.C(n_570),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1129),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1070),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1081),
.A2(n_740),
.B(n_790),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1170),
.B(n_740),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1209),
.A2(n_1115),
.B1(n_1099),
.B2(n_1074),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1209),
.A2(n_583),
.B1(n_570),
.B2(n_571),
.Y(n_1353)
);

O2A1O1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1147),
.A2(n_576),
.B(n_571),
.C(n_572),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1199),
.B(n_572),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1186),
.B(n_810),
.Y(n_1356)
);

OAI22x1_ASAP7_75t_L g1357 ( 
.A1(n_1109),
.A2(n_595),
.B1(n_593),
.B2(n_592),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1220),
.A2(n_825),
.B(n_817),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1168),
.A2(n_790),
.B(n_812),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1221),
.B(n_573),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1084),
.A2(n_1093),
.B(n_1220),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1188),
.A2(n_817),
.B(n_816),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1186),
.B(n_810),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1086),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1196),
.B(n_816),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1152),
.B(n_573),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1144),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1119),
.A2(n_812),
.B(n_790),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1196),
.B(n_704),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1091),
.B(n_790),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1098),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1103),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1046),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1104),
.B(n_582),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1148),
.A2(n_593),
.B(n_585),
.C(n_590),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1163),
.A2(n_595),
.B(n_585),
.C(n_590),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1133),
.B(n_790),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1133),
.B(n_812),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1084),
.A2(n_1093),
.B(n_1106),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1115),
.A2(n_583),
.B1(n_591),
.B2(n_592),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1182),
.A2(n_812),
.B(n_615),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1102),
.A2(n_812),
.B(n_615),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1177),
.A2(n_741),
.B(n_738),
.C(n_734),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1218),
.B(n_713),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1113),
.A2(n_615),
.B(n_738),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1149),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1064),
.A2(n_1219),
.B(n_1205),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1210),
.A2(n_741),
.B(n_734),
.Y(n_1388)
);

OA22x2_ASAP7_75t_L g1389 ( 
.A1(n_1109),
.A2(n_591),
.B1(n_485),
.B2(n_486),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1099),
.A2(n_514),
.B1(n_485),
.B2(n_486),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1045),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1226),
.B(n_0),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1114),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1149),
.B(n_1),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1205),
.B(n_713),
.Y(n_1395)
);

NOR3xp33_ASAP7_75t_SL g1396 ( 
.A(n_1213),
.B(n_483),
.C(n_494),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1110),
.B(n_1),
.Y(n_1397)
);

AOI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1284),
.A2(n_1067),
.B(n_1076),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_SL g1399 ( 
.A1(n_1274),
.A2(n_1206),
.B(n_1211),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1251),
.A2(n_1219),
.A3(n_1135),
.B(n_1164),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1344),
.A2(n_1067),
.B(n_1183),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1228),
.A2(n_1073),
.B(n_1076),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_SL g1403 ( 
.A(n_1261),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_SL g1404 ( 
.A(n_1392),
.B(n_1159),
.C(n_1218),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1316),
.A2(n_1079),
.B(n_1077),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1271),
.A2(n_1192),
.B(n_1190),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1237),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1340),
.A2(n_1183),
.B(n_1097),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1229),
.B(n_1172),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1352),
.B(n_1146),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1352),
.B(n_1157),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1255),
.A2(n_1073),
.B(n_1060),
.Y(n_1412)
);

AO31x2_ASAP7_75t_L g1413 ( 
.A1(n_1241),
.A2(n_1167),
.A3(n_1162),
.B(n_1158),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1333),
.Y(n_1414)
);

OAI22x1_ASAP7_75t_L g1415 ( 
.A1(n_1394),
.A2(n_1184),
.B1(n_1083),
.B2(n_1041),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1317),
.B(n_1165),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1289),
.A2(n_1097),
.B(n_1087),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1267),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1321),
.A2(n_1074),
.B1(n_1096),
.B2(n_1065),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1387),
.B(n_1195),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1236),
.A2(n_1204),
.B(n_1200),
.Y(n_1421)
);

INVxp67_ASAP7_75t_L g1422 ( 
.A(n_1232),
.Y(n_1422)
);

AOI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1357),
.A2(n_1159),
.B1(n_1041),
.B2(n_1083),
.C(n_1208),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1230),
.A2(n_1088),
.B(n_1085),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1312),
.B(n_1114),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1280),
.A2(n_1217),
.B(n_1070),
.Y(n_1426)
);

AO31x2_ASAP7_75t_L g1427 ( 
.A1(n_1241),
.A2(n_1038),
.A3(n_1035),
.B(n_1054),
.Y(n_1427)
);

OR2x2_ASAP7_75t_SL g1428 ( 
.A(n_1276),
.B(n_1108),
.Y(n_1428)
);

NOR4xp25_ASAP7_75t_L g1429 ( 
.A(n_1375),
.B(n_1110),
.C(n_1171),
.D(n_1225),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1387),
.B(n_1194),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1239),
.A2(n_1260),
.B(n_1233),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1386),
.B(n_1194),
.Y(n_1432)
);

NOR3xp33_ASAP7_75t_SL g1433 ( 
.A(n_1281),
.B(n_1127),
.C(n_1078),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1245),
.Y(n_1434)
);

AO31x2_ASAP7_75t_L g1435 ( 
.A1(n_1306),
.A2(n_1035),
.A3(n_1038),
.B(n_1054),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1379),
.A2(n_1073),
.B(n_1096),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1306),
.A2(n_1107),
.B(n_1112),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1367),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1244),
.A2(n_1155),
.B(n_1131),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1360),
.B(n_1194),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1291),
.A2(n_1073),
.B(n_1065),
.Y(n_1441)
);

NOR2xp67_ASAP7_75t_L g1442 ( 
.A(n_1301),
.B(n_1123),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1367),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1368),
.A2(n_1155),
.B(n_1128),
.Y(n_1444)
);

INVxp67_ASAP7_75t_SL g1445 ( 
.A(n_1242),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1282),
.Y(n_1446)
);

NAND2xp33_ASAP7_75t_L g1447 ( 
.A(n_1278),
.B(n_1288),
.Y(n_1447)
);

AOI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1258),
.A2(n_1116),
.B(n_1131),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1234),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1233),
.A2(n_1217),
.B(n_1145),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1247),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1231),
.B(n_1194),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1298),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1331),
.A2(n_1069),
.B(n_1105),
.C(n_1090),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1243),
.B(n_1140),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1389),
.A2(n_1105),
.B1(n_1227),
.B2(n_1198),
.Y(n_1456)
);

AOI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1389),
.A2(n_1142),
.B(n_1161),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1345),
.A2(n_1142),
.B(n_1161),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1355),
.B(n_1328),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1333),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1291),
.A2(n_1361),
.B(n_1259),
.Y(n_1461)
);

AO31x2_ASAP7_75t_L g1462 ( 
.A1(n_1343),
.A2(n_1045),
.A3(n_1112),
.B(n_1145),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1297),
.B(n_1140),
.Y(n_1463)
);

AO31x2_ASAP7_75t_L g1464 ( 
.A1(n_1368),
.A2(n_1116),
.A3(n_1126),
.B(n_1128),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1259),
.A2(n_1198),
.B(n_1126),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1275),
.A2(n_1140),
.B(n_1160),
.C(n_1123),
.Y(n_1466)
);

AO32x2_ASAP7_75t_L g1467 ( 
.A1(n_1353),
.A2(n_1198),
.A3(n_1160),
.B1(n_4),
.B2(n_6),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1235),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1333),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1383),
.A2(n_1198),
.B(n_732),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1367),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1246),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1249),
.B(n_1250),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1377),
.A2(n_1154),
.B(n_732),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1325),
.B(n_494),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1350),
.A2(n_514),
.B(n_526),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1378),
.A2(n_1154),
.B(n_654),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1279),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1264),
.A2(n_1154),
.B(n_654),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1304),
.A2(n_513),
.B(n_526),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1303),
.A2(n_1154),
.B1(n_517),
.B2(n_513),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1319),
.B(n_496),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1338),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1388),
.A2(n_1358),
.B(n_1359),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1265),
.A2(n_1388),
.B(n_1385),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1346),
.Y(n_1486)
);

AOI221x1_ASAP7_75t_L g1487 ( 
.A1(n_1397),
.A2(n_517),
.B1(n_499),
.B2(n_507),
.C(n_525),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1358),
.A2(n_496),
.B(n_525),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1262),
.B(n_2),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1308),
.B(n_499),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1295),
.B(n_507),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1326),
.Y(n_1492)
);

BUFx8_ASAP7_75t_L g1493 ( 
.A(n_1277),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1381),
.A2(n_509),
.B(n_518),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1372),
.B(n_509),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1346),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1264),
.A2(n_654),
.B(n_646),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1256),
.B(n_518),
.Y(n_1498)
);

AOI31xp67_ASAP7_75t_L g1499 ( 
.A1(n_1384),
.A2(n_654),
.A3(n_646),
.B(n_632),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1364),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1371),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1373),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1382),
.A2(n_166),
.B(n_91),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1391),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1315),
.A2(n_173),
.B(n_93),
.Y(n_1505)
);

AO31x2_ASAP7_75t_L g1506 ( 
.A1(n_1353),
.A2(n_3),
.A3(n_11),
.B(n_15),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1287),
.B(n_632),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1266),
.B(n_632),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1267),
.A2(n_654),
.B(n_646),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1315),
.A2(n_654),
.B(n_646),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1253),
.A2(n_174),
.B(n_95),
.Y(n_1511)
);

A2O1A1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1396),
.A2(n_646),
.B(n_632),
.C(n_19),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1268),
.A2(n_646),
.B(n_632),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1309),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1266),
.A2(n_632),
.B(n_223),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1273),
.A2(n_220),
.B(n_219),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1290),
.B(n_11),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1330),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1273),
.A2(n_215),
.B(n_214),
.Y(n_1519)
);

NAND2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1278),
.B(n_210),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1356),
.B(n_16),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1330),
.A2(n_206),
.B(n_199),
.Y(n_1522)
);

OAI22x1_ASAP7_75t_L g1523 ( 
.A1(n_1248),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1374),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1356),
.A2(n_194),
.B(n_190),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1369),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1366),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1363),
.A2(n_1365),
.B(n_1369),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1287),
.Y(n_1529)
);

OAI21xp33_ASAP7_75t_L g1530 ( 
.A1(n_1272),
.A2(n_24),
.B(n_27),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1252),
.B(n_28),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1363),
.A2(n_188),
.B(n_185),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1318),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1318),
.B(n_29),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1351),
.A2(n_184),
.B(n_176),
.Y(n_1535)
);

BUFx4f_ASAP7_75t_SL g1536 ( 
.A(n_1346),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1314),
.B(n_31),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1365),
.A2(n_165),
.B(n_161),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1395),
.A2(n_159),
.B(n_153),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1395),
.B(n_1238),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1362),
.Y(n_1541)
);

AOI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1362),
.A2(n_143),
.B(n_140),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1294),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1242),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1296),
.A2(n_1269),
.B1(n_1283),
.B2(n_1263),
.Y(n_1545)
);

AOI221x1_ASAP7_75t_L g1546 ( 
.A1(n_1327),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.C(n_37),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1349),
.B(n_34),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1270),
.A2(n_139),
.B(n_126),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1339),
.A2(n_116),
.B(n_107),
.Y(n_1549)
);

NOR2xp67_ASAP7_75t_L g1550 ( 
.A(n_1329),
.B(n_105),
.Y(n_1550)
);

NAND2x1_ASAP7_75t_L g1551 ( 
.A(n_1348),
.B(n_104),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1296),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1348),
.Y(n_1553)
);

CKINVDCx16_ASAP7_75t_R g1554 ( 
.A(n_1293),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1278),
.B(n_101),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1341),
.A2(n_96),
.B(n_89),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1349),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1285),
.A2(n_39),
.B(n_41),
.Y(n_1558)
);

OAI22x1_ASAP7_75t_L g1559 ( 
.A1(n_1335),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_1334),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1242),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1370),
.A2(n_44),
.B(n_45),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1324),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1275),
.B(n_46),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1302),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1376),
.A2(n_47),
.B(n_51),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1337),
.A2(n_54),
.B(n_57),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1286),
.A2(n_58),
.B(n_59),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1254),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1380),
.A2(n_58),
.A3(n_59),
.B(n_60),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1257),
.A2(n_61),
.B(n_64),
.Y(n_1571)
);

O2A1O1Ixp5_ASAP7_75t_L g1572 ( 
.A1(n_1311),
.A2(n_65),
.B(n_72),
.C(n_74),
.Y(n_1572)
);

AOI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1322),
.A2(n_65),
.B(n_72),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1310),
.A2(n_1313),
.B(n_1320),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1354),
.A2(n_1307),
.B(n_1347),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1336),
.B(n_1299),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1299),
.B(n_78),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1300),
.B(n_84),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1342),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1390),
.A2(n_78),
.B(n_79),
.Y(n_1580)
);

AO31x2_ASAP7_75t_L g1581 ( 
.A1(n_1390),
.A2(n_80),
.A3(n_82),
.B(n_1240),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1485),
.A2(n_1305),
.B(n_1393),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1440),
.B(n_1288),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1430),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1461),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1292),
.C(n_1293),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1408),
.A2(n_1323),
.B(n_1332),
.Y(n_1587)
);

AOI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1439),
.A2(n_1293),
.B(n_1288),
.Y(n_1588)
);

AOI21xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1415),
.A2(n_80),
.B(n_1323),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1431),
.A2(n_1254),
.B(n_1332),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1424),
.A2(n_1254),
.B(n_1402),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1530),
.A2(n_1404),
.B1(n_1566),
.B2(n_1580),
.C(n_1517),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1440),
.B(n_1409),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1500),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1580),
.A2(n_1566),
.B1(n_1564),
.B2(n_1578),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1458),
.A2(n_1401),
.B(n_1417),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1412),
.A2(n_1426),
.B(n_1398),
.Y(n_1597)
);

NOR2x1_ASAP7_75t_R g1598 ( 
.A(n_1514),
.B(n_1560),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1407),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1438),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1459),
.B(n_1475),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1416),
.B(n_1524),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1430),
.Y(n_1603)
);

AO21x2_ASAP7_75t_L g1604 ( 
.A1(n_1429),
.A2(n_1556),
.B(n_1421),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1535),
.B(n_1466),
.Y(n_1605)
);

AOI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1465),
.A2(n_1574),
.B(n_1448),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1554),
.A2(n_1419),
.B1(n_1463),
.B2(n_1489),
.Y(n_1607)
);

OAI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1497),
.A2(n_1513),
.B(n_1542),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1503),
.A2(n_1436),
.B(n_1476),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1434),
.Y(n_1610)
);

AOI21xp33_ASAP7_75t_SL g1611 ( 
.A1(n_1545),
.A2(n_1523),
.B(n_1455),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1416),
.B(n_1432),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1528),
.A2(n_1494),
.B(n_1479),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1575),
.A2(n_1421),
.B(n_1454),
.Y(n_1614)
);

AOI22x1_ASAP7_75t_L g1615 ( 
.A1(n_1559),
.A2(n_1543),
.B1(n_1562),
.B2(n_1575),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1546),
.A2(n_1419),
.B1(n_1411),
.B2(n_1410),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1451),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1527),
.B(n_1498),
.Y(n_1618)
);

AO31x2_ASAP7_75t_L g1619 ( 
.A1(n_1487),
.A2(n_1441),
.A3(n_1420),
.B(n_1456),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1429),
.A2(n_1556),
.B(n_1510),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1438),
.Y(n_1621)
);

CKINVDCx11_ASAP7_75t_R g1622 ( 
.A(n_1414),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1443),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1548),
.A2(n_1420),
.B(n_1450),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1510),
.A2(n_1450),
.B(n_1406),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1423),
.A2(n_1571),
.B1(n_1399),
.B2(n_1522),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1444),
.Y(n_1627)
);

AND2x6_ASAP7_75t_L g1628 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1522),
.A2(n_1537),
.B1(n_1456),
.B2(n_1529),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1444),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1526),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1567),
.A2(n_1531),
.B1(n_1533),
.B2(n_1534),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1529),
.B(n_1432),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1406),
.A2(n_1512),
.B(n_1481),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1428),
.A2(n_1425),
.B1(n_1446),
.B2(n_1520),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1505),
.A2(n_1488),
.B(n_1539),
.Y(n_1636)
);

INVx8_ASAP7_75t_L g1637 ( 
.A(n_1403),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1558),
.A2(n_1493),
.B1(n_1403),
.B2(n_1555),
.Y(n_1638)
);

OA21x2_ASAP7_75t_L g1639 ( 
.A1(n_1568),
.A2(n_1470),
.B(n_1525),
.Y(n_1639)
);

BUFx2_ASAP7_75t_SL g1640 ( 
.A(n_1442),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1532),
.A2(n_1538),
.B(n_1515),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1470),
.A2(n_1508),
.B(n_1540),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1518),
.B(n_1452),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1452),
.B(n_1540),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1558),
.A2(n_1565),
.B1(n_1579),
.B2(n_1521),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1563),
.A2(n_1572),
.B1(n_1422),
.B2(n_1453),
.C(n_1502),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1474),
.A2(n_1477),
.B(n_1521),
.Y(n_1647)
);

AO31x2_ASAP7_75t_L g1648 ( 
.A1(n_1508),
.A2(n_1499),
.A3(n_1547),
.B(n_1516),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1425),
.B(n_1490),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1483),
.A2(n_1576),
.B1(n_1492),
.B2(n_1501),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1437),
.A2(n_1484),
.B(n_1509),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1471),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1550),
.A2(n_1482),
.B1(n_1449),
.B2(n_1468),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1462),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1418),
.B(n_1553),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1462),
.Y(n_1656)
);

CKINVDCx6p67_ASAP7_75t_R g1657 ( 
.A(n_1414),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1437),
.A2(n_1484),
.B(n_1405),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1472),
.Y(n_1659)
);

CKINVDCx11_ASAP7_75t_R g1660 ( 
.A(n_1414),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1464),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1576),
.A2(n_1507),
.B1(n_1433),
.B2(n_1577),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1405),
.A2(n_1519),
.B(n_1495),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1520),
.B(n_1555),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1478),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1464),
.Y(n_1666)
);

AO31x2_ASAP7_75t_L g1667 ( 
.A1(n_1547),
.A2(n_1577),
.A3(n_1495),
.B(n_1413),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1473),
.A2(n_1460),
.B1(n_1496),
.B2(n_1553),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1464),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1557),
.B(n_1504),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1544),
.Y(n_1671)
);

OAI21x1_ASAP7_75t_L g1672 ( 
.A1(n_1519),
.A2(n_1573),
.B(n_1491),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_SL g1673 ( 
.A1(n_1549),
.A2(n_1457),
.B(n_1473),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1544),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1418),
.A2(n_1445),
.B1(n_1469),
.B2(n_1486),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1491),
.B(n_1486),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1469),
.B(n_1486),
.Y(n_1677)
);

INVx5_ASAP7_75t_L g1678 ( 
.A(n_1418),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1469),
.B(n_1569),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1551),
.A2(n_1435),
.B(n_1427),
.Y(n_1680)
);

OR2x6_ASAP7_75t_L g1681 ( 
.A(n_1544),
.B(n_1561),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1435),
.A2(n_1427),
.B(n_1480),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1506),
.B(n_1581),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1435),
.A2(n_1427),
.B(n_1480),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1457),
.A2(n_1467),
.B(n_1447),
.C(n_1418),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1467),
.A2(n_1561),
.B1(n_1570),
.B2(n_1506),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_SL g1687 ( 
.A(n_1467),
.B(n_1493),
.C(n_1570),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1561),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1400),
.A2(n_1413),
.B(n_1511),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_SL g1690 ( 
.A(n_1581),
.B(n_1570),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1511),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1400),
.A2(n_1413),
.B(n_1581),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1506),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1400),
.A2(n_1485),
.B(n_1431),
.Y(n_1694)
);

NOR2xp67_ASAP7_75t_L g1695 ( 
.A(n_1422),
.B(n_1039),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_SL g1696 ( 
.A(n_1418),
.B(n_1040),
.Y(n_1696)
);

INVx8_ASAP7_75t_L g1697 ( 
.A(n_1403),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1459),
.B(n_1120),
.Y(n_1699)
);

OA21x2_ASAP7_75t_L g1700 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1316),
.Y(n_1700)
);

NOR2xp67_ASAP7_75t_L g1701 ( 
.A(n_1422),
.B(n_1039),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1416),
.A2(n_1180),
.B1(n_735),
.B2(n_1317),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1438),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_SL g1704 ( 
.A1(n_1580),
.A2(n_1466),
.B(n_1399),
.Y(n_1704)
);

AO21x2_ASAP7_75t_L g1705 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1429),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_SL g1706 ( 
.A(n_1514),
.B(n_1039),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1430),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1404),
.A2(n_1180),
.B1(n_1150),
.B2(n_1530),
.Y(n_1709)
);

INVx4_ASAP7_75t_L g1710 ( 
.A(n_1536),
.Y(n_1710)
);

NOR2xp67_ASAP7_75t_SL g1711 ( 
.A(n_1535),
.B(n_1191),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1404),
.A2(n_1180),
.B1(n_1150),
.B2(n_1530),
.Y(n_1712)
);

INVxp67_ASAP7_75t_L g1713 ( 
.A(n_1483),
.Y(n_1713)
);

OAI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1404),
.A2(n_1180),
.B1(n_1150),
.B2(n_1530),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1316),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1536),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1440),
.B(n_1452),
.Y(n_1719)
);

CKINVDCx6p67_ASAP7_75t_R g1720 ( 
.A(n_1403),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1416),
.A2(n_1180),
.B1(n_735),
.B2(n_1317),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1404),
.A2(n_1150),
.B(n_1180),
.C(n_964),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1409),
.B(n_1120),
.Y(n_1724)
);

OR2x6_ASAP7_75t_L g1725 ( 
.A(n_1535),
.B(n_1466),
.Y(n_1725)
);

AOI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1439),
.A2(n_1402),
.B(n_1412),
.Y(n_1726)
);

AO31x2_ASAP7_75t_L g1727 ( 
.A1(n_1541),
.A2(n_1251),
.A3(n_1487),
.B(n_1546),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1728)
);

OAI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1580),
.A2(n_1180),
.B1(n_1352),
.B2(n_1546),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1438),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1316),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1536),
.Y(n_1732)
);

OAI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1580),
.A2(n_1180),
.B1(n_1352),
.B2(n_1546),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1416),
.A2(n_1180),
.B1(n_735),
.B2(n_1317),
.Y(n_1735)
);

AOI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1439),
.A2(n_1402),
.B(n_1412),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1409),
.B(n_1120),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1500),
.Y(n_1738)
);

BUFx8_ASAP7_75t_SL g1739 ( 
.A(n_1514),
.Y(n_1739)
);

OAI22x1_ASAP7_75t_L g1740 ( 
.A1(n_1455),
.A2(n_1150),
.B1(n_1392),
.B2(n_1180),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1500),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1536),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1409),
.B(n_1180),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1535),
.B(n_1466),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1524),
.B(n_1490),
.Y(n_1745)
);

BUFx4f_ASAP7_75t_L g1746 ( 
.A(n_1414),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1404),
.A2(n_488),
.B1(n_516),
.B2(n_498),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1500),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1416),
.A2(n_1180),
.B1(n_735),
.B2(n_1317),
.Y(n_1749)
);

NOR4xp25_ASAP7_75t_L g1750 ( 
.A(n_1404),
.B(n_1150),
.C(n_1180),
.D(n_1274),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1500),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1316),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1404),
.A2(n_1180),
.B(n_1150),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1438),
.Y(n_1754)
);

OAI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1459),
.B(n_1120),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1500),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1409),
.B(n_1120),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1493),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1544),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1409),
.B(n_1180),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1500),
.Y(n_1762)
);

OAI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1530),
.A2(n_1180),
.B1(n_1150),
.B2(n_964),
.C(n_731),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1404),
.B(n_1180),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1404),
.A2(n_1180),
.B1(n_1150),
.B2(n_1530),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1446),
.Y(n_1766)
);

OA21x2_ASAP7_75t_L g1767 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1316),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1446),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_SL g1773 ( 
.A1(n_1580),
.A2(n_1466),
.B(n_1399),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1500),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1541),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1500),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1580),
.A2(n_1180),
.B1(n_1352),
.B2(n_1546),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1500),
.Y(n_1778)
);

AO21x2_ASAP7_75t_L g1779 ( 
.A1(n_1485),
.A2(n_1431),
.B(n_1429),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1408),
.A2(n_1439),
.B(n_1230),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1404),
.B(n_1180),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1594),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1601),
.B(n_1699),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1595),
.A2(n_1607),
.B1(n_1763),
.B2(n_1592),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1593),
.B(n_1612),
.Y(n_1785)
);

O2A1O1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1729),
.A2(n_1777),
.B(n_1733),
.C(n_1764),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1729),
.A2(n_1777),
.B(n_1733),
.Y(n_1787)
);

AOI21x1_ASAP7_75t_SL g1788 ( 
.A1(n_1683),
.A2(n_1737),
.B(n_1724),
.Y(n_1788)
);

O2A1O1Ixp5_ASAP7_75t_L g1789 ( 
.A1(n_1614),
.A2(n_1616),
.B(n_1634),
.C(n_1690),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1593),
.B(n_1612),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1756),
.B(n_1618),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1764),
.A2(n_1781),
.B1(n_1750),
.B2(n_1595),
.C(n_1723),
.Y(n_1792)
);

O2A1O1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1781),
.A2(n_1761),
.B(n_1743),
.C(n_1753),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1739),
.Y(n_1794)
);

BUFx8_ASAP7_75t_SL g1795 ( 
.A(n_1759),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1599),
.Y(n_1796)
);

OA21x2_ASAP7_75t_L g1797 ( 
.A1(n_1689),
.A2(n_1692),
.B(n_1663),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1746),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1738),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1702),
.A2(n_1735),
.B(n_1722),
.Y(n_1800)
);

AND2x2_ASAP7_75t_SL g1801 ( 
.A(n_1585),
.B(n_1582),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1719),
.B(n_1740),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1585),
.A2(n_1616),
.B(n_1749),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1741),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1748),
.Y(n_1805)
);

A2O1A1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1685),
.A2(n_1629),
.B(n_1626),
.C(n_1709),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1610),
.Y(n_1807)
);

OR2x6_ASAP7_75t_L g1808 ( 
.A(n_1605),
.B(n_1725),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1746),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1696),
.A2(n_1664),
.B(n_1743),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1718),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1719),
.B(n_1633),
.Y(n_1812)
);

OA21x2_ASAP7_75t_L g1813 ( 
.A1(n_1689),
.A2(n_1692),
.B(n_1663),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1617),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1739),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1649),
.B(n_1583),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1583),
.B(n_1670),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1670),
.B(n_1679),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1664),
.A2(n_1761),
.B(n_1758),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1644),
.B(n_1602),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1745),
.B(n_1650),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1710),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1647),
.A2(n_1603),
.B(n_1584),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1584),
.B(n_1603),
.Y(n_1824)
);

OA22x2_ASAP7_75t_L g1825 ( 
.A1(n_1635),
.A2(n_1662),
.B1(n_1747),
.B2(n_1704),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1708),
.B(n_1643),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1670),
.B(n_1677),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1709),
.B(n_1712),
.Y(n_1828)
);

OAI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1712),
.A2(n_1765),
.B(n_1715),
.C(n_1611),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1715),
.A2(n_1765),
.B1(n_1626),
.B2(n_1586),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1708),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1751),
.B(n_1757),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1762),
.B(n_1774),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1605),
.A2(n_1725),
.B(n_1744),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1776),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1664),
.A2(n_1685),
.B(n_1605),
.Y(n_1836)
);

AOI21x1_ASAP7_75t_SL g1837 ( 
.A1(n_1676),
.A2(n_1711),
.B(n_1687),
.Y(n_1837)
);

CKINVDCx6p67_ASAP7_75t_R g1838 ( 
.A(n_1759),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1778),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1589),
.A2(n_1773),
.B(n_1632),
.C(n_1713),
.Y(n_1840)
);

OA21x2_ASAP7_75t_L g1841 ( 
.A1(n_1682),
.A2(n_1684),
.B(n_1658),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1659),
.B(n_1665),
.Y(n_1842)
);

AOI31xp33_ASAP7_75t_L g1843 ( 
.A1(n_1638),
.A2(n_1598),
.A3(n_1632),
.B(n_1646),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1628),
.B(n_1631),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1631),
.B(n_1766),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1628),
.B(n_1771),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1688),
.B(n_1681),
.Y(n_1847)
);

O2A1O1Ixp5_ASAP7_75t_L g1848 ( 
.A1(n_1691),
.A2(n_1726),
.B(n_1736),
.C(n_1606),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1667),
.B(n_1582),
.Y(n_1849)
);

AOI211xp5_ASAP7_75t_L g1850 ( 
.A1(n_1695),
.A2(n_1701),
.B(n_1668),
.C(n_1693),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1725),
.A2(n_1744),
.B(n_1582),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1686),
.A2(n_1645),
.B(n_1653),
.C(n_1624),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1628),
.B(n_1653),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1744),
.A2(n_1675),
.B(n_1655),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1640),
.A2(n_1615),
.B1(n_1645),
.B2(n_1720),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1600),
.B(n_1621),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1628),
.B(n_1667),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1710),
.A2(n_1703),
.B1(n_1730),
.B2(n_1623),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1710),
.A2(n_1703),
.B1(n_1730),
.B2(n_1623),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1652),
.A2(n_1754),
.B1(n_1637),
.B2(n_1697),
.Y(n_1860)
);

AOI21x1_ASAP7_75t_SL g1861 ( 
.A1(n_1604),
.A2(n_1620),
.B(n_1779),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1628),
.B(n_1667),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1667),
.B(n_1705),
.Y(n_1863)
);

AOI21x1_ASAP7_75t_SL g1864 ( 
.A1(n_1604),
.A2(n_1620),
.B(n_1705),
.Y(n_1864)
);

AND2x2_ASAP7_75t_SL g1865 ( 
.A(n_1625),
.B(n_1700),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1622),
.B(n_1660),
.Y(n_1866)
);

OA22x2_ASAP7_75t_L g1867 ( 
.A1(n_1681),
.A2(n_1673),
.B1(n_1742),
.B2(n_1732),
.Y(n_1867)
);

A2O1A1Ixp33_ASAP7_75t_L g1868 ( 
.A1(n_1624),
.A2(n_1672),
.B(n_1678),
.C(n_1641),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1681),
.B(n_1671),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_SL g1870 ( 
.A1(n_1655),
.A2(n_1678),
.B(n_1642),
.Y(n_1870)
);

INVx8_ASAP7_75t_L g1871 ( 
.A(n_1637),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1779),
.B(n_1642),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1700),
.B(n_1752),
.Y(n_1873)
);

A2O1A1Ixp33_ASAP7_75t_L g1874 ( 
.A1(n_1672),
.A2(n_1678),
.B(n_1641),
.C(n_1609),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1775),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1671),
.B(n_1674),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1694),
.A2(n_1697),
.B1(n_1691),
.B2(n_1656),
.C(n_1654),
.Y(n_1877)
);

O2A1O1Ixp5_ASAP7_75t_L g1878 ( 
.A1(n_1691),
.A2(n_1588),
.B(n_1656),
.C(n_1654),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1609),
.A2(n_1651),
.B(n_1608),
.C(n_1680),
.Y(n_1879)
);

INVx4_ASAP7_75t_L g1880 ( 
.A(n_1622),
.Y(n_1880)
);

INVx1_ASAP7_75t_SL g1881 ( 
.A(n_1660),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1657),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1642),
.A2(n_1625),
.B(n_1590),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1700),
.A2(n_1752),
.B(n_1731),
.Y(n_1884)
);

INVxp33_ASAP7_75t_SL g1885 ( 
.A(n_1706),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1694),
.A2(n_1716),
.B(n_1767),
.C(n_1669),
.Y(n_1886)
);

NOR2x1_ASAP7_75t_SL g1887 ( 
.A(n_1661),
.B(n_1666),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1760),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1760),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1590),
.Y(n_1890)
);

OA21x2_ASAP7_75t_L g1891 ( 
.A1(n_1597),
.A2(n_1707),
.B(n_1772),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1767),
.A2(n_1625),
.B1(n_1590),
.B2(n_1639),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1767),
.Y(n_1893)
);

NOR2xp67_ASAP7_75t_L g1894 ( 
.A(n_1627),
.B(n_1630),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1619),
.B(n_1727),
.Y(n_1895)
);

AOI21x1_ASAP7_75t_SL g1896 ( 
.A1(n_1619),
.A2(n_1727),
.B(n_1648),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1619),
.B(n_1727),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1619),
.B(n_1727),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1648),
.B(n_1587),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1591),
.B(n_1680),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1591),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1639),
.A2(n_1613),
.B(n_1630),
.Y(n_1902)
);

OAI31xp33_ASAP7_75t_L g1903 ( 
.A1(n_1627),
.A2(n_1648),
.A3(n_1639),
.B(n_1636),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1698),
.B(n_1734),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1707),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1714),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_SL g1907 ( 
.A1(n_1714),
.A2(n_1755),
.B(n_1717),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1721),
.Y(n_1908)
);

BUFx2_ASAP7_75t_L g1909 ( 
.A(n_1721),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1780),
.B(n_1768),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1728),
.B(n_1734),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1728),
.B(n_1755),
.Y(n_1912)
);

AOI21x1_ASAP7_75t_SL g1913 ( 
.A1(n_1769),
.A2(n_1770),
.B(n_1772),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1596),
.A2(n_1352),
.B(n_1580),
.Y(n_1914)
);

O2A1O1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1592),
.A2(n_1150),
.B(n_1180),
.C(n_1763),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1766),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1601),
.B(n_1699),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1595),
.A2(n_1180),
.B1(n_1607),
.B2(n_1763),
.Y(n_1918)
);

O2A1O1Ixp33_ASAP7_75t_L g1919 ( 
.A1(n_1592),
.A2(n_1150),
.B(n_1180),
.C(n_1763),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1729),
.A2(n_1150),
.B(n_735),
.Y(n_1920)
);

INVx2_ASAP7_75t_SL g1921 ( 
.A(n_1637),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1622),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1595),
.A2(n_1180),
.B1(n_1607),
.B2(n_1763),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1637),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1594),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1583),
.B(n_1719),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1702),
.A2(n_1352),
.B(n_1580),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1729),
.A2(n_1150),
.B(n_735),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1601),
.B(n_1699),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1584),
.Y(n_1930)
);

BUFx3_ASAP7_75t_L g1931 ( 
.A(n_1718),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1702),
.A2(n_1352),
.B(n_1580),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1601),
.B(n_1699),
.Y(n_1933)
);

O2A1O1Ixp5_ASAP7_75t_L g1934 ( 
.A1(n_1729),
.A2(n_1733),
.B(n_1777),
.C(n_1614),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1595),
.A2(n_1180),
.B1(n_1607),
.B2(n_1763),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1584),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1593),
.B(n_1612),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1729),
.A2(n_1150),
.B(n_735),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1593),
.B(n_1612),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_SL g1940 ( 
.A1(n_1702),
.A2(n_1352),
.B(n_1580),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1622),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1831),
.Y(n_1942)
);

AO21x1_ASAP7_75t_L g1943 ( 
.A1(n_1787),
.A2(n_1784),
.B(n_1786),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1930),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1802),
.B(n_1812),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1857),
.B(n_1862),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1863),
.B(n_1849),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1848),
.A2(n_1789),
.B(n_1884),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1865),
.B(n_1801),
.Y(n_1949)
);

BUFx2_ASAP7_75t_L g1950 ( 
.A(n_1936),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1936),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1865),
.B(n_1801),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1872),
.B(n_1824),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1844),
.B(n_1808),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1915),
.A2(n_1919),
.B(n_1934),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1887),
.Y(n_1956)
);

AO21x2_ASAP7_75t_L g1957 ( 
.A1(n_1874),
.A2(n_1879),
.B(n_1868),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1797),
.Y(n_1958)
);

AO21x2_ASAP7_75t_L g1959 ( 
.A1(n_1874),
.A2(n_1879),
.B(n_1868),
.Y(n_1959)
);

BUFx2_ASAP7_75t_L g1960 ( 
.A(n_1906),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1813),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1808),
.B(n_1900),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1826),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1808),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_SL g1965 ( 
.A1(n_1918),
.A2(n_1923),
.B1(n_1935),
.B2(n_1825),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1796),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1785),
.B(n_1790),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1900),
.B(n_1894),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1821),
.Y(n_1969)
);

OAI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1915),
.A2(n_1919),
.B(n_1934),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1807),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1926),
.B(n_1814),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1890),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1783),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1871),
.Y(n_1975)
);

OAI21x1_ASAP7_75t_L g1976 ( 
.A1(n_1913),
.A2(n_1848),
.B(n_1902),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1841),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1895),
.B(n_1897),
.Y(n_1978)
);

OR2x6_ASAP7_75t_L g1979 ( 
.A(n_1851),
.B(n_1836),
.Y(n_1979)
);

INVxp33_ASAP7_75t_L g1980 ( 
.A(n_1795),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1786),
.A2(n_1806),
.B(n_1843),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1937),
.B(n_1939),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1841),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1901),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1841),
.Y(n_1985)
);

OR2x6_ASAP7_75t_L g1986 ( 
.A(n_1834),
.B(n_1870),
.Y(n_1986)
);

AO21x2_ASAP7_75t_L g1987 ( 
.A1(n_1803),
.A2(n_1907),
.B(n_1852),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1901),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1875),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1926),
.B(n_1846),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1899),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1845),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1898),
.B(n_1893),
.Y(n_1993)
);

AO21x2_ASAP7_75t_L g1994 ( 
.A1(n_1852),
.A2(n_1892),
.B(n_1883),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1817),
.B(n_1816),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1782),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1799),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1867),
.Y(n_1998)
);

BUFx2_ASAP7_75t_L g1999 ( 
.A(n_1867),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1823),
.B(n_1853),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1910),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1804),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1905),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1818),
.B(n_1827),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1891),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1911),
.B(n_1904),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1805),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1835),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1839),
.B(n_1925),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1878),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1878),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1873),
.B(n_1909),
.Y(n_2012)
);

OAI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1825),
.A2(n_1806),
.B1(n_1792),
.B2(n_1830),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1789),
.B(n_1832),
.Y(n_2014)
);

INVx4_ASAP7_75t_L g2015 ( 
.A(n_1871),
.Y(n_2015)
);

NAND3xp33_ASAP7_75t_L g2016 ( 
.A(n_1829),
.B(n_1793),
.C(n_1840),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1916),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1833),
.B(n_1842),
.Y(n_2018)
);

AO21x2_ASAP7_75t_L g2019 ( 
.A1(n_1920),
.A2(n_1928),
.B(n_1938),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1791),
.B(n_1877),
.Y(n_2020)
);

CKINVDCx16_ASAP7_75t_R g2021 ( 
.A(n_1922),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1912),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1908),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1888),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1889),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1856),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1886),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1869),
.B(n_1856),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1886),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_L g2030 ( 
.A(n_1793),
.B(n_1840),
.C(n_1850),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1914),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1917),
.B(n_1933),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_2013),
.A2(n_1855),
.B1(n_1940),
.B2(n_1932),
.C(n_1927),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1967),
.B(n_1885),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1949),
.B(n_1929),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1953),
.B(n_1903),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1949),
.B(n_1876),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1963),
.B(n_1820),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1953),
.B(n_1800),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1988),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1966),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1971),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1971),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1942),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1952),
.B(n_1847),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_2001),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2000),
.B(n_1819),
.Y(n_2047)
);

OAI211xp5_ASAP7_75t_SL g2048 ( 
.A1(n_1981),
.A2(n_1828),
.B(n_1810),
.C(n_1881),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_2003),
.Y(n_2049)
);

BUFx12f_ASAP7_75t_L g2050 ( 
.A(n_1975),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2000),
.B(n_1860),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1981),
.A2(n_1970),
.B(n_1955),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1942),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1947),
.B(n_1861),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_2003),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1947),
.B(n_1864),
.Y(n_2056)
);

INVxp67_ASAP7_75t_L g2057 ( 
.A(n_2017),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1950),
.Y(n_2058)
);

INVxp67_ASAP7_75t_SL g2059 ( 
.A(n_1969),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1965),
.A2(n_1880),
.B1(n_1922),
.B2(n_1941),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_1968),
.Y(n_2061)
);

OAI211xp5_ASAP7_75t_SL g2062 ( 
.A1(n_2016),
.A2(n_1854),
.B(n_1921),
.C(n_1924),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1973),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1973),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_1946),
.B(n_1864),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2005),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1945),
.B(n_1941),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2005),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2022),
.B(n_1991),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_1943),
.A2(n_1880),
.B1(n_1838),
.B2(n_1941),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_2006),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1991),
.B(n_1922),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_2012),
.B(n_1896),
.Y(n_2073)
);

INVx4_ASAP7_75t_L g2074 ( 
.A(n_1979),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2014),
.B(n_1866),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1992),
.B(n_1858),
.Y(n_2076)
);

INVxp67_ASAP7_75t_SL g2077 ( 
.A(n_1993),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1974),
.Y(n_2078)
);

INVxp67_ASAP7_75t_L g2079 ( 
.A(n_2024),
.Y(n_2079)
);

INVx4_ASAP7_75t_L g2080 ( 
.A(n_1979),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2014),
.B(n_1866),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_1976),
.A2(n_1837),
.B(n_1788),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_2006),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1944),
.Y(n_2084)
);

OAI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2030),
.A2(n_1822),
.B1(n_1859),
.B2(n_1931),
.C(n_1811),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_1978),
.B(n_1871),
.Y(n_2086)
);

OAI332xp33_ASAP7_75t_L g2087 ( 
.A1(n_2060),
.A2(n_1982),
.A3(n_2021),
.B1(n_1943),
.B2(n_2029),
.B3(n_2027),
.C1(n_2031),
.C2(n_2011),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2075),
.B(n_1994),
.Y(n_2088)
);

A2O1A1Ixp33_ASAP7_75t_L g2089 ( 
.A1(n_2052),
.A2(n_2031),
.B(n_1999),
.C(n_1998),
.Y(n_2089)
);

OAI211xp5_ASAP7_75t_L g2090 ( 
.A1(n_2033),
.A2(n_1998),
.B(n_1999),
.C(n_2020),
.Y(n_2090)
);

BUFx2_ASAP7_75t_L g2091 ( 
.A(n_2055),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2075),
.B(n_1994),
.Y(n_2092)
);

OAI221xp5_ASAP7_75t_L g2093 ( 
.A1(n_2070),
.A2(n_2047),
.B1(n_2048),
.B2(n_2062),
.C(n_2085),
.Y(n_2093)
);

OAI221xp5_ASAP7_75t_L g2094 ( 
.A1(n_2051),
.A2(n_1979),
.B1(n_1986),
.B2(n_1960),
.C(n_1964),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2049),
.Y(n_2095)
);

OAI33xp33_ASAP7_75t_L g2096 ( 
.A1(n_2065),
.A2(n_1978),
.A3(n_2029),
.B1(n_2027),
.B2(n_1951),
.B3(n_2011),
.Y(n_2096)
);

AO21x2_ASAP7_75t_L g2097 ( 
.A1(n_2066),
.A2(n_2010),
.B(n_1983),
.Y(n_2097)
);

OAI21xp5_ASAP7_75t_SL g2098 ( 
.A1(n_2081),
.A2(n_1980),
.B(n_2020),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_R g2099 ( 
.A(n_2050),
.B(n_1794),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2041),
.Y(n_2100)
);

BUFx2_ASAP7_75t_L g2101 ( 
.A(n_2055),
.Y(n_2101)
);

AO21x2_ASAP7_75t_L g2102 ( 
.A1(n_2066),
.A2(n_2010),
.B(n_1977),
.Y(n_2102)
);

NAND3xp33_ASAP7_75t_L g2103 ( 
.A(n_2039),
.B(n_1956),
.C(n_1954),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_2081),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2041),
.Y(n_2105)
);

NAND2x1_ASAP7_75t_L g2106 ( 
.A(n_2061),
.B(n_1979),
.Y(n_2106)
);

NAND3xp33_ASAP7_75t_L g2107 ( 
.A(n_2039),
.B(n_2065),
.C(n_2036),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_2049),
.Y(n_2108)
);

OAI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_2074),
.A2(n_1986),
.B1(n_1964),
.B2(n_2021),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2042),
.Y(n_2110)
);

OAI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2038),
.A2(n_1986),
.B1(n_1960),
.B2(n_1964),
.C(n_1956),
.Y(n_2111)
);

OAI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_2086),
.A2(n_1986),
.B1(n_1954),
.B2(n_2015),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_2044),
.Y(n_2113)
);

INVxp67_ASAP7_75t_L g2114 ( 
.A(n_2059),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2061),
.B(n_1994),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_2040),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2043),
.Y(n_2117)
);

AOI211xp5_ASAP7_75t_SL g2118 ( 
.A1(n_2036),
.A2(n_1962),
.B(n_1954),
.C(n_1984),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2083),
.B(n_1990),
.Y(n_2119)
);

NAND4xp25_ASAP7_75t_SL g2120 ( 
.A(n_2067),
.B(n_2032),
.C(n_1972),
.D(n_1795),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_2083),
.Y(n_2121)
);

NOR4xp25_ASAP7_75t_SL g2122 ( 
.A(n_2077),
.B(n_1815),
.C(n_2026),
.D(n_1882),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_2057),
.B(n_2032),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2034),
.A2(n_2019),
.B1(n_1987),
.B2(n_1954),
.Y(n_2124)
);

NAND2xp33_ASAP7_75t_R g2125 ( 
.A(n_2054),
.B(n_1986),
.Y(n_2125)
);

OAI211xp5_ASAP7_75t_L g2126 ( 
.A1(n_2076),
.A2(n_1948),
.B(n_2025),
.C(n_2007),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_2078),
.A2(n_2019),
.B1(n_1987),
.B2(n_1972),
.Y(n_2127)
);

AOI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_2074),
.A2(n_2080),
.B1(n_2079),
.B2(n_2072),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_2074),
.A2(n_2004),
.B1(n_2008),
.B2(n_1996),
.Y(n_2129)
);

INVxp67_ASAP7_75t_SL g2130 ( 
.A(n_2053),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2083),
.B(n_1962),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_SL g2132 ( 
.A1(n_2074),
.A2(n_1962),
.B1(n_1957),
.B2(n_1959),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2037),
.B(n_2028),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2071),
.B(n_2045),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_2058),
.B(n_2023),
.Y(n_2135)
);

AOI221xp5_ASAP7_75t_L g2136 ( 
.A1(n_2035),
.A2(n_2008),
.B1(n_1996),
.B2(n_1997),
.C(n_2002),
.Y(n_2136)
);

OAI221xp5_ASAP7_75t_L g2137 ( 
.A1(n_2080),
.A2(n_1975),
.B1(n_2026),
.B2(n_2015),
.C(n_2002),
.Y(n_2137)
);

BUFx3_ASAP7_75t_L g2138 ( 
.A(n_2050),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2037),
.B(n_2028),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_2080),
.A2(n_2004),
.B1(n_1997),
.B2(n_2007),
.Y(n_2140)
);

AOI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2035),
.A2(n_2018),
.B1(n_2009),
.B2(n_1995),
.C(n_1989),
.Y(n_2141)
);

OAI211xp5_ASAP7_75t_SL g2142 ( 
.A1(n_2056),
.A2(n_2073),
.B(n_2086),
.C(n_2084),
.Y(n_2142)
);

AO21x2_ASAP7_75t_L g2143 ( 
.A1(n_2068),
.A2(n_1983),
.B(n_1985),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2107),
.B(n_2046),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_2115),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_2116),
.Y(n_2146)
);

AO21x1_ASAP7_75t_L g2147 ( 
.A1(n_2098),
.A2(n_2063),
.B(n_2064),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_2097),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_2143),
.Y(n_2149)
);

INVx4_ASAP7_75t_L g2150 ( 
.A(n_2138),
.Y(n_2150)
);

INVx4_ASAP7_75t_SL g2151 ( 
.A(n_2116),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_2115),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2088),
.B(n_2069),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_2091),
.Y(n_2154)
);

HB1xp67_ASAP7_75t_L g2155 ( 
.A(n_2102),
.Y(n_2155)
);

BUFx2_ASAP7_75t_L g2156 ( 
.A(n_2121),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2100),
.Y(n_2157)
);

INVx4_ASAP7_75t_L g2158 ( 
.A(n_2138),
.Y(n_2158)
);

INVx4_ASAP7_75t_SL g2159 ( 
.A(n_2116),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2105),
.Y(n_2160)
);

OA21x2_ASAP7_75t_L g2161 ( 
.A1(n_2126),
.A2(n_1961),
.B(n_1958),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_2110),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_2101),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_2106),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_2099),
.Y(n_2165)
);

INVx4_ASAP7_75t_L g2166 ( 
.A(n_2116),
.Y(n_2166)
);

OR2x6_ASAP7_75t_L g2167 ( 
.A(n_2089),
.B(n_2080),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_SL g2168 ( 
.A1(n_2094),
.A2(n_2015),
.B(n_1962),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2117),
.Y(n_2169)
);

AOI21xp5_ASAP7_75t_L g2170 ( 
.A1(n_2087),
.A2(n_1959),
.B(n_1957),
.Y(n_2170)
);

INVxp67_ASAP7_75t_SL g2171 ( 
.A(n_2095),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2121),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_2137),
.Y(n_2173)
);

NOR2x1p5_ASAP7_75t_L g2174 ( 
.A(n_2103),
.B(n_2015),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2092),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2162),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2149),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2164),
.B(n_2092),
.Y(n_2178)
);

INVx1_ASAP7_75t_SL g2179 ( 
.A(n_2165),
.Y(n_2179)
);

AND4x1_ASAP7_75t_L g2180 ( 
.A(n_2170),
.B(n_2118),
.C(n_2096),
.D(n_2124),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2170),
.A2(n_2090),
.B1(n_2125),
.B2(n_2124),
.Y(n_2181)
);

NAND3xp33_ASAP7_75t_SL g2182 ( 
.A(n_2147),
.B(n_2122),
.C(n_2093),
.Y(n_2182)
);

INVx1_ASAP7_75t_SL g2183 ( 
.A(n_2165),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2162),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2149),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2164),
.B(n_2131),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2164),
.B(n_2131),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2144),
.B(n_2135),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2149),
.Y(n_2189)
);

INVxp67_ASAP7_75t_SL g2190 ( 
.A(n_2147),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_2151),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2164),
.B(n_2119),
.Y(n_2192)
);

INVx1_ASAP7_75t_SL g2193 ( 
.A(n_2154),
.Y(n_2193)
);

INVx3_ASAP7_75t_SL g2194 ( 
.A(n_2150),
.Y(n_2194)
);

OAI21xp5_ASAP7_75t_SL g2195 ( 
.A1(n_2154),
.A2(n_2132),
.B(n_2127),
.Y(n_2195)
);

BUFx3_ASAP7_75t_L g2196 ( 
.A(n_2150),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2173),
.B(n_2104),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2174),
.B(n_2119),
.Y(n_2198)
);

INVx4_ASAP7_75t_L g2199 ( 
.A(n_2150),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2157),
.Y(n_2200)
);

OAI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_2168),
.A2(n_2127),
.B(n_2111),
.Y(n_2201)
);

OAI22xp5_ASAP7_75t_L g2202 ( 
.A1(n_2173),
.A2(n_2128),
.B1(n_2129),
.B2(n_2140),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2174),
.B(n_2134),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2157),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2149),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2157),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2145),
.B(n_2134),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2173),
.B(n_2141),
.Y(n_2208)
);

OR2x6_ASAP7_75t_L g2209 ( 
.A(n_2167),
.B(n_2082),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_2150),
.B(n_2120),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2160),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2145),
.B(n_2108),
.Y(n_2212)
);

OR2x6_ASAP7_75t_L g2213 ( 
.A(n_2167),
.B(n_2112),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2145),
.B(n_2133),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2160),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_2150),
.B(n_2099),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_2151),
.B(n_2159),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2152),
.B(n_2139),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2173),
.B(n_2123),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2160),
.Y(n_2220)
);

AOI33xp33_ASAP7_75t_L g2221 ( 
.A1(n_2175),
.A2(n_2140),
.A3(n_2129),
.B1(n_2128),
.B2(n_2136),
.B3(n_2109),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_R g2222 ( 
.A(n_2158),
.B(n_2125),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2158),
.B(n_2123),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2169),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2151),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_2158),
.B(n_2114),
.Y(n_2226)
);

AOI222xp33_ASAP7_75t_L g2227 ( 
.A1(n_2158),
.A2(n_2142),
.B1(n_2130),
.B2(n_2067),
.C1(n_2113),
.C2(n_2072),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2217),
.B(n_2151),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2200),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2193),
.B(n_2219),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2179),
.B(n_2158),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2183),
.B(n_2216),
.Y(n_2232)
);

NAND3xp33_ASAP7_75t_L g2233 ( 
.A(n_2180),
.B(n_2167),
.C(n_2161),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2217),
.B(n_2151),
.Y(n_2234)
);

NAND2x1p5_ASAP7_75t_L g2235 ( 
.A(n_2180),
.B(n_2166),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2208),
.B(n_2163),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2217),
.B(n_2151),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2221),
.B(n_2163),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2188),
.B(n_2144),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2200),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_R g2241 ( 
.A(n_2182),
.B(n_1798),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2204),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2223),
.B(n_2147),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2204),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2206),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2217),
.B(n_2151),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2188),
.B(n_2144),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2177),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2203),
.B(n_2159),
.Y(n_2249)
);

NOR2x1_ASAP7_75t_L g2250 ( 
.A(n_2199),
.B(n_2166),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2203),
.B(n_2159),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2206),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2197),
.B(n_2171),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2177),
.Y(n_2254)
);

INVx1_ASAP7_75t_SL g2255 ( 
.A(n_2194),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2211),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2211),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2186),
.B(n_2159),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2215),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2186),
.B(n_2187),
.Y(n_2260)
);

OAI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2181),
.A2(n_2167),
.B(n_2171),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2187),
.B(n_2159),
.Y(n_2262)
);

OR2x2_ASAP7_75t_L g2263 ( 
.A(n_2176),
.B(n_2175),
.Y(n_2263)
);

NAND2x1_ASAP7_75t_L g2264 ( 
.A(n_2191),
.B(n_2152),
.Y(n_2264)
);

AOI22xp33_ASAP7_75t_L g2265 ( 
.A1(n_2201),
.A2(n_2167),
.B1(n_1957),
.B2(n_1959),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2215),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2192),
.B(n_2159),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2195),
.B(n_2153),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2176),
.B(n_2175),
.Y(n_2269)
);

NOR3xp33_ASAP7_75t_L g2270 ( 
.A(n_2232),
.B(n_2199),
.C(n_2190),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2229),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2235),
.B(n_2222),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2229),
.Y(n_2273)
);

CKINVDCx16_ASAP7_75t_R g2274 ( 
.A(n_2241),
.Y(n_2274)
);

INVx1_ASAP7_75t_SL g2275 ( 
.A(n_2258),
.Y(n_2275)
);

AOI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2238),
.A2(n_2202),
.B1(n_2210),
.B2(n_2226),
.Y(n_2276)
);

HB1xp67_ASAP7_75t_L g2277 ( 
.A(n_2264),
.Y(n_2277)
);

AO21x2_ASAP7_75t_L g2278 ( 
.A1(n_2233),
.A2(n_2261),
.B(n_2243),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2258),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2264),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2240),
.Y(n_2281)
);

INVx1_ASAP7_75t_SL g2282 ( 
.A(n_2262),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2265),
.A2(n_2167),
.B1(n_2213),
.B2(n_2194),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2240),
.Y(n_2284)
);

BUFx3_ASAP7_75t_L g2285 ( 
.A(n_2235),
.Y(n_2285)
);

INVx1_ASAP7_75t_SL g2286 ( 
.A(n_2262),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2260),
.B(n_2191),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2230),
.B(n_2199),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_2267),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2242),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2242),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2260),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2244),
.Y(n_2293)
);

HB1xp67_ASAP7_75t_L g2294 ( 
.A(n_2239),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2267),
.B(n_2225),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2239),
.B(n_2184),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2235),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_2247),
.B(n_2184),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2255),
.B(n_2214),
.Y(n_2299)
);

AOI21xp5_ASAP7_75t_L g2300 ( 
.A1(n_2278),
.A2(n_2236),
.B(n_2268),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_2292),
.B(n_2253),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2294),
.Y(n_2302)
);

AOI222xp33_ASAP7_75t_L g2303 ( 
.A1(n_2272),
.A2(n_2231),
.B1(n_2249),
.B2(n_2251),
.C1(n_2228),
.C2(n_2237),
.Y(n_2303)
);

OAI221xp5_ASAP7_75t_L g2304 ( 
.A1(n_2276),
.A2(n_2213),
.B1(n_2250),
.B2(n_2194),
.C(n_2225),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2292),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2292),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2280),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2296),
.Y(n_2308)
);

OAI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2276),
.A2(n_2213),
.B1(n_2209),
.B2(n_2251),
.C(n_2249),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2296),
.Y(n_2310)
);

NAND3xp33_ASAP7_75t_L g2311 ( 
.A(n_2270),
.B(n_2247),
.C(n_2196),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2274),
.B(n_2227),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2295),
.B(n_2228),
.Y(n_2313)
);

AOI21xp33_ASAP7_75t_SL g2314 ( 
.A1(n_2274),
.A2(n_2278),
.B(n_2288),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2275),
.B(n_2279),
.Y(n_2315)
);

AOI32xp33_ASAP7_75t_L g2316 ( 
.A1(n_2282),
.A2(n_2237),
.A3(n_2234),
.B1(n_2246),
.B2(n_2178),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2278),
.A2(n_2246),
.B(n_2234),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2286),
.B(n_2214),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2298),
.Y(n_2319)
);

AOI222xp33_ASAP7_75t_L g2320 ( 
.A1(n_2283),
.A2(n_2212),
.B1(n_2152),
.B2(n_2178),
.C1(n_2259),
.C2(n_2257),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2298),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2285),
.A2(n_2213),
.B1(n_2167),
.B2(n_2209),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2313),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2305),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2302),
.B(n_2289),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2300),
.B(n_2287),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_2314),
.B(n_2285),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2300),
.B(n_2287),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2318),
.B(n_2299),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2306),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2308),
.B(n_2295),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2310),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2319),
.Y(n_2333)
);

OA21x2_ASAP7_75t_L g2334 ( 
.A1(n_2312),
.A2(n_2297),
.B(n_2280),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2321),
.B(n_2285),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2307),
.Y(n_2336)
);

INVx1_ASAP7_75t_SL g2337 ( 
.A(n_2315),
.Y(n_2337)
);

AOI221xp5_ASAP7_75t_SL g2338 ( 
.A1(n_2326),
.A2(n_2304),
.B1(n_2317),
.B2(n_2309),
.C(n_2322),
.Y(n_2338)
);

AOI211xp5_ASAP7_75t_L g2339 ( 
.A1(n_2328),
.A2(n_2311),
.B(n_2317),
.C(n_2301),
.Y(n_2339)
);

OAI21xp5_ASAP7_75t_SL g2340 ( 
.A1(n_2337),
.A2(n_2303),
.B(n_2316),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2323),
.B(n_2297),
.Y(n_2341)
);

O2A1O1Ixp33_ASAP7_75t_L g2342 ( 
.A1(n_2327),
.A2(n_2297),
.B(n_2277),
.C(n_2320),
.Y(n_2342)
);

OAI211xp5_ASAP7_75t_L g2343 ( 
.A1(n_2334),
.A2(n_2327),
.B(n_2335),
.C(n_2331),
.Y(n_2343)
);

AOI222xp33_ASAP7_75t_L g2344 ( 
.A1(n_2335),
.A2(n_2322),
.B1(n_2280),
.B2(n_2291),
.C1(n_2290),
.C2(n_2284),
.Y(n_2344)
);

NOR4xp25_ASAP7_75t_L g2345 ( 
.A(n_2332),
.B(n_2333),
.C(n_2325),
.D(n_2336),
.Y(n_2345)
);

OAI221xp5_ASAP7_75t_L g2346 ( 
.A1(n_2334),
.A2(n_2213),
.B1(n_2209),
.B2(n_2196),
.C(n_2291),
.Y(n_2346)
);

AOI211x1_ASAP7_75t_SL g2347 ( 
.A1(n_2334),
.A2(n_2248),
.B(n_2254),
.C(n_2185),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2329),
.B(n_2324),
.Y(n_2348)
);

AOI222xp33_ASAP7_75t_L g2349 ( 
.A1(n_2330),
.A2(n_2293),
.B1(n_2271),
.B2(n_2273),
.C1(n_2290),
.C2(n_2284),
.Y(n_2349)
);

OAI21xp33_ASAP7_75t_L g2350 ( 
.A1(n_2337),
.A2(n_2273),
.B(n_2271),
.Y(n_2350)
);

AOI211x1_ASAP7_75t_SL g2351 ( 
.A1(n_2338),
.A2(n_2248),
.B(n_2254),
.C(n_2185),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2339),
.B(n_2281),
.Y(n_2352)
);

OAI22xp5_ASAP7_75t_L g2353 ( 
.A1(n_2340),
.A2(n_2209),
.B1(n_2198),
.B2(n_2192),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2341),
.Y(n_2354)
);

A2O1A1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_2342),
.A2(n_2293),
.B(n_2281),
.C(n_2252),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2348),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2344),
.B(n_2218),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2343),
.A2(n_2209),
.B1(n_2198),
.B2(n_2212),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2346),
.A2(n_2269),
.B1(n_2263),
.B2(n_2207),
.Y(n_2359)
);

XNOR2x1_ASAP7_75t_L g2360 ( 
.A(n_2353),
.B(n_2345),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2356),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2354),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2351),
.B(n_2350),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2357),
.B(n_2349),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2355),
.B(n_2347),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2352),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2358),
.B(n_2218),
.Y(n_2367)
);

AOI221xp5_ASAP7_75t_L g2368 ( 
.A1(n_2364),
.A2(n_2359),
.B1(n_2245),
.B2(n_2266),
.C(n_2244),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2361),
.Y(n_2369)
);

INVxp67_ASAP7_75t_L g2370 ( 
.A(n_2360),
.Y(n_2370)
);

AND2x4_ASAP7_75t_L g2371 ( 
.A(n_2362),
.B(n_2207),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2367),
.B(n_2245),
.Y(n_2372)
);

NOR2xp67_ASAP7_75t_L g2373 ( 
.A(n_2366),
.B(n_2365),
.Y(n_2373)
);

OR5x1_ASAP7_75t_L g2374 ( 
.A(n_2373),
.B(n_2363),
.C(n_2365),
.D(n_2205),
.E(n_2189),
.Y(n_2374)
);

NOR3xp33_ASAP7_75t_SL g2375 ( 
.A(n_2369),
.B(n_2266),
.C(n_2256),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2371),
.B(n_2256),
.Y(n_2376)
);

AND4x2_ASAP7_75t_L g2377 ( 
.A(n_2368),
.B(n_2159),
.C(n_2189),
.D(n_2205),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2376),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2378),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2379),
.B(n_2370),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2379),
.Y(n_2381)
);

OAI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2381),
.A2(n_2372),
.B1(n_2375),
.B2(n_2377),
.Y(n_2382)
);

XNOR2xp5_ASAP7_75t_L g2383 ( 
.A(n_2380),
.B(n_2374),
.Y(n_2383)
);

NOR3xp33_ASAP7_75t_L g2384 ( 
.A(n_2382),
.B(n_2166),
.C(n_2269),
.Y(n_2384)
);

OAI22xp33_ASAP7_75t_L g2385 ( 
.A1(n_2383),
.A2(n_2263),
.B1(n_2166),
.B2(n_2224),
.Y(n_2385)
);

AOI22x1_ASAP7_75t_L g2386 ( 
.A1(n_2384),
.A2(n_2166),
.B1(n_2220),
.B2(n_2224),
.Y(n_2386)
);

OAI21x1_ASAP7_75t_L g2387 ( 
.A1(n_2386),
.A2(n_2385),
.B(n_2220),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2387),
.B(n_2146),
.Y(n_2388)
);

AOI22x1_ASAP7_75t_L g2389 ( 
.A1(n_2388),
.A2(n_2146),
.B1(n_2148),
.B2(n_2155),
.Y(n_2389)
);

OAI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2389),
.A2(n_2146),
.B1(n_2156),
.B2(n_2172),
.Y(n_2390)
);

AOI211xp5_ASAP7_75t_L g2391 ( 
.A1(n_2390),
.A2(n_1798),
.B(n_1809),
.C(n_2146),
.Y(n_2391)
);


endmodule