module fake_aes_511_n_710 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_710);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_710;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g80 ( .A(n_40), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_38), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_59), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_77), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_5), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_30), .Y(n_85) );
CKINVDCx14_ASAP7_75t_R g86 ( .A(n_2), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_1), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_10), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_37), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_49), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_36), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_64), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_11), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_67), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_39), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_35), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_20), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_46), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_32), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_75), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_26), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_56), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_44), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_27), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_50), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_16), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_4), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_71), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_41), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_52), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_78), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_6), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_3), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_61), .Y(n_122) );
CKINVDCx14_ASAP7_75t_R g123 ( .A(n_33), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_79), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_65), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_23), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_53), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_16), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_111), .B(n_0), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_126), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_126), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_111), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_126), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_126), .B(n_25), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
INVxp67_ASAP7_75t_SL g136 ( .A(n_84), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_80), .B(n_0), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_81), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_81), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_98), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_86), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_108), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_90), .B(n_1), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_93), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_112), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_112), .B(n_3), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_87), .B(n_4), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_93), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_100), .B(n_29), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_87), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_97), .B(n_5), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_97), .B(n_6), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_90), .B(n_7), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_102), .B(n_7), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_100), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
BUFx8_ASAP7_75t_L g167 ( .A(n_113), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_115), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_115), .Y(n_169) );
BUFx8_ASAP7_75t_L g170 ( .A(n_116), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_102), .B(n_8), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_101), .B(n_9), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
INVx6_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_136), .B(n_117), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_148), .B(n_119), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_135), .B(n_123), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_135), .B(n_82), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_138), .B(n_119), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_167), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_138), .B(n_83), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
NOR2x1_ASAP7_75t_L g192 ( .A(n_140), .B(n_116), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_140), .B(n_127), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
AO22x2_ASAP7_75t_L g198 ( .A1(n_172), .A2(n_171), .B1(n_163), .B2(n_164), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_160), .B(n_128), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_172), .B(n_124), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_131), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_145), .B(n_127), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_130), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_131), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_131), .B(n_124), .Y(n_205) );
AO22x2_ASAP7_75t_L g206 ( .A1(n_163), .A2(n_128), .B1(n_101), .B2(n_106), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_145), .B(n_114), .Y(n_207) );
NAND3xp33_ASAP7_75t_L g208 ( .A(n_167), .B(n_170), .C(n_129), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_130), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_133), .B(n_125), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_130), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_129), .B(n_88), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_164), .B(n_106), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_141), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_133), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_133), .B(n_125), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_152), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_152), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_165), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_147), .B(n_85), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_171), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_147), .B(n_121), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_154), .B(n_121), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_154), .B(n_120), .Y(n_224) );
INVx1_ASAP7_75t_SL g225 ( .A(n_151), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_152), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_158), .Y(n_227) );
OR2x2_ASAP7_75t_L g228 ( .A(n_161), .B(n_114), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_143), .Y(n_229) );
AND2x6_ASAP7_75t_L g230 ( .A(n_143), .B(n_120), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_141), .Y(n_231) );
INVx4_ASAP7_75t_L g232 ( .A(n_134), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_141), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_232), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_178), .B(n_170), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_198), .A2(n_170), .B1(n_167), .B2(n_94), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_178), .B(n_167), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_232), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_184), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_213), .B(n_166), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_188), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_198), .A2(n_221), .B1(n_213), .B2(n_206), .Y(n_243) );
INVx4_ASAP7_75t_L g244 ( .A(n_188), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_183), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_183), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_230), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_198), .A2(n_170), .B1(n_107), .B2(n_166), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_173), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_195), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_173), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_185), .B(n_189), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_206), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_199), .B(n_161), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_222), .B(n_162), .Y(n_256) );
BUFx4f_ASAP7_75t_L g257 ( .A(n_200), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_230), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_221), .A2(n_159), .B1(n_134), .B2(n_162), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_222), .B(n_155), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_229), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_228), .A2(n_118), .B(n_169), .C(n_158), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_223), .B(n_159), .Y(n_263) );
INVx8_ASAP7_75t_L g264 ( .A(n_200), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_223), .B(n_200), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_207), .B(n_118), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_230), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_176), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_200), .B(n_159), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_204), .Y(n_271) );
AND3x1_ASAP7_75t_L g272 ( .A(n_180), .B(n_155), .C(n_139), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_230), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_176), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_225), .B(n_155), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_207), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_207), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_215), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_208), .B(n_155), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_175), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_179), .A2(n_169), .B1(n_158), .B2(n_159), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_206), .B(n_169), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_217), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_180), .B(n_110), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_191), .A2(n_159), .B1(n_134), .B2(n_122), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_173), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_182), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_173), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_193), .B(n_168), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_212), .Y(n_292) );
OAI22xp5_ASAP7_75t_SL g293 ( .A1(n_197), .A2(n_104), .B1(n_96), .B2(n_103), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_218), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
BUFx4f_ASAP7_75t_L g297 ( .A(n_205), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_196), .B(n_159), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_192), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_256), .B(n_255), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_295), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_277), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_250), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_283), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_240), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_268), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_292), .B(n_181), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_283), .A2(n_254), .B1(n_255), .B2(n_256), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_264), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_241), .B(n_186), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_257), .B(n_196), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_250), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_298), .A2(n_220), .B(n_190), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_271), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_241), .B(n_202), .Y(n_318) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_257), .B(n_202), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_283), .B(n_187), .Y(n_320) );
BUFx12f_ASAP7_75t_L g321 ( .A(n_261), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_277), .B(n_194), .Y(n_322) );
NOR2x1_ASAP7_75t_SL g323 ( .A(n_277), .B(n_194), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_254), .A2(n_210), .B1(n_216), .B2(n_205), .Y(n_324) );
INVx5_ASAP7_75t_L g325 ( .A(n_264), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_247), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_285), .A2(n_187), .B(n_142), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_279), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_285), .B(n_99), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_245), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_266), .B(n_205), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_247), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_244), .B(n_134), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
OAI22x1_ASAP7_75t_L g335 ( .A1(n_248), .A2(n_137), .B1(n_142), .B2(n_144), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_243), .A2(n_205), .B1(n_216), .B2(n_210), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_298), .A2(n_209), .B(n_203), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_234), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_284), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_266), .B(n_144), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_236), .B(n_205), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_294), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_276), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_234), .Y(n_344) );
INVxp67_ASAP7_75t_L g345 ( .A(n_260), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_260), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_273), .B(n_168), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_278), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_236), .B(n_210), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_234), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_244), .B(n_134), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_238), .B(n_105), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_303), .A2(n_238), .B1(n_280), .B2(n_293), .Y(n_353) );
INVx5_ASAP7_75t_L g354 ( .A(n_325), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_306), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_312), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_309), .A2(n_272), .B1(n_259), .B2(n_237), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_314), .A2(n_280), .B1(n_242), .B2(n_291), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_320), .A2(n_242), .B1(n_275), .B2(n_265), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_325), .Y(n_360) );
AO21x2_ASAP7_75t_L g361 ( .A1(n_315), .A2(n_286), .B(n_263), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_320), .A2(n_275), .B1(n_265), .B2(n_235), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_312), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_337), .A2(n_262), .B(n_282), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_304), .A2(n_282), .B1(n_262), .B2(n_296), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_325), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
AOI21xp5_ASAP7_75t_SL g369 ( .A1(n_304), .A2(n_273), .B(n_258), .Y(n_369) );
NOR2xp33_ASAP7_75t_SL g370 ( .A(n_325), .B(n_247), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g371 ( .A1(n_300), .A2(n_263), .B(n_270), .Y(n_371) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_325), .B(n_252), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
INVxp33_ASAP7_75t_L g374 ( .A(n_307), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_305), .A2(n_274), .B1(n_269), .B2(n_299), .Y(n_375) );
NOR4xp25_ASAP7_75t_L g376 ( .A(n_327), .B(n_137), .C(n_142), .D(n_144), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_301), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_341), .A2(n_270), .B(n_253), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_301), .Y(n_380) );
NAND3xp33_ASAP7_75t_L g381 ( .A(n_349), .B(n_146), .C(n_141), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_305), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_318), .A2(n_253), .B1(n_137), .B2(n_150), .C(n_290), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_348), .B(n_252), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_357), .A2(n_335), .B1(n_352), .B2(n_329), .Y(n_386) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_358), .A2(n_345), .B(n_311), .C(n_346), .Y(n_387) );
AOI22xp5_ASAP7_75t_SL g388 ( .A1(n_357), .A2(n_335), .B1(n_351), .B2(n_333), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_374), .A2(n_340), .B(n_331), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_383), .A2(n_319), .B1(n_321), .B2(n_333), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_353), .A2(n_343), .B1(n_348), .B2(n_317), .C(n_328), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
NAND2x1p5_ASAP7_75t_L g393 ( .A(n_354), .B(n_326), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_383), .A2(n_340), .B1(n_336), .B2(n_321), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_359), .A2(n_319), .B1(n_351), .B2(n_333), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_354), .B(n_317), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_356), .B(n_328), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_364), .A2(n_342), .B1(n_324), .B2(n_334), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_364), .A2(n_377), .B1(n_368), .B2(n_378), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_354), .A2(n_351), .B1(n_323), .B2(n_308), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g404 ( .A1(n_375), .A2(n_150), .B(n_290), .C(n_165), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_368), .A2(n_342), .B1(n_134), .B2(n_159), .Y(n_405) );
NOR2x1_ASAP7_75t_SL g406 ( .A(n_354), .B(n_326), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_355), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_377), .A2(n_134), .B1(n_159), .B2(n_334), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_366), .A2(n_216), .B1(n_210), .B2(n_134), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_378), .A2(n_330), .B1(n_210), .B2(n_216), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_362), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_380), .A2(n_150), .B1(n_297), .B2(n_330), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_354), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_380), .B(n_323), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_398), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_392), .B(n_362), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_387), .A2(n_366), .B1(n_363), .B2(n_376), .C(n_384), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_392), .B(n_362), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_392), .B(n_373), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_394), .B(n_373), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_394), .B(n_373), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_396), .A2(n_361), .B1(n_384), .B2(n_354), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_391), .A2(n_376), .B1(n_371), .B2(n_168), .C(n_165), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_395), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_409), .A2(n_382), .B1(n_385), .B2(n_371), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_386), .A2(n_361), .B1(n_367), .B2(n_360), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_394), .A2(n_382), .B(n_381), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_390), .A2(n_385), .B1(n_313), .B2(n_381), .C(n_360), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
NAND4xp25_ASAP7_75t_SL g432 ( .A(n_397), .B(n_369), .C(n_382), .D(n_11), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_389), .A2(n_361), .B1(n_367), .B2(n_216), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_407), .B(n_365), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_361), .B1(n_367), .B2(n_330), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g436 ( .A1(n_398), .A2(n_369), .B(n_165), .C(n_168), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_407), .B(n_365), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_403), .A2(n_365), .B1(n_379), .B2(n_165), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_403), .A2(n_165), .B1(n_168), .B2(n_350), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_388), .A2(n_370), .B1(n_372), .B2(n_313), .Y(n_440) );
OA222x2_ASAP7_75t_L g441 ( .A1(n_403), .A2(n_308), .B1(n_350), .B2(n_344), .C1(n_338), .C2(n_302), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_413), .Y(n_442) );
AOI33xp33_ASAP7_75t_L g443 ( .A1(n_401), .A2(n_214), .A3(n_231), .B1(n_233), .B2(n_209), .B3(n_203), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_411), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_411), .B(n_168), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_388), .B(n_9), .C(n_10), .D(n_12), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_411), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_409), .A2(n_372), .B1(n_297), .B2(n_313), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
AO221x2_ASAP7_75t_L g450 ( .A1(n_427), .A2(n_412), .B1(n_400), .B2(n_414), .C(n_15), .Y(n_450) );
OAI21xp5_ASAP7_75t_SL g451 ( .A1(n_446), .A2(n_402), .B(n_393), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_416), .B(n_413), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_446), .B(n_404), .C(n_400), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_437), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_416), .B(n_413), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_431), .B(n_406), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_437), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_426), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_431), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_444), .B(n_406), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_444), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_426), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_447), .B(n_393), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_419), .A2(n_412), .B(n_408), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_432), .A2(n_410), .B1(n_370), .B2(n_405), .Y(n_465) );
AOI33xp33_ASAP7_75t_L g466 ( .A1(n_428), .A2(n_231), .A3(n_233), .B1(n_214), .B2(n_17), .B3(n_18), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_449), .B(n_393), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_432), .A2(n_149), .B1(n_146), .B2(n_141), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_449), .B(n_149), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_427), .A2(n_149), .B1(n_146), .B2(n_141), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_448), .B(n_372), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_447), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_417), .B(n_149), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_417), .B(n_149), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_420), .B(n_149), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_420), .B(n_12), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
OAI21x1_ASAP7_75t_L g478 ( .A1(n_429), .A2(n_347), .B(n_322), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_434), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_421), .B(n_13), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_421), .B(n_13), .Y(n_481) );
AOI211xp5_ASAP7_75t_SL g482 ( .A1(n_436), .A2(n_350), .B(n_344), .C(n_338), .Y(n_482) );
NAND2xp33_ASAP7_75t_SL g483 ( .A(n_418), .B(n_267), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_422), .B(n_14), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_423), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_415), .B(n_14), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_425), .A2(n_344), .B1(n_338), .B2(n_322), .Y(n_488) );
AND2x2_ASAP7_75t_SL g489 ( .A(n_424), .B(n_267), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_423), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_415), .B(n_17), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_442), .B(n_19), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_442), .B(n_19), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_442), .B(n_20), .Y(n_495) );
OAI221xp5_ASAP7_75t_L g496 ( .A1(n_433), .A2(n_322), .B1(n_347), .B2(n_146), .C(n_109), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_442), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_458), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_479), .B(n_477), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g501 ( .A(n_466), .B(n_436), .C(n_440), .D(n_435), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_459), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_456), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_479), .B(n_438), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_498), .B(n_443), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_477), .B(n_441), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_477), .B(n_441), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_458), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_462), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_476), .B(n_21), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_462), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_476), .B(n_21), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_495), .B(n_430), .C(n_448), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_480), .B(n_146), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_472), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_454), .B(n_146), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_454), .B(n_439), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_480), .B(n_246), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_454), .B(n_22), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_459), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_457), .B(n_24), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_457), .B(n_28), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_453), .A2(n_219), .B1(n_177), .B2(n_211), .C(n_174), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_481), .B(n_31), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_481), .B(n_34), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_457), .B(n_42), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_459), .B(n_43), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_461), .B(n_45), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_461), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_485), .B(n_47), .Y(n_532) );
NAND4xp75_ASAP7_75t_L g533 ( .A(n_489), .B(n_310), .C(n_51), .D(n_55), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_485), .B(n_48), .Y(n_534) );
AOI211xp5_ASAP7_75t_L g535 ( .A1(n_451), .A2(n_177), .B(n_211), .C(n_174), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_461), .B(n_211), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_484), .Y(n_537) );
AOI211xp5_ASAP7_75t_SL g538 ( .A1(n_451), .A2(n_302), .B(n_58), .C(n_60), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_484), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_486), .B(n_57), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_486), .B(n_490), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_490), .B(n_62), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_460), .B(n_66), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_469), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_460), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g546 ( .A1(n_482), .A2(n_302), .B(n_177), .C(n_174), .Y(n_546) );
NOR2x1p5_ASAP7_75t_L g547 ( .A(n_452), .B(n_252), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_463), .B(n_68), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_469), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_463), .B(n_72), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_494), .B(n_73), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_492), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_455), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_467), .B(n_74), .Y(n_554) );
NAND5xp2_ASAP7_75t_L g555 ( .A(n_482), .B(n_347), .C(n_76), .D(n_310), .E(n_258), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_452), .B(n_267), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_467), .B(n_174), .Y(n_557) );
NAND4xp25_ASAP7_75t_L g558 ( .A(n_538), .B(n_468), .C(n_464), .D(n_465), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_506), .A2(n_489), .B(n_470), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_499), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_545), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_541), .B(n_497), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_541), .B(n_497), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_503), .B(n_455), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_503), .B(n_515), .Y(n_565) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_555), .A2(n_493), .B(n_492), .C(n_491), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_501), .A2(n_450), .B1(n_489), .B2(n_464), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_553), .B(n_494), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_502), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_545), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_553), .B(n_450), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_552), .B(n_487), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_513), .A2(n_450), .B1(n_493), .B2(n_491), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_502), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_499), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_510), .A2(n_450), .B1(n_471), .B2(n_487), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_508), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_508), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_500), .B(n_475), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_539), .B(n_475), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_509), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_506), .B(n_471), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_552), .B(n_474), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_509), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_502), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_537), .B(n_474), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_511), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_539), .B(n_473), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_500), .B(n_473), .Y(n_589) );
NOR2xp67_ASAP7_75t_L g590 ( .A(n_546), .B(n_496), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_537), .B(n_471), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_522), .Y(n_592) );
NOR4xp75_ASAP7_75t_L g593 ( .A(n_533), .B(n_471), .C(n_483), .D(n_465), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_522), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_507), .B(n_471), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_535), .B(n_488), .C(n_211), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_511), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_537), .B(n_488), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_531), .B(n_478), .Y(n_599) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_533), .B(n_332), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_516), .B(n_478), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_512), .B(n_219), .C(n_251), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_507), .B(n_177), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_531), .B(n_332), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_535), .A2(n_332), .B(n_326), .Y(n_605) );
OAI211xp5_ASAP7_75t_L g606 ( .A1(n_538), .A2(n_258), .B(n_332), .C(n_326), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_543), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_504), .B(n_326), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_504), .B(n_332), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_516), .B(n_249), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_544), .A2(n_287), .B1(n_289), .B2(n_251), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_562), .B(n_520), .Y(n_612) );
NAND2xp33_ASAP7_75t_SL g613 ( .A(n_565), .B(n_547), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_596), .A2(n_505), .B(n_543), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_563), .B(n_520), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_574), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_595), .B(n_517), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_560), .Y(n_618) );
OA211x2_ASAP7_75t_L g619 ( .A1(n_567), .A2(n_532), .B(n_526), .C(n_527), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_575), .Y(n_620) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_567), .B(n_550), .C(n_548), .D(n_534), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_577), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_578), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_581), .Y(n_624) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_569), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_571), .B(n_544), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_558), .B(n_514), .C(n_540), .Y(n_627) );
CKINVDCx14_ASAP7_75t_R g628 ( .A(n_579), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_568), .B(n_549), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_584), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_587), .B(n_549), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_606), .B(n_521), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_561), .B(n_519), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_607), .B(n_521), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_597), .B(n_517), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_576), .A2(n_548), .B(n_550), .C(n_542), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_570), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_589), .B(n_518), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_595), .B(n_518), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_572), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_592), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_592), .B(n_542), .Y(n_642) );
OAI32xp33_ASAP7_75t_L g643 ( .A1(n_564), .A2(n_551), .A3(n_529), .B1(n_530), .B2(n_554), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_594), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_569), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_594), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_559), .B(n_521), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_580), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_583), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_588), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_576), .B(n_525), .C(n_556), .D(n_551), .Y(n_651) );
XNOR2x2_ASAP7_75t_L g652 ( .A(n_593), .B(n_524), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_574), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_585), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_573), .A2(n_530), .B(n_529), .C(n_524), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_573), .A2(n_547), .B1(n_521), .B2(n_528), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_585), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_599), .Y(n_658) );
INVxp67_ASAP7_75t_SL g659 ( .A(n_603), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_586), .B(n_536), .Y(n_660) );
XOR2xp5_ASAP7_75t_L g661 ( .A(n_582), .B(n_523), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_591), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_582), .A2(n_523), .B1(n_528), .B2(n_557), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_582), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_601), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_598), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_610), .Y(n_667) );
XNOR2xp5_ASAP7_75t_L g668 ( .A(n_566), .B(n_536), .Y(n_668) );
AO21x1_ASAP7_75t_L g669 ( .A1(n_605), .A2(n_249), .B(n_287), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_610), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_590), .A2(n_239), .B1(n_287), .B2(n_289), .Y(n_671) );
AOI22xp5_ASAP7_75t_SL g672 ( .A1(n_608), .A2(n_239), .B1(n_289), .B2(n_600), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_609), .A2(n_604), .B1(n_608), .B2(n_602), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g674 ( .A1(n_602), .A2(n_239), .B(n_611), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_662), .B(n_666), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_628), .A2(n_636), .B1(n_656), .B2(n_664), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_621), .A2(n_619), .B1(n_628), .B2(n_647), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_641), .Y(n_678) );
CKINVDCx16_ASAP7_75t_R g679 ( .A(n_637), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_674), .A2(n_614), .B(n_647), .C(n_656), .Y(n_680) );
OAI21xp5_ASAP7_75t_SL g681 ( .A1(n_668), .A2(n_655), .B(n_632), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_613), .A2(n_632), .B(n_659), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_613), .A2(n_659), .B1(n_640), .B2(n_627), .C(n_626), .Y(n_683) );
AOI221x1_ASAP7_75t_L g684 ( .A1(n_633), .A2(n_651), .B1(n_648), .B2(n_650), .C(n_630), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g685 ( .A1(n_637), .A2(n_634), .B(n_671), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_612), .A2(n_615), .B1(n_649), .B2(n_643), .C(n_638), .Y(n_686) );
INVxp67_ASAP7_75t_SL g687 ( .A(n_645), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g688 ( .A1(n_645), .A2(n_663), .B1(n_642), .B2(n_634), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_676), .A2(n_673), .B1(n_658), .B2(n_625), .C(n_629), .Y(n_689) );
OAI311xp33_ASAP7_75t_L g690 ( .A1(n_681), .A2(n_652), .A3(n_639), .B1(n_631), .C1(n_635), .Y(n_690) );
OAI211xp5_ASAP7_75t_L g691 ( .A1(n_680), .A2(n_661), .B(n_658), .C(n_665), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_675), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_683), .A2(n_667), .B1(n_670), .B2(n_673), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_677), .A2(n_671), .B(n_624), .C(n_618), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g695 ( .A1(n_688), .A2(n_669), .B(n_617), .C(n_665), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_679), .A2(n_672), .B1(n_660), .B2(n_617), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_692), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_693), .B(n_684), .Y(n_698) );
OAI211xp5_ASAP7_75t_SL g699 ( .A1(n_695), .A2(n_686), .B(n_682), .C(n_687), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_691), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_690), .A2(n_687), .B(n_685), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_697), .B(n_678), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_701), .A2(n_689), .B1(n_694), .B2(n_696), .C(n_622), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_700), .B(n_611), .C(n_623), .D(n_620), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_702), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_703), .A2(n_698), .B1(n_699), .B2(n_646), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_704), .B1(n_644), .B2(n_653), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_SL g708 ( .A1(n_707), .A2(n_705), .B(n_657), .C(n_654), .Y(n_708) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_708), .B(n_616), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g710 ( .A1(n_709), .A2(n_616), .B(n_654), .Y(n_710) );
endmodule