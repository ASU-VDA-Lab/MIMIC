module fake_jpeg_4157_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_16),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_55),
.B1(n_33),
.B2(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_29),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_52),
.B(n_68),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_67),
.B1(n_26),
.B2(n_24),
.Y(n_85)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_65),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_31),
.B1(n_41),
.B2(n_35),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_18),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_18),
.B(n_17),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_21),
.B1(n_29),
.B2(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_27),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_41),
.B1(n_27),
.B2(n_45),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_85),
.B1(n_21),
.B2(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_46),
.B1(n_45),
.B2(n_38),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_53),
.B1(n_59),
.B2(n_57),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_24),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_76),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_36),
.B1(n_19),
.B2(n_24),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_36),
.B1(n_21),
.B2(n_26),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_69),
.B(n_56),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_116),
.B1(n_75),
.B2(n_87),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_50),
.B1(n_66),
.B2(n_59),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_101),
.A2(n_122),
.B1(n_94),
.B2(n_99),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_120),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_127),
.B1(n_85),
.B2(n_83),
.Y(n_144)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_117),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_68),
.C(n_61),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_81),
.C(n_75),
.Y(n_145)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_123),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_59),
.B1(n_46),
.B2(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_126),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_56),
.B(n_39),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_116),
.B(n_126),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_84),
.A2(n_54),
.B1(n_20),
.B2(n_22),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_131),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_88),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_108),
.Y(n_172)
);

BUFx4f_ASAP7_75t_SL g131 ( 
.A(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_133),
.B(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_154),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_146),
.B(n_155),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_89),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_145),
.C(n_149),
.Y(n_161)
);

BUFx24_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_77),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_151),
.B1(n_122),
.B2(n_109),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_98),
.B(n_91),
.C(n_93),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_157),
.B1(n_74),
.B2(n_63),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_87),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_150),
.B(n_63),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_96),
.B1(n_72),
.B2(n_74),
.Y(n_151)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_96),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_72),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_110),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_39),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_164),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_124),
.B1(n_99),
.B2(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_178),
.B1(n_190),
.B2(n_128),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_125),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_165),
.B(n_167),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_110),
.C(n_100),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_155),
.A3(n_152),
.B1(n_153),
.B2(n_61),
.Y(n_205)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_171),
.B1(n_183),
.B2(n_185),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_109),
.B1(n_108),
.B2(n_63),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_186),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_119),
.B(n_20),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_131),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_174),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_90),
.B(n_1),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_177),
.CI(n_0),
.CON(n_204),
.SN(n_204)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_141),
.B(n_12),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_22),
.B1(n_25),
.B2(n_37),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_145),
.C(n_149),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_144),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_25),
.B1(n_37),
.B2(n_61),
.Y(n_190)
);

AND2x4_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_146),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_205),
.B(n_209),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_161),
.B1(n_179),
.B2(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_211),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_196),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_201),
.C(n_202),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_163),
.B(n_130),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_217),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_212),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_30),
.B(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_71),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_215),
.C(n_140),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_142),
.B1(n_30),
.B2(n_9),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_214),
.A2(n_190),
.B1(n_164),
.B2(n_165),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_161),
.B(n_140),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_238),
.Y(n_248)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_185),
.B1(n_183),
.B2(n_172),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_231),
.B(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_192),
.A2(n_178),
.B1(n_167),
.B2(n_169),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_236),
.B1(n_195),
.B2(n_193),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_194),
.B1(n_208),
.B2(n_209),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_246),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_159),
.B1(n_172),
.B2(n_176),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_173),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_242),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_177),
.B1(n_180),
.B2(n_174),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_180),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_3),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_215),
.C(n_204),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_197),
.B(n_30),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_266),
.B1(n_233),
.B2(n_231),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_201),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_255),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_258),
.C(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_204),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_238),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_1),
.C(n_2),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_7),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_241),
.B1(n_227),
.B2(n_221),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_234),
.C(n_237),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_8),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_221),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_3),
.B(n_4),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_282),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_274),
.C(n_266),
.Y(n_289)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_278),
.B(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_243),
.C(n_226),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_252),
.C(n_259),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_225),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_283),
.Y(n_290)
);

NOR4xp25_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_225),
.C(n_223),
.D(n_228),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_276),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_242),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_281),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_247),
.A2(n_223),
.B(n_229),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_229),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_230),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_260),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_295),
.B(n_5),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_254),
.C(n_250),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_249),
.B1(n_247),
.B2(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_256),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_268),
.B1(n_271),
.B2(n_275),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_258),
.B1(n_265),
.B2(n_3),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_296),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_280),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_306),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_4),
.Y(n_301)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_286),
.C(n_290),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_305),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_4),
.Y(n_304)
);

AOI32xp33_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_8),
.A3(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_285),
.B(n_6),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_288),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_287),
.A2(n_6),
.B(n_7),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_16),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_311),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_10),
.B1(n_12),
.B2(n_15),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_10),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_316),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.C(n_300),
.Y(n_322)
);

AOI31xp33_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_304),
.A3(n_303),
.B(n_300),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_320),
.A2(n_312),
.B(n_314),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_299),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_317),
.B(n_315),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_321),
.B(n_328),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_327),
.C(n_324),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_16),
.Y(n_332)
);


endmodule