module fake_jpeg_15173_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_15),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_44),
.C(n_45),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_14),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_16),
.B1(n_31),
.B2(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_18),
.B1(n_24),
.B2(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_56),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_46),
.C(n_38),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_25),
.C(n_22),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_17),
.B1(n_16),
.B2(n_31),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_42),
.B1(n_24),
.B2(n_34),
.Y(n_91)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_23),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_26),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_27),
.B1(n_25),
.B2(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_16),
.B1(n_19),
.B2(n_33),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_76),
.B1(n_51),
.B2(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_75),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_81),
.Y(n_120)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_47),
.B1(n_18),
.B2(n_33),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_82),
.A2(n_89),
.B1(n_91),
.B2(n_94),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_33),
.B1(n_24),
.B2(n_26),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_23),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_95),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_48),
.B1(n_42),
.B2(n_47),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_88),
.A2(n_96),
.B1(n_101),
.B2(n_103),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_47),
.B1(n_18),
.B2(n_33),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_104),
.C(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_22),
.Y(n_95)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_45),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_29),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_25),
.B1(n_22),
.B2(n_46),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_111),
.Y(n_138)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_27),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_27),
.B1(n_22),
.B2(n_34),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_34),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_21),
.B1(n_30),
.B2(n_29),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_20),
.B(n_32),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_53),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_77),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_122),
.C(n_114),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_88),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_77),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_124),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_75),
.B(n_21),
.C(n_20),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_137),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_20),
.B(n_29),
.C(n_30),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_111),
.B(n_105),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_70),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_88),
.Y(n_165)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_84),
.A3(n_101),
.B1(n_108),
.B2(n_90),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_171),
.A3(n_163),
.B1(n_149),
.B2(n_169),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_84),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_149),
.B(n_167),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_104),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_134),
.C(n_132),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_91),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_162),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_103),
.B1(n_88),
.B2(n_50),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_177),
.B1(n_144),
.B2(n_119),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_170),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_103),
.B1(n_110),
.B2(n_81),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_117),
.B1(n_119),
.B2(n_127),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_171),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_99),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_166),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_99),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_93),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_169),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_140),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

XOR2x2_ASAP7_75t_SL g171 ( 
.A(n_122),
.B(n_78),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_86),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_59),
.Y(n_203)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_86),
.B(n_80),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_137),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_115),
.B(n_0),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_50),
.B1(n_79),
.B2(n_97),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_181),
.B(n_187),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_189),
.B1(n_211),
.B2(n_178),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_162),
.B1(n_175),
.B2(n_146),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_191),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_132),
.B1(n_131),
.B2(n_124),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g190 ( 
.A(n_156),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_190),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_155),
.C(n_174),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_213),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_135),
.B1(n_128),
.B2(n_118),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_202),
.B1(n_205),
.B2(n_184),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_128),
.B1(n_118),
.B2(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_206),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_59),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_126),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_150),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_53),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_62),
.B1(n_59),
.B2(n_49),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_214),
.B(n_216),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_151),
.C(n_161),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_215),
.B(n_238),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_192),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_220),
.B1(n_223),
.B2(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_236),
.C(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_162),
.B1(n_185),
.B2(n_194),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_221),
.A2(n_226),
.B1(n_200),
.B2(n_212),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_175),
.B1(n_177),
.B2(n_158),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_148),
.B1(n_153),
.B2(n_147),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_153),
.B1(n_166),
.B2(n_172),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_147),
.B1(n_154),
.B2(n_173),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_230),
.B1(n_204),
.B2(n_187),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_154),
.B1(n_145),
.B2(n_62),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_12),
.C(n_11),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_11),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_9),
.C(n_8),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g241 ( 
.A1(n_195),
.A2(n_9),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_197),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_209),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_SL g285 ( 
.A1(n_243),
.A2(n_241),
.B(n_2),
.C(n_3),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_193),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_263),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_184),
.B(n_180),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_251),
.B1(n_257),
.B2(n_264),
.Y(n_277)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_206),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_210),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_259),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_198),
.C(n_202),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_256),
.C(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_199),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_182),
.B1(n_188),
.B2(n_197),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_234),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_224),
.B(n_203),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_235),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_262),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_230),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_212),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_225),
.A2(n_0),
.B(n_1),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_228),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_283),
.C(n_252),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_273),
.B(n_243),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_1),
.B(n_2),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_281),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_285),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_1),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_256),
.C(n_254),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_284),
.C(n_252),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_231),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_240),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_245),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_215),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_236),
.C(n_229),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_289),
.C(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_263),
.C(n_249),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.C(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_248),
.C(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_243),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_242),
.C(n_258),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_298),
.C(n_276),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_222),
.Y(n_297)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_288),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_306),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_270),
.C(n_271),
.Y(n_306)
);

XOR2x2_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_280),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_286),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_314),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_268),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_287),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_285),
.Y(n_323)
);

XOR2x1_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_280),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_296),
.B1(n_295),
.B2(n_298),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_267),
.C(n_285),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_320),
.C(n_4),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_299),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_325),
.C(n_303),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_285),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_3),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_2),
.Y(n_325)
);

AOI322xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_313),
.A3(n_308),
.B1(n_305),
.B2(n_306),
.C1(n_314),
.C2(n_315),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_330),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_322),
.C(n_325),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_7),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_3),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_332),
.B(n_318),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_333),
.B(n_332),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_4),
.C(n_5),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_338),
.A2(n_334),
.B(n_337),
.Y(n_340)
);

AOI321xp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_5),
.A3(n_6),
.B1(n_339),
.B2(n_333),
.C(n_302),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_5),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_6),
.Y(n_343)
);


endmodule