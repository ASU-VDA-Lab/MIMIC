module real_jpeg_30419_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_216;
wire n_179;
wire n_167;
wire n_244;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_0),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_0),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_1),
.B(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_6),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_1),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_1),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_6),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_7),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_8),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_8),
.B(n_110),
.Y(n_109)
);

NAND2x1_ASAP7_75t_L g124 ( 
.A(n_8),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_8),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_8),
.B(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_10),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_10),
.B(n_128),
.Y(n_127)
);

AND2x4_ASAP7_75t_SL g148 ( 
.A(n_10),
.B(n_29),
.Y(n_148)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_11),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_12),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_13),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_14),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_165),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_162),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_19),
.B(n_137),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_77),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_40),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_30),
.C(n_33),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_22),
.A2(n_23),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_24),
.A2(n_27),
.B1(n_28),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_24),
.Y(n_161)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_30),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_59),
.Y(n_40)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_52),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVxp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

NOR2x1_ASAP7_75t_R g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_61),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_61),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_76),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_69),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

OR2x2_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_118),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.C(n_102),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_85),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_84),
.Y(n_213)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_97),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_252)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_94),
.B(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_109),
.C(n_113),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_117),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_115),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_133),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_127),
.Y(n_132)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.C(n_146),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_138),
.A2(n_139),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_142),
.B(n_146),
.Y(n_264)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.C(n_159),
.Y(n_146)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_147),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_148),
.B(n_150),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_154),
.A2(n_159),
.B1(n_160),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_154),
.Y(n_256)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_260),
.B(n_265),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_244),
.B(n_259),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_222),
.B(n_243),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_204),
.B(n_221),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_195),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_195),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_182),
.B2(n_183),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_178),
.C(n_182),
.Y(n_223)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_190),
.B2(n_191),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_190),
.Y(n_227)
);

NOR2x1_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx4f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_214),
.B(n_220),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_219),
.Y(n_220)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_224),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_236),
.C(n_238),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_246),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_253),
.B1(n_257),
.B2(n_258),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_250),
.C(n_258),
.Y(n_261)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);


endmodule