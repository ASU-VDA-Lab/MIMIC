module fake_jpeg_2524_n_149 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_149);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_2),
.B(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_30),
.B(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_41),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_23),
.B(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_11),
.B(n_3),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_25),
.B1(n_5),
.B2(n_6),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_14),
.Y(n_57)
);

OA22x2_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_19),
.B1(n_25),
.B2(n_27),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_52),
.B(n_66),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_27),
.C(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_76),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_18),
.B1(n_25),
.B2(n_12),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_73),
.B1(n_34),
.B2(n_36),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_30),
.A2(n_18),
.B1(n_21),
.B2(n_12),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_11),
.B1(n_14),
.B2(n_21),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_32),
.B1(n_43),
.B2(n_28),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_45),
.B1(n_33),
.B2(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_45),
.B1(n_32),
.B2(n_43),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_82),
.B1(n_69),
.B2(n_56),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_85),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_88),
.C(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_37),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_68),
.B1(n_59),
.B2(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_51),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_79),
.C(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_50),
.B1(n_56),
.B2(n_74),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_79),
.B1(n_84),
.B2(n_95),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_93),
.B(n_90),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_121),
.B(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_118),
.B(n_120),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_54),
.C(n_81),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_81),
.B(n_100),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_126),
.B(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_97),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_129),
.B1(n_114),
.B2(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_105),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_134),
.B1(n_136),
.B2(n_132),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_119),
.B(n_122),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_103),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_108),
.C(n_118),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_103),
.C(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_117),
.B1(n_112),
.B2(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_112),
.B1(n_110),
.B2(n_98),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_135),
.B1(n_124),
.B2(n_129),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_139),
.C(n_140),
.Y(n_142)
);

XOR2x2_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_139),
.Y(n_144)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_144),
.A2(n_142),
.B(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_111),
.C(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_101),
.Y(n_149)
);


endmodule