module fake_jpeg_6248_n_232 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_30),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_20),
.B1(n_27),
.B2(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_22),
.C(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_17),
.B1(n_27),
.B2(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_15),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_26),
.B(n_25),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_18),
.B(n_21),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_28),
.B1(n_37),
.B2(n_22),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_72),
.Y(n_76)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_28),
.B1(n_37),
.B2(n_20),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_17),
.B1(n_27),
.B2(n_24),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_65),
.B1(n_72),
.B2(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_61),
.B1(n_18),
.B2(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_36),
.B1(n_15),
.B2(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_40),
.B1(n_47),
.B2(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_26),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_70),
.C(n_21),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_32),
.A3(n_31),
.B1(n_33),
.B2(n_14),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_84),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_66),
.B1(n_23),
.B2(n_69),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_26),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_44),
.C(n_38),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_68),
.B(n_64),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_66),
.B(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_14),
.B(n_32),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_33),
.C(n_25),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_100),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_106),
.C(n_116),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_94),
.Y(n_103)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_86),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_112),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_26),
.B1(n_25),
.B2(n_31),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_88),
.B(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_80),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_92),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_132),
.C(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_83),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_114),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_138),
.B(n_109),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_83),
.A3(n_88),
.B1(n_82),
.B2(n_74),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_139),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_117),
.B(n_108),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_33),
.A3(n_39),
.B1(n_26),
.B2(n_25),
.C1(n_19),
.C2(n_63),
.Y(n_135)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_103),
.A3(n_116),
.B1(n_107),
.B2(n_110),
.C1(n_111),
.C2(n_113),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_39),
.B1(n_19),
.B2(n_33),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_140),
.B1(n_99),
.B2(n_98),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_19),
.B(n_0),
.Y(n_138)
);

NOR4xp25_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_0),
.C(n_2),
.D(n_3),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_95),
.B1(n_4),
.B2(n_5),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_147),
.C(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_121),
.B1(n_127),
.B2(n_136),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_117),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_153),
.B(n_155),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_154),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_114),
.B(n_109),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_129),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_95),
.C(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_160),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_136),
.B1(n_120),
.B2(n_126),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_167),
.B(n_122),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_164),
.Y(n_177)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_168),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_140),
.B1(n_138),
.B2(n_122),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_142),
.C(n_150),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_179),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_155),
.Y(n_179)
);

AOI21x1_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_148),
.B(n_141),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_160),
.B1(n_143),
.B2(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_143),
.C(n_158),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_170),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_166),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_133),
.B1(n_134),
.B2(n_5),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_134),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_198),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_173),
.B1(n_166),
.B2(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_200),
.B1(n_195),
.B2(n_190),
.Y(n_203)
);

AOI21x1_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_187),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_206),
.Y(n_214)
);

AO221x1_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_189),
.B1(n_165),
.B2(n_179),
.C(n_182),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_208),
.B(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_174),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_178),
.C(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_216),
.C(n_206),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_209),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_186),
.B1(n_188),
.B2(n_175),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_213),
.B(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_218),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_221),
.B1(n_6),
.B2(n_9),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_203),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_3),
.B(n_4),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_6),
.Y(n_226)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_214),
.B(n_8),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_225),
.B(n_9),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_9),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.C(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_10),
.C(n_11),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_10),
.C(n_11),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_12),
.B(n_210),
.Y(n_232)
);


endmodule