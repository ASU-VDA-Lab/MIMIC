module fake_jpeg_18680_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_35),
.B1(n_22),
.B2(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_39),
.B1(n_35),
.B2(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_85),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_71),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_84),
.B1(n_104),
.B2(n_105),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_87),
.Y(n_117)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_45),
.B1(n_50),
.B2(n_29),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_81),
.B(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_49),
.B1(n_45),
.B2(n_29),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_88),
.B1(n_93),
.B2(n_28),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_17),
.B1(n_35),
.B2(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_29),
.B1(n_46),
.B2(n_23),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_22),
.B1(n_34),
.B2(n_23),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_41),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_101),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_63),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_48),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_44),
.C(n_28),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_59),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_17),
.B1(n_25),
.B2(n_37),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_74),
.B1(n_90),
.B2(n_100),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_48),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_123),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_17),
.B1(n_37),
.B2(n_25),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_48),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_128),
.B(n_82),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_78),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_118),
.C(n_132),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_48),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_37),
.B1(n_20),
.B2(n_36),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_128),
.B1(n_114),
.B2(n_135),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_44),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_24),
.B(n_31),
.C(n_27),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_141),
.B(n_146),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_107),
.B(n_110),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_31),
.B(n_27),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_83),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_139),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_99),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_149),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_88),
.B(n_89),
.C(n_76),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_142),
.B(n_150),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_89),
.B(n_90),
.C(n_94),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_86),
.B(n_1),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_163),
.B(n_32),
.Y(n_191)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_80),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_92),
.C(n_98),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_160),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_111),
.B(n_80),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_153),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_77),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_154),
.B(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_92),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_161),
.B1(n_141),
.B2(n_138),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_109),
.A2(n_125),
.B1(n_119),
.B2(n_135),
.Y(n_159)
);

OAI22x1_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_40),
.B1(n_131),
.B2(n_18),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_77),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_128),
.B1(n_114),
.B2(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_33),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_169),
.B1(n_175),
.B2(n_184),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_0),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_106),
.B(n_20),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_181),
.B(n_187),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_130),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_168),
.A2(n_173),
.B(n_180),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_141),
.A2(n_127),
.B1(n_126),
.B2(n_125),
.Y(n_169)
);

AO21x2_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_131),
.B(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_126),
.B1(n_119),
.B2(n_120),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_186),
.B1(n_195),
.B2(n_146),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_158),
.B1(n_161),
.B2(n_144),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_120),
.B1(n_33),
.B2(n_40),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_163),
.B1(n_148),
.B2(n_153),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_179),
.B(n_185),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_19),
.B(n_33),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_145),
.B1(n_159),
.B2(n_143),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_33),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_19),
.B(n_33),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_38),
.B1(n_32),
.B2(n_26),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_32),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_191),
.B(n_192),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

XNOR2x2_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_38),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_163),
.B(n_146),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_0),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_221),
.B1(n_169),
.B2(n_180),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_162),
.C(n_149),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_224),
.C(n_227),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_204),
.Y(n_233)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_188),
.A3(n_175),
.B1(n_194),
.B2(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_210),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_171),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_207),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_163),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_208),
.A2(n_10),
.B1(n_14),
.B2(n_6),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_182),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_212),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_153),
.B1(n_148),
.B2(n_38),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_222),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_220),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_164),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

AOI32xp33_ASAP7_75t_L g223 ( 
.A1(n_167),
.A2(n_9),
.A3(n_15),
.B1(n_14),
.B2(n_6),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_172),
.B(n_181),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_9),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_196),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_9),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_226),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_8),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_229),
.A2(n_247),
.B1(n_16),
.B2(n_12),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_170),
.B(n_176),
.C(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_235),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_173),
.B1(n_165),
.B2(n_170),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_228),
.A2(n_197),
.B(n_225),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_197),
.B(n_205),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_187),
.C(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_199),
.C(n_228),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_206),
.A2(n_165),
.B1(n_170),
.B2(n_191),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_242),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_13),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_206),
.A2(n_170),
.B1(n_172),
.B2(n_5),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_198),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_203),
.B1(n_221),
.B2(n_207),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_255),
.C(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_200),
.C(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_257),
.A2(n_271),
.B(n_272),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_222),
.B1(n_214),
.B2(n_200),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_251),
.B1(n_247),
.B2(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_264),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_227),
.C(n_224),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_7),
.C(n_10),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_265),
.C(n_273),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_274),
.B1(n_244),
.B2(n_248),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_269),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_231),
.B(n_232),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_248),
.B(n_13),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_275),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_229),
.A2(n_2),
.B1(n_4),
.B2(n_13),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_253),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_278),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_253),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_285),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_232),
.B1(n_239),
.B2(n_235),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_291),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_241),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_258),
.A2(n_245),
.B(n_243),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_289),
.B(n_256),
.Y(n_306)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_258),
.B(n_272),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_307),
.B(n_308),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_267),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_299),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_266),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_292),
.B(n_289),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_271),
.C(n_263),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_282),
.C(n_286),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_293),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_316),
.Y(n_325)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_293),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_297),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_298),
.C(n_296),
.Y(n_323)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_323),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_290),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_329),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_233),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_325),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_323),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_313),
.B1(n_300),
.B2(n_281),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_310),
.B1(n_307),
.B2(n_317),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_279),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_333),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_244),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_334),
.C(n_333),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_316),
.C(n_331),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_336),
.B(n_321),
.C(n_322),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_314),
.B(n_262),
.Y(n_342)
);

A2O1A1O1Ixp25_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_283),
.B(n_230),
.C(n_337),
.D(n_260),
.Y(n_343)
);

OAI321xp33_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_244),
.A3(n_275),
.B1(n_284),
.B2(n_252),
.C(n_297),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_268),
.C(n_274),
.Y(n_345)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_319),
.B(n_311),
.Y(n_346)
);


endmodule