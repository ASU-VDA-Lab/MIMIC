module real_jpeg_11946_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_288, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_288;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_249;
wire n_83;
wire n_176;
wire n_166;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_211;
wire n_45;
wire n_160;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_258;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_20),
.B1(n_22),
.B2(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_0),
.A2(n_48),
.B1(n_55),
.B2(n_56),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_0),
.A2(n_8),
.B(n_27),
.C(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_48),
.B1(n_65),
.B2(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_0),
.B(n_25),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_0),
.B(n_63),
.C(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_0),
.B(n_54),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_0),
.B(n_28),
.C(n_30),
.Y(n_170)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_20),
.B1(n_22),
.B2(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_37),
.B1(n_65),
.B2(n_66),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_6),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_23),
.B1(n_55),
.B2(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_23),
.B1(n_65),
.B2(n_66),
.Y(n_205)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_11),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B(n_284),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_12),
.B(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_20),
.B1(n_22),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_13),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_39),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_38),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_34),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_24),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_19),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_22),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_24),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_32),
.B1(n_44),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_26),
.A2(n_36),
.B(n_76),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_26),
.A2(n_45),
.B(n_76),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

O2A1O1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_52),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_34),
.B(n_41),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_77),
.B(n_283),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_71),
.C(n_75),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_42),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.C(n_58),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_43),
.A2(n_110),
.B1(n_120),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_43),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_43),
.B(n_120),
.C(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_43),
.A2(n_86),
.B1(n_87),
.B2(n_185),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_43),
.A2(n_185),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_47),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_48),
.A2(n_52),
.B(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_48),
.B(n_106),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_48),
.B(n_69),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_49),
.A2(n_58),
.B1(n_258),
.B2(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_49),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_49)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_50),
.Y(n_260)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_56),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_58),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_58),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_58),
.B(n_173),
.C(n_259),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_59),
.A2(n_69),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_95),
.Y(n_94)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_60),
.A2(n_64),
.B1(n_93),
.B2(n_95),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_60),
.A2(n_64),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_65),
.B(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_92),
.B(n_94),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_69),
.A2(n_94),
.B(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_70),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_71),
.B(n_75),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_74),
.B1(n_88),
.B2(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_73),
.A2(n_74),
.B(n_111),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_74),
.A2(n_89),
.B(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_278),
.B(n_282),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_250),
.B(n_275),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_229),
.B(n_249),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_212),
.B(n_228),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_180),
.A3(n_207),
.B1(n_210),
.B2(n_211),
.C(n_288),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_162),
.B(n_179),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_128),
.B(n_161),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_107),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_85),
.B(n_107),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.C(n_96),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_145),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_86),
.A2(n_87),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_87),
.B(n_172),
.C(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_87),
.B(n_185),
.C(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_91),
.A2(n_132),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_91),
.A2(n_145),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_95),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_96),
.A2(n_97),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_102),
.B(n_205),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_105),
.A2(n_106),
.B1(n_188),
.B2(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_106),
.A2(n_118),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_122),
.B2(n_123),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_125),
.C(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_120),
.B2(n_121),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_113),
.C(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_120),
.A2(n_244),
.B(n_247),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_120),
.B(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_127),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_137),
.C(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_125),
.A2(n_127),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_125),
.B(n_204),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_155),
.B(n_160),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_141),
.B(n_154),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_139),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_168),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_146),
.B(n_153),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_187),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B(n_152),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_167),
.C(n_171),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_173),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_195),
.C(n_200),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_172),
.A2(n_173),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_172),
.A2(n_173),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_173),
.B(n_269),
.C(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_191),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_190),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_182),
.B(n_186),
.CI(n_190),
.CON(n_209),
.SN(n_209)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_206),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_201),
.B2(n_202),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_202),
.C(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_209),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_227),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_227),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_216),
.C(n_221),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_224),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_222),
.A2(n_226),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_235),
.B(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_231),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_248),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_242),
.B2(n_243),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_242),
.C(n_248),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_254),
.B1(n_255),
.B2(n_262),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_247),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_265),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_264),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_264),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_262),
.C(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_259),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_274),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_274),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_273),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_281),
.Y(n_282)
);


endmodule