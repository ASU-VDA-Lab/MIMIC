module fake_jpeg_6711_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_44),
.B(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_19),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_52),
.B1(n_65),
.B2(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_31),
.B1(n_19),
.B2(n_30),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_34),
.Y(n_55)
);

OR2x4_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_18),
.B1(n_27),
.B2(n_34),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_29),
.B(n_28),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_27),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_33),
.B(n_38),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_72),
.B(n_51),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_33),
.B(n_38),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_82),
.B1(n_32),
.B2(n_21),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_39),
.B1(n_20),
.B2(n_24),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_77),
.B1(n_85),
.B2(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_39),
.B1(n_43),
.B2(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_86),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_24),
.B1(n_39),
.B2(n_23),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_38),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_67),
.B(n_38),
.C(n_36),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_59),
.B1(n_55),
.B2(n_63),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_44),
.A2(n_39),
.B1(n_25),
.B2(n_43),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_98),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_51),
.C(n_65),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_83),
.Y(n_125)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_103),
.B(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_43),
.B(n_38),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_108),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_36),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_72),
.B1(n_80),
.B2(n_91),
.Y(n_140)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_69),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_28),
.Y(n_165)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_128),
.B(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_84),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_135),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_83),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_0),
.B(n_32),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_142),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_149),
.B1(n_91),
.B2(n_102),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_77),
.B1(n_84),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_114),
.B1(n_109),
.B2(n_97),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_79),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_145),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_75),
.B(n_80),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_114),
.B(n_89),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_154),
.B(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_172),
.B1(n_175),
.B2(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_165),
.Y(n_185)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_169),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_111),
.C(n_108),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_168),
.C(n_177),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_118),
.B(n_116),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_45),
.B(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_173),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_134),
.A2(n_45),
.B(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_178),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_176),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_0),
.B(n_21),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_91),
.B1(n_45),
.B2(n_66),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_81),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_21),
.A3(n_66),
.B1(n_64),
.B2(n_0),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_182),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_139),
.B(n_133),
.C(n_143),
.D(n_144),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_157),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_132),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_177),
.C(n_163),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_127),
.B1(n_122),
.B2(n_140),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_193),
.A2(n_194),
.B1(n_200),
.B2(n_168),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_147),
.B1(n_141),
.B2(n_123),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_199),
.Y(n_223)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_146),
.B1(n_126),
.B2(n_145),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_188),
.B1(n_137),
.B2(n_102),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_154),
.B(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_151),
.B(n_128),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_214),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_167),
.C(n_166),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_221),
.C(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_225),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_178),
.B1(n_153),
.B2(n_179),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_218),
.B1(n_224),
.B2(n_226),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_158),
.B1(n_155),
.B2(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_203),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_165),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_175),
.C(n_81),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_190),
.A2(n_1),
.B(n_2),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_64),
.B1(n_81),
.B2(n_73),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_73),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_228),
.A2(n_184),
.B1(n_181),
.B2(n_202),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_73),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_200),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_232),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_235),
.C(n_239),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_184),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_244),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_237),
.B(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_206),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_216),
.B1(n_218),
.B2(n_221),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_198),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_247),
.C(n_248),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_183),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_5),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_195),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_224),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_210),
.B(n_187),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_113),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_208),
.B1(n_213),
.B2(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_261),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_228),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_262),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_258),
.B(n_259),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_229),
.B(n_220),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_2),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_64),
.B1(n_113),
.B2(n_7),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_264),
.C(n_268),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_230),
.C(n_248),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_256),
.A2(n_230),
.B1(n_6),
.B2(n_8),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_270),
.A2(n_260),
.B1(n_249),
.B2(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_5),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_272),
.B(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_16),
.C(n_6),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_5),
.C(n_8),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_9),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_277),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_282),
.B(n_268),
.C(n_13),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_262),
.B(n_10),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_278),
.A2(n_274),
.B(n_12),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_12),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_9),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_11),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_278),
.B(n_279),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_282),
.Y(n_294)
);

OAI21x1_ASAP7_75t_SL g295 ( 
.A1(n_288),
.A2(n_290),
.B(n_291),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_284),
.B1(n_15),
.B2(n_14),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_13),
.B(n_14),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_281),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_288),
.B(n_295),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_297),
.C(n_293),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_281),
.C(n_296),
.Y(n_301)
);


endmodule