module real_jpeg_10341_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_325, n_11, n_14, n_7, n_3, n_5, n_4, n_324, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_325;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_324;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_1),
.A2(n_23),
.B1(n_61),
.B2(n_62),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_1),
.A2(n_23),
.B1(n_46),
.B2(n_47),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_46),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_3),
.B(n_46),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_3),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_3),
.A2(n_32),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_3),
.B(n_32),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_3),
.B(n_36),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_29),
.B(n_33),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_107),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_4),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_141),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_141),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_141),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_5),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_56),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_8),
.A2(n_46),
.B(n_59),
.C(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_11),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_82),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_82),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_82),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_12),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_123),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_123),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_123),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_13),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_94),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_94),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_15),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_54),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_16),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_16),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_17),
.A2(n_61),
.B1(n_62),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_17),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_17),
.A2(n_46),
.B1(n_47),
.B2(n_87),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_87),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_87),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_316),
.B(n_319),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_69),
.B(n_315),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_21),
.B(n_37),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_21),
.B(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_21),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_22),
.A2(n_26),
.B1(n_36),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_24),
.A2(n_28),
.B(n_107),
.C(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_26),
.A2(n_36),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_26),
.A2(n_34),
.B(n_36),
.Y(n_318)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_27),
.A2(n_31),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_27),
.A2(n_31),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_27),
.A2(n_31),
.B1(n_211),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_27),
.A2(n_31),
.B1(n_229),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_27),
.A2(n_31),
.B1(n_246),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_27),
.A2(n_31),
.B1(n_53),
.B2(n_267),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_65),
.C(n_67),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_38),
.A2(n_39),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_51),
.C(n_57),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_40),
.A2(n_41),
.B1(n_57),
.B2(n_293),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_45),
.B(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_42),
.A2(n_45),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_42),
.A2(n_45),
.B1(n_132),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_42),
.A2(n_45),
.B1(n_149),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_42),
.A2(n_45),
.B1(n_189),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_42),
.A2(n_45),
.B1(n_207),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_42),
.A2(n_45),
.B1(n_226),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_42),
.A2(n_45),
.B1(n_243),
.B2(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_42),
.A2(n_45),
.B1(n_49),
.B2(n_260),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_44),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_45),
.B(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_46),
.B(n_48),
.Y(n_136)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_47),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_51),
.A2(n_52),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_57),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_57),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_60),
.B(n_64),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_60),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_60),
.B1(n_93),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_58),
.A2(n_60),
.B1(n_120),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_58),
.A2(n_60),
.B1(n_128),
.B2(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_58),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_58),
.A2(n_60),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_58),
.A2(n_60),
.B1(n_202),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_58),
.A2(n_60),
.B1(n_221),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_58),
.A2(n_60),
.B1(n_64),
.B2(n_252),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_60),
.B(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_60),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_61),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_61),
.B(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_65),
.A2(n_67),
.B1(n_68),
.B2(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_65),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_308),
.B(n_314),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_285),
.A3(n_303),
.B1(n_306),
.B2(n_307),
.C(n_324),
.Y(n_70)
);

AOI321xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_236),
.A3(n_273),
.B1(n_279),
.B2(n_284),
.C(n_325),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_194),
.C(n_233),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_164),
.B(n_193),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_143),
.B(n_163),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_125),
.B(n_142),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_114),
.B(n_124),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_100),
.B(n_113),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_88),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_83),
.A2(n_84),
.B1(n_140),
.B2(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_104),
.B1(n_105),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_99),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_99),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_108),
.B(n_112),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_106),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_105),
.B1(n_122),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_104),
.A2(n_105),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_104),
.A2(n_105),
.B1(n_175),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_104),
.A2(n_105),
.B1(n_199),
.B2(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_104),
.A2(n_105),
.B(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_107),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_126),
.Y(n_142)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.CI(n_121),
.CON(n_117),
.SN(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.CI(n_133),
.CON(n_126),
.SN(n_126)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_145),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_156),
.B2(n_157),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_159),
.C(n_161),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_155),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_166),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_179),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_178),
.C(n_179),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_173),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_190),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_187),
.B2(n_188),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_187),
.C(n_190),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_195),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_214),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_196),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_196),
.B(n_214),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_203),
.CI(n_204),
.CON(n_196),
.SN(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_200),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_213),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_212),
.C(n_213),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_231),
.B2(n_232),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_217),
.B(n_222),
.C(n_232),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_220),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_227),
.C(n_230),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_231),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_235),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_255),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_237),
.B(n_255),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_248),
.C(n_254),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_239),
.B1(n_248),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_244),
.C(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_242),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_248),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_250),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_249),
.A2(n_266),
.B(n_269),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_251),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_251),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_271),
.B2(n_272),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_263),
.C(n_272),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_261),
.B(n_262),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_287),
.C(n_295),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_262),
.B(n_287),
.CI(n_295),
.CON(n_305),
.SN(n_305)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_269),
.B2(n_270),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_271),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_280),
.B(n_283),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_296),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_296),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_289),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_293),
.C(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_298),
.C(n_302),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_313),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_310),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);


endmodule