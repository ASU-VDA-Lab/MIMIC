module fake_jpeg_4199_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_17),
.B1(n_21),
.B2(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_14),
.B1(n_22),
.B2(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_34),
.B1(n_20),
.B2(n_17),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_14),
.B1(n_17),
.B2(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_17),
.B1(n_15),
.B2(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_43),
.Y(n_44)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_20),
.B1(n_38),
.B2(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_18),
.Y(n_68)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_15),
.B(n_18),
.C(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_57),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_20),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_35),
.B(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_43),
.B1(n_33),
.B2(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_62),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_64),
.B1(n_72),
.B2(n_33),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_68),
.B1(n_55),
.B2(n_54),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_28),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_53),
.B1(n_57),
.B2(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_37),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_28),
.B(n_12),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

AOI32xp33_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_40),
.A3(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_77),
.B1(n_80),
.B2(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_55),
.B1(n_48),
.B2(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_83),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_54),
.B1(n_20),
.B2(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_58),
.B(n_70),
.Y(n_87)
);

AOI321xp33_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_92),
.A3(n_40),
.B1(n_37),
.B2(n_16),
.C(n_71),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_72),
.B(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_89),
.B1(n_85),
.B2(n_84),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_69),
.B(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_96),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_69),
.B(n_40),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_40),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_92),
.C(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_74),
.B1(n_86),
.B2(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_114),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_87),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_110),
.C(n_99),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_79),
.B1(n_78),
.B2(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_19),
.B1(n_22),
.B2(n_18),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_75),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_40),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_71),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_114),
.B(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_97),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_123),
.C(n_130),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_99),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_120),
.B(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_37),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_127),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_40),
.C(n_37),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_33),
.B1(n_18),
.B2(n_12),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_19),
.B1(n_16),
.B2(n_7),
.Y(n_139)
);

NOR4xp25_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_8),
.C(n_11),
.D(n_10),
.Y(n_128)
);

OAI322xp33_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_124),
.A3(n_118),
.B1(n_19),
.B2(n_130),
.C1(n_10),
.C2(n_9),
.Y(n_134)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_56),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_0),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_R g152 ( 
.A(n_134),
.B(n_8),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_101),
.C(n_29),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_9),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_8),
.B1(n_7),
.B2(n_2),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_149),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_29),
.B1(n_16),
.B2(n_2),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_151),
.B1(n_153),
.B2(n_136),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_16),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_136),
.B1(n_142),
.B2(n_139),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_1),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_140),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_163),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_140),
.C(n_132),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_161),
.B(n_4),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_3),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_149),
.B1(n_152),
.B2(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_2),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_13),
.C(n_3),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_13),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_166),
.B(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_3),
.Y(n_166)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_158),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_157),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_4),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_4),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_164),
.C(n_6),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_173),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_156),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_176),
.C(n_5),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_6),
.C(n_13),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_5),
.C(n_6),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_5),
.B(n_6),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_13),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_184),
.B(n_13),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_13),
.B(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_182),
.Y(n_186)
);


endmodule