module fake_jpeg_5493_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_13),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_43),
.Y(n_72)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_0),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_15),
.B(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_52),
.Y(n_80)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_53),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_23),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_46),
.B1(n_47),
.B2(n_59),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_90),
.B1(n_109),
.B2(n_31),
.Y(n_117)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_76),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_33),
.B1(n_32),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_82),
.B1(n_87),
.B2(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_79),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_83),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_33),
.B1(n_37),
.B2(n_28),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_39),
.A2(n_33),
.B1(n_37),
.B2(n_23),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_22),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_17),
.B1(n_27),
.B2(n_18),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_28),
.B1(n_21),
.B2(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_16),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_26),
.B1(n_21),
.B2(n_24),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_108),
.B1(n_9),
.B2(n_2),
.Y(n_135)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_45),
.A2(n_28),
.B1(n_26),
.B2(n_17),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_105),
.B1(n_106),
.B2(n_29),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_44),
.B(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_36),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_48),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_48),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_52),
.A2(n_15),
.B1(n_22),
.B2(n_25),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_112),
.Y(n_164)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_116),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_118),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_139),
.B1(n_64),
.B2(n_87),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_125),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_84),
.B1(n_81),
.B2(n_107),
.Y(n_158)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_25),
.A3(n_22),
.B1(n_11),
.B2(n_10),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_80),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_63),
.A2(n_9),
.B1(n_22),
.B2(n_3),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_130),
.B(n_84),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_138),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_130),
.B1(n_139),
.B2(n_126),
.Y(n_162)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_73),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_89),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_63),
.Y(n_157)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_64),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_147),
.Y(n_187)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_158),
.B1(n_162),
.B2(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_151),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_67),
.B1(n_123),
.B2(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_92),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_179),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_118),
.B(n_75),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_169),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_137),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_161),
.B(n_171),
.Y(n_216)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_170),
.Y(n_193)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_70),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_130),
.B(n_1),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_93),
.C(n_83),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_110),
.B(n_121),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_9),
.Y(n_202)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_178),
.B1(n_153),
.B2(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_78),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_183),
.Y(n_243)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_185),
.B(n_206),
.CI(n_209),
.CON(n_220),
.SN(n_220)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_186),
.B(n_189),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_170),
.A2(n_62),
.B1(n_71),
.B2(n_104),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_192),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_67),
.B1(n_136),
.B2(n_98),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_200),
.B1(n_66),
.B2(n_3),
.Y(n_239)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_162),
.A2(n_99),
.B1(n_62),
.B2(n_120),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_204),
.B1(n_159),
.B2(n_123),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_211),
.B(n_213),
.Y(n_223)
);

AOI22x1_ASAP7_75t_L g204 ( 
.A1(n_157),
.A2(n_116),
.B1(n_114),
.B2(n_96),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_208),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_116),
.B(n_131),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_207),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_154),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_111),
.B(n_113),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_1),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_156),
.Y(n_217)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_156),
.B(n_163),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_241),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_222),
.B1(n_229),
.B2(n_240),
.Y(n_247)
);

NAND2x1_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_216),
.Y(n_224)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_210),
.B(n_192),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_150),
.B1(n_148),
.B2(n_171),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_166),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_202),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_180),
.A2(n_178),
.B(n_155),
.Y(n_229)
);

OAI32xp33_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_145),
.A3(n_151),
.B1(n_149),
.B2(n_165),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_232),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_166),
.A3(n_147),
.B1(n_176),
.B2(n_96),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_147),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_237),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_120),
.B1(n_141),
.B2(n_167),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_131),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_112),
.B1(n_153),
.B2(n_66),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_2),
.B(n_3),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_194),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_204),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_4),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_185),
.C(n_198),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_248),
.C(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_250),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_251),
.B(n_254),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_214),
.B(n_195),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_213),
.C(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_263),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_233),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_193),
.C(n_196),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_262),
.C(n_237),
.Y(n_286)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_188),
.C(n_183),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

BUFx12_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_217),
.Y(n_285)
);

NOR4xp25_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_232),
.C(n_218),
.D(n_205),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_229),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_277),
.B(n_283),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_268),
.B1(n_255),
.B2(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_272),
.B(n_281),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_268),
.A2(n_222),
.B1(n_227),
.B2(n_243),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_276),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_247),
.A2(n_227),
.B1(n_244),
.B2(n_225),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_220),
.B1(n_241),
.B2(n_230),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_230),
.B1(n_186),
.B2(n_219),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_240),
.B(n_189),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_253),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_245),
.C(n_246),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_293),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_249),
.B(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_296),
.C(n_278),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_256),
.A3(n_260),
.B1(n_262),
.B2(n_265),
.C1(n_248),
.C2(n_258),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_281),
.Y(n_304)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_234),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_257),
.C(n_263),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_187),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_182),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_236),
.B(n_264),
.C(n_212),
.D(n_197),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_285),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_276),
.B1(n_277),
.B2(n_270),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_306),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_300),
.A2(n_270),
.B1(n_269),
.B2(n_283),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_273),
.B1(n_282),
.B2(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_308),
.C(n_310),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_298),
.B1(n_289),
.B2(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_297),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_264),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_299),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_274),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_314),
.A2(n_315),
.B(n_316),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_293),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_296),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_199),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_321),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_278),
.C(n_284),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_309),
.B(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_311),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_323),
.B1(n_326),
.B2(n_190),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_306),
.B1(n_208),
.B2(n_236),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_SL g328 ( 
.A(n_325),
.B(n_321),
.C(n_319),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_312),
.B(n_182),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_330),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_203),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_332),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_324),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_331),
.Y(n_337)
);


endmodule