module fake_netlist_6_2792_n_1755 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1755);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1755;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_5),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_33),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_11),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_69),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_108),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_89),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_51),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_23),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_68),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_26),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_95),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_20),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_10),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_75),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_26),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_56),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_41),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_71),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_4),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_101),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_10),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_2),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_54),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_28),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_84),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_78),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_0),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_140),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_70),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_111),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_29),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_2),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_7),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_40),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_13),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_93),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_53),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_98),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_62),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_29),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_42),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_81),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_64),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_83),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_16),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_38),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_43),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_67),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_66),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_11),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_138),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_19),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_30),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_141),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_58),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_43),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_25),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_41),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_63),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_46),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_35),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_74),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_22),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_90),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_19),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_17),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_54),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_1),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_119),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_143),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_96),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_79),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_61),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_4),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_14),
.Y(n_254)
);

BUFx8_ASAP7_75t_SL g255 ( 
.A(n_44),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_80),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_132),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_120),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_82),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_59),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_33),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_100),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_5),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_12),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_18),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_55),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_105),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_38),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_32),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_52),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_123),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_109),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_94),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_135),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_113),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_60),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_107),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_103),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_104),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_27),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_99),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_73),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_121),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_65),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_7),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_55),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_36),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_3),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_106),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_22),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_50),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_118),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_51),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_53),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_32),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_1),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_77),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_13),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_102),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_91),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_125),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_17),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_217),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_169),
.B(n_0),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_255),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_217),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_173),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_216),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_161),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_162),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_237),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_217),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_168),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_221),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_257),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_171),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_175),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_285),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_169),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_217),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_176),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_306),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_178),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_180),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_6),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_159),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_159),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_182),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_157),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_184),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_288),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_194),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_184),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_196),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_181),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_181),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_272),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_187),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_198),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_210),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_166),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_166),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_199),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_183),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_200),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_185),
.B(n_6),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_206),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_210),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_183),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_185),
.B(n_8),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_226),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_207),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_214),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_215),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_191),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_191),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_271),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_220),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_223),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_271),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_227),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_192),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_232),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_238),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_179),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_192),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_310),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_380),
.A2(n_187),
.B(n_179),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_353),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_363),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_275),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_380),
.A2(n_187),
.B(n_251),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_190),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

AND3x2_ASAP7_75t_L g402 ( 
.A(n_311),
.B(n_225),
.C(n_251),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_190),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_275),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_336),
.B(n_224),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_335),
.B(n_296),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_314),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_349),
.B(n_296),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_359),
.B(n_302),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_280),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_280),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_315),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_370),
.A2(n_212),
.B(n_208),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_371),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_324),
.Y(n_434)
);

AND2x2_ASAP7_75t_SL g435 ( 
.A(n_361),
.B(n_302),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_155),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_343),
.B(n_361),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_366),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_375),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_155),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_328),
.B(n_160),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_381),
.B(n_156),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_350),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_156),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_435),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_385),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_431),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_396),
.B(n_317),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_386),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_445),
.B(n_343),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_445),
.B(n_318),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_386),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_385),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_437),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_391),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_391),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_398),
.B(n_165),
.Y(n_469)
);

BUFx6f_ASAP7_75t_SL g470 ( 
.A(n_435),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_398),
.B(n_165),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_401),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_345),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

CKINVDCx6p67_ASAP7_75t_R g476 ( 
.A(n_411),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_321),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_431),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

AND3x2_ASAP7_75t_L g483 ( 
.A(n_392),
.B(n_337),
.C(n_330),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_431),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_408),
.B(n_325),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_435),
.A2(n_319),
.B1(n_301),
.B2(n_292),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

INVx11_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_435),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_409),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_407),
.Y(n_492)
);

BUFx6f_ASAP7_75t_SL g493 ( 
.A(n_435),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_398),
.B(n_186),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_386),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_386),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_351),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_326),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_438),
.B(n_331),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_437),
.B(n_333),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_434),
.B(n_339),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_398),
.B(n_334),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_434),
.B(n_341),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_398),
.B(n_346),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_447),
.A2(n_236),
.B1(n_188),
.B2(n_170),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_386),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_382),
.Y(n_511)
);

BUFx4f_ASAP7_75t_L g512 ( 
.A(n_436),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_382),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g514 ( 
.A(n_443),
.B(n_193),
.C(n_186),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_443),
.B(n_197),
.C(n_193),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_382),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_389),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_389),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_398),
.B(n_404),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_384),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_404),
.B(n_348),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_411),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_386),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_386),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_399),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_447),
.B(n_354),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_387),
.B(n_339),
.C(n_284),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_402),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_399),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_386),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_402),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_403),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_387),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_412),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_429),
.B(n_358),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_429),
.B(n_360),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_384),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_403),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_403),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_415),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_429),
.B(n_197),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_430),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_394),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_429),
.B(n_362),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_413),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_429),
.B(n_367),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_415),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_415),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_429),
.B(n_374),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_413),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_R g556 ( 
.A(n_387),
.B(n_393),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_443),
.A2(n_240),
.B1(n_189),
.B2(n_208),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_404),
.B(n_379),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_443),
.B(n_211),
.C(n_209),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_415),
.Y(n_560)
);

INVx11_ASAP7_75t_L g561 ( 
.A(n_410),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_413),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_394),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_394),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_394),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_428),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_443),
.B(n_368),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_418),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_384),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_384),
.Y(n_572)
);

AND3x2_ASAP7_75t_L g573 ( 
.A(n_440),
.B(n_211),
.C(n_209),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_383),
.B(n_164),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_443),
.A2(n_240),
.B1(n_189),
.B2(n_308),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_428),
.B(n_312),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_394),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_418),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_418),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_428),
.B(n_228),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_446),
.B(n_369),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_414),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_414),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_L g584 ( 
.A(n_428),
.B(n_239),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_446),
.B(n_228),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_446),
.B(n_378),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_446),
.A2(n_201),
.B1(n_299),
.B2(n_307),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_414),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_394),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_436),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_446),
.B(n_234),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_393),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_446),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_393),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_582),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_521),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_590),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_590),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_436),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_450),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_449),
.B(n_394),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_568),
.B(n_436),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_449),
.B(n_394),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_479),
.B(n_373),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_485),
.B(n_405),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_527),
.B(n_436),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_488),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_490),
.B(n_394),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_490),
.B(n_456),
.Y(n_609)
);

OAI221xp5_ASAP7_75t_L g610 ( 
.A1(n_557),
.A2(n_252),
.B1(n_219),
.B2(n_212),
.C(n_254),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_495),
.B(n_436),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_489),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_583),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_495),
.B(n_436),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_495),
.B(n_293),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_474),
.B(n_383),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_474),
.B(n_383),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_470),
.A2(n_252),
.B1(n_219),
.B2(n_254),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_522),
.B(n_383),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_470),
.A2(n_376),
.B1(n_323),
.B2(n_327),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_450),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_488),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_454),
.A2(n_283),
.B(n_290),
.C(n_291),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_491),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_521),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_491),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_558),
.B(n_158),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_593),
.B(n_383),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_L g630 ( 
.A(n_501),
.B(n_405),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_502),
.B(n_163),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_593),
.B(n_390),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_529),
.B(n_440),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_521),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_500),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_580),
.B(n_390),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_470),
.A2(n_322),
.B1(n_332),
.B2(n_247),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_512),
.B(n_293),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_458),
.B(n_167),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_451),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_451),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_486),
.B(n_174),
.C(n_172),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_500),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_594),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_580),
.B(n_390),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_571),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_452),
.B(n_395),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_571),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_454),
.B(n_390),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_448),
.A2(n_294),
.B1(n_291),
.B2(n_297),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_486),
.B(n_195),
.C(n_177),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_461),
.B(n_390),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_512),
.B(n_520),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_461),
.B(n_390),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_462),
.B(n_426),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_503),
.B(n_203),
.C(n_202),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_493),
.A2(n_256),
.B1(n_241),
.B2(n_248),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_494),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_462),
.B(n_426),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_468),
.B(n_426),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_493),
.A2(n_294),
.B1(n_297),
.B2(n_290),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_494),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_468),
.B(n_426),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_477),
.B(n_426),
.Y(n_665)
);

INVxp33_ASAP7_75t_L g666 ( 
.A(n_464),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_477),
.B(n_426),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_452),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_476),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_588),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_480),
.B(n_444),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_498),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_512),
.B(n_293),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_480),
.B(n_484),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_484),
.B(n_293),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_493),
.A2(n_448),
.B1(n_581),
.B2(n_569),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_498),
.B(n_444),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_504),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_511),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_588),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_448),
.A2(n_250),
.B1(n_235),
.B2(n_253),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_591),
.B(n_293),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_511),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_540),
.B(n_444),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_513),
.Y(n_685)
);

NOR2xp67_ASAP7_75t_L g686 ( 
.A(n_592),
.B(n_405),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_513),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_585),
.A2(n_587),
.B(n_551),
.C(n_591),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_516),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_585),
.B(n_444),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_516),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_505),
.B(n_293),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_591),
.B(n_444),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_504),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_591),
.B(n_444),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_469),
.B(n_293),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_574),
.B(n_469),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_576),
.B(n_420),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_448),
.A2(n_235),
.B1(n_234),
.B2(n_250),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_448),
.A2(n_283),
.B1(n_308),
.B2(n_258),
.Y(n_700)
);

AND2x6_ASAP7_75t_SL g701 ( 
.A(n_476),
.B(n_253),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_L g702 ( 
.A1(n_509),
.A2(n_258),
.B1(n_274),
.B2(n_304),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_469),
.B(n_419),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_455),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_469),
.B(n_293),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_472),
.B(n_293),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_489),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_455),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_472),
.B(n_541),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_517),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_518),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_459),
.B(n_204),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_508),
.A2(n_287),
.B1(n_274),
.B2(n_278),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_529),
.B(n_205),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_556),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_576),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_463),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_535),
.B(n_249),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_472),
.B(n_400),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_472),
.B(n_572),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_587),
.A2(n_278),
.B1(n_282),
.B2(n_287),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_525),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_571),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_518),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_525),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_535),
.B(n_400),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_519),
.B(n_419),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_519),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_526),
.B(n_419),
.Y(n_729)
);

INVxp33_ASAP7_75t_L g730 ( 
.A(n_537),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_526),
.B(n_419),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_530),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_530),
.B(n_419),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_523),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_463),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_523),
.B(n_440),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_586),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_531),
.B(n_419),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_531),
.B(n_282),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_536),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_525),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_536),
.B(n_304),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_543),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_543),
.B(n_424),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_544),
.B(n_424),
.Y(n_745)
);

BUFx8_ASAP7_75t_L g746 ( 
.A(n_547),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_509),
.B(n_395),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_544),
.B(n_424),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_528),
.B(n_395),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_525),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_550),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_546),
.Y(n_752)
);

INVx5_ASAP7_75t_L g753 ( 
.A(n_525),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_584),
.A2(n_263),
.B1(n_267),
.B2(n_270),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_550),
.B(n_422),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_555),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_555),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_539),
.B(n_213),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_549),
.A2(n_397),
.B(n_388),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_554),
.B(n_218),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_SL g761 ( 
.A(n_575),
.B(n_222),
.Y(n_761)
);

INVxp67_ASAP7_75t_SL g762 ( 
.A(n_532),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_514),
.A2(n_388),
.B1(n_397),
.B2(n_224),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_674),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_662),
.B(n_547),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_609),
.B(n_563),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_635),
.B(n_430),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_573),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_499),
.B(n_457),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_741),
.Y(n_770)
);

NOR2x1_ASAP7_75t_L g771 ( 
.A(n_605),
.B(n_514),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_722),
.A2(n_499),
.B(n_457),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_631),
.B(n_563),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_722),
.A2(n_499),
.B(n_457),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_643),
.B(n_647),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_722),
.A2(n_499),
.B(n_457),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_710),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_700),
.A2(n_546),
.B(n_515),
.C(n_559),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_630),
.B(n_546),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_712),
.A2(n_515),
.B(n_559),
.C(n_397),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_700),
.A2(n_546),
.B(n_579),
.C(n_578),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_759),
.A2(n_397),
.B(n_388),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_734),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_722),
.A2(n_548),
.B(n_532),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_741),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_753),
.A2(n_548),
.B(n_532),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_698),
.B(n_532),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_644),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_712),
.A2(n_388),
.B(n_589),
.C(n_460),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_628),
.B(n_597),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_753),
.A2(n_548),
.B(n_532),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_740),
.Y(n_792)
);

O2A1O1Ixp5_ASAP7_75t_L g793 ( 
.A1(n_638),
.A2(n_510),
.B(n_460),
.C(n_497),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_668),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_740),
.Y(n_795)
);

AO21x1_ASAP7_75t_L g796 ( 
.A1(n_616),
.A2(n_553),
.B(n_552),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_678),
.B(n_546),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_628),
.B(n_460),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_753),
.A2(n_548),
.B(n_453),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_753),
.A2(n_453),
.B(n_524),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_598),
.B(n_497),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_599),
.B(n_497),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_744),
.B(n_589),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_715),
.B(n_483),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_653),
.A2(n_453),
.B(n_524),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_745),
.B(n_510),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_611),
.A2(n_561),
.B1(n_577),
.B2(n_567),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_694),
.B(n_510),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_604),
.B(n_564),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_748),
.B(n_589),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_596),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_653),
.A2(n_453),
.B(n_524),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_621),
.B(n_276),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_730),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_686),
.B(n_224),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_606),
.A2(n_453),
.B(n_524),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_614),
.A2(n_453),
.B(n_524),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_679),
.B(n_564),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_614),
.A2(n_524),
.B(n_534),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_762),
.A2(n_534),
.B(n_562),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_617),
.A2(n_534),
.B(n_562),
.Y(n_821)
);

OAI21xp33_ASAP7_75t_L g822 ( 
.A1(n_639),
.A2(n_229),
.B(n_262),
.Y(n_822)
);

INVx11_ASAP7_75t_L g823 ( 
.A(n_746),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_716),
.B(n_420),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_675),
.A2(n_564),
.B(n_565),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_618),
.A2(n_534),
.B(n_562),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_709),
.A2(n_534),
.B(n_562),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_666),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_720),
.A2(n_534),
.B(n_562),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_620),
.A2(n_562),
.B(n_565),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_683),
.B(n_565),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_639),
.A2(n_567),
.B(n_577),
.C(n_578),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_746),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_685),
.B(n_567),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_751),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_741),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_636),
.A2(n_570),
.B(n_566),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_633),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_645),
.A2(n_570),
.B(n_566),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_687),
.B(n_465),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_688),
.A2(n_467),
.B(n_560),
.C(n_553),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_604),
.B(n_224),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_688),
.A2(n_561),
.B1(n_277),
.B2(n_279),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_689),
.B(n_465),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_599),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_691),
.B(n_466),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_711),
.B(n_466),
.Y(n_847)
);

INVx5_ASAP7_75t_L g848 ( 
.A(n_741),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_702),
.B(n_676),
.C(n_651),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_723),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_612),
.B(n_707),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_684),
.A2(n_560),
.B(n_552),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_642),
.B(n_714),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_624),
.A2(n_545),
.B(n_542),
.C(n_538),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_602),
.A2(n_545),
.B(n_542),
.Y(n_855)
);

NOR2x1_ASAP7_75t_L g856 ( 
.A(n_656),
.B(n_467),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_675),
.A2(n_603),
.B(n_601),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_649),
.A2(n_538),
.B(n_533),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_724),
.B(n_728),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_758),
.A2(n_533),
.B(n_507),
.C(n_496),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_652),
.A2(n_507),
.B(n_496),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_596),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_654),
.A2(n_492),
.B(n_487),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_714),
.B(n_230),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_601),
.A2(n_492),
.B(n_487),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_732),
.B(n_743),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_690),
.B(n_471),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_756),
.B(n_471),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_757),
.B(n_634),
.Y(n_869)
);

AOI21xp33_ASAP7_75t_L g870 ( 
.A1(n_758),
.A2(n_231),
.B(n_242),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_736),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_603),
.A2(n_482),
.B(n_481),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_608),
.A2(n_482),
.B(n_481),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_608),
.A2(n_478),
.B(n_475),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_SL g875 ( 
.A(n_669),
.B(n_298),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_616),
.A2(n_298),
.B1(n_478),
.B2(n_473),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_634),
.A2(n_475),
.B(n_473),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_607),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_747),
.B(n_233),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_693),
.B(n_400),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_646),
.B(n_281),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_760),
.B(n_298),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_657),
.B(n_286),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_646),
.B(n_305),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_760),
.B(n_243),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_655),
.A2(n_660),
.B(n_659),
.Y(n_886)
);

NAND2x1_ASAP7_75t_L g887 ( 
.A(n_612),
.B(n_400),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_619),
.B(n_420),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_664),
.A2(n_417),
.B(n_410),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_637),
.B(n_427),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_623),
.B(n_422),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_619),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_625),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_627),
.B(n_422),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_665),
.A2(n_400),
.B(n_425),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_633),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_595),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_658),
.B(n_422),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_667),
.A2(n_671),
.B(n_632),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_629),
.A2(n_400),
.B(n_423),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_613),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_661),
.B(n_427),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_663),
.B(n_423),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_726),
.B(n_749),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_726),
.B(n_265),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_672),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_723),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_661),
.B(n_423),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_752),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_626),
.B(n_423),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_633),
.B(n_298),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_626),
.B(n_425),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_626),
.B(n_648),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_613),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_626),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_615),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_702),
.B(n_721),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_752),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_719),
.A2(n_400),
.B(n_425),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_695),
.A2(n_703),
.B(n_677),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_648),
.B(n_425),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_761),
.A2(n_442),
.B(n_441),
.C(n_439),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_719),
.A2(n_400),
.B(n_406),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_638),
.A2(n_400),
.B(n_406),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_648),
.B(n_615),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_624),
.A2(n_442),
.B(n_441),
.C(n_439),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_673),
.A2(n_400),
.B(n_406),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_673),
.A2(n_416),
.B(n_406),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_650),
.A2(n_442),
.B(n_441),
.C(n_439),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_727),
.A2(n_410),
.B(n_417),
.Y(n_930)
);

OAI21xp33_ASAP7_75t_L g931 ( 
.A1(n_737),
.A2(n_309),
.B(n_289),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_648),
.A2(n_273),
.B1(n_295),
.B2(n_300),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_681),
.A2(n_433),
.B(n_427),
.C(n_303),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_682),
.B(n_433),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_692),
.A2(n_416),
.B(n_406),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_650),
.A2(n_433),
.B(n_9),
.C(n_12),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_699),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_729),
.A2(n_417),
.B(n_410),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_725),
.A2(n_416),
.B(n_406),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_718),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_701),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_670),
.B(n_432),
.Y(n_942)
);

BUFx12f_ASAP7_75t_L g943 ( 
.A(n_783),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_764),
.A2(n_755),
.B(n_738),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_764),
.A2(n_707),
.B1(n_725),
.B2(n_750),
.Y(n_945)
);

AOI22x1_ASAP7_75t_L g946 ( 
.A1(n_882),
.A2(n_670),
.B1(n_680),
.B2(n_640),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_792),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_798),
.A2(n_731),
.B(n_733),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_885),
.A2(n_713),
.B(n_739),
.C(n_742),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_790),
.A2(n_682),
.B(n_680),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_789),
.A2(n_696),
.B(n_705),
.Y(n_951)
);

NOR2xp67_ASAP7_75t_R g952 ( 
.A(n_896),
.B(n_750),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_795),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_886),
.A2(n_899),
.B(n_766),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_833),
.Y(n_955)
);

XNOR2x2_ASAP7_75t_SL g956 ( 
.A(n_842),
.B(n_754),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_920),
.A2(n_705),
.B(n_696),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_767),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_885),
.A2(n_706),
.B(n_610),
.C(n_717),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_904),
.B(n_600),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_864),
.A2(n_706),
.B(n_735),
.C(n_708),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_848),
.A2(n_806),
.B(n_803),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_848),
.A2(n_704),
.B(n_641),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_918),
.B(n_622),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_848),
.A2(n_763),
.B(n_416),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_853),
.A2(n_763),
.B1(n_432),
.B2(n_421),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_853),
.B(n_432),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_814),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_904),
.A2(n_421),
.B1(n_432),
.B2(n_416),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_823),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_810),
.A2(n_416),
.B(n_406),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_864),
.B(n_432),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_SL g973 ( 
.A(n_804),
.B(n_8),
.C(n_14),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_775),
.B(n_768),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_879),
.B(n_15),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_777),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_768),
.B(n_432),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_809),
.A2(n_421),
.B1(n_432),
.B2(n_416),
.Y(n_978)
);

OAI22x1_ASAP7_75t_L g979 ( 
.A1(n_917),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_811),
.B(n_86),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_913),
.A2(n_416),
.B(n_406),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_788),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_862),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_917),
.A2(n_432),
.B(n_421),
.C(n_416),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_809),
.B(n_432),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_870),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_782),
.A2(n_406),
.B(n_421),
.Y(n_987)
);

INVx6_ASAP7_75t_L g988 ( 
.A(n_862),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_940),
.A2(n_432),
.B1(n_421),
.B2(n_76),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_879),
.A2(n_21),
.B(n_24),
.C(n_25),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_SL g991 ( 
.A(n_849),
.B(n_822),
.C(n_875),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_828),
.B(n_421),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_835),
.Y(n_993)
);

OAI22xp33_ASAP7_75t_L g994 ( 
.A1(n_871),
.A2(n_421),
.B1(n_30),
.B2(n_31),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_781),
.A2(n_421),
.B(n_417),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_918),
.B(n_88),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_SL g997 ( 
.A1(n_941),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_878),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_769),
.A2(n_421),
.B(n_92),
.Y(n_999)
);

INVx8_ASAP7_75t_L g1000 ( 
.A(n_770),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_794),
.B(n_34),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_772),
.A2(n_776),
.B(n_774),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_940),
.B(n_97),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_845),
.B(n_87),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_849),
.A2(n_845),
.B1(n_905),
.B2(n_937),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_937),
.A2(n_37),
.B(n_39),
.C(n_42),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_794),
.B(n_37),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_788),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_893),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_862),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_773),
.A2(n_417),
.B(n_410),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_857),
.A2(n_417),
.B(n_410),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_862),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_SL g1014 ( 
.A1(n_780),
.A2(n_115),
.B(n_151),
.C(n_150),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_905),
.B(n_417),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_906),
.B(n_417),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_910),
.A2(n_417),
.B(n_410),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_770),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_765),
.B(n_39),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_838),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_914),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_804),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_912),
.A2(n_417),
.B(n_410),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_921),
.A2(n_417),
.B(n_410),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_859),
.B(n_417),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_797),
.B(n_57),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_915),
.B(n_110),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_779),
.A2(n_410),
.B(n_148),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_866),
.B(n_410),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_815),
.B(n_45),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_909),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_925),
.A2(n_137),
.B(n_130),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_869),
.A2(n_867),
.B(n_841),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_SL g1034 ( 
.A1(n_832),
.A2(n_144),
.B(n_128),
.C(n_47),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_936),
.A2(n_933),
.B(n_931),
.C(n_922),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_932),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_867),
.A2(n_45),
.B(n_46),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_850),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_SL g1039 ( 
.A(n_770),
.B(n_48),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_SL g1040 ( 
.A(n_892),
.B(n_49),
.C(n_50),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_793),
.A2(n_52),
.B(n_860),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_897),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_911),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_808),
.B(n_850),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_824),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_901),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_907),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_907),
.B(n_808),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_890),
.B(n_811),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_915),
.B(n_883),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_813),
.B(n_888),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_916),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_902),
.A2(n_929),
.B(n_843),
.C(n_778),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_908),
.A2(n_926),
.B(n_868),
.C(n_846),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_915),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_915),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_881),
.B(n_884),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_934),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_856),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_840),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_784),
.A2(n_791),
.B(n_786),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_934),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_796),
.A2(n_787),
.B(n_816),
.C(n_852),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_SL g1064 ( 
.A(n_771),
.B(n_770),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_807),
.A2(n_880),
.B(n_855),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_802),
.B(n_880),
.C(n_938),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_876),
.B(n_847),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_785),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_802),
.A2(n_934),
.B1(n_876),
.B2(n_844),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_785),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_818),
.B(n_831),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_834),
.B(n_801),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_891),
.B(n_903),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_825),
.A2(n_889),
.B(n_930),
.C(n_894),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_898),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_785),
.B(n_836),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_785),
.B(n_836),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_SL g1078 ( 
.A(n_854),
.B(n_851),
.C(n_837),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_942),
.Y(n_1079)
);

AO32x2_ASAP7_75t_L g1080 ( 
.A1(n_966),
.A2(n_1038),
.A3(n_945),
.B1(n_1062),
.B2(n_989),
.Y(n_1080)
);

OA21x2_ASAP7_75t_L g1081 ( 
.A1(n_984),
.A2(n_839),
.B(n_863),
.Y(n_1081)
);

OR2x6_ASAP7_75t_L g1082 ( 
.A(n_1000),
.B(n_836),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_1000),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_982),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_968),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1005),
.A2(n_836),
.B1(n_851),
.B2(n_817),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_998),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_L g1088 ( 
.A(n_975),
.B(n_900),
.C(n_919),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_958),
.B(n_865),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1049),
.B(n_874),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1000),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_991),
.A2(n_873),
.B1(n_872),
.B2(n_895),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_990),
.A2(n_858),
.B(n_861),
.C(n_877),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_943),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_954),
.A2(n_830),
.B(n_799),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_1010),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_974),
.A2(n_928),
.B(n_935),
.C(n_927),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_986),
.A2(n_924),
.B(n_923),
.C(n_827),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1065),
.A2(n_805),
.A3(n_812),
.B(n_829),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_954),
.A2(n_819),
.B(n_887),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1019),
.A2(n_939),
.B(n_821),
.C(n_826),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1002),
.A2(n_820),
.B(n_800),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1057),
.A2(n_972),
.B(n_944),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_957),
.A2(n_949),
.B(n_1067),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_944),
.A2(n_957),
.B(n_1061),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_1018),
.B(n_1008),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1009),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1021),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1078),
.A2(n_948),
.B(n_1073),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1047),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_959),
.A2(n_1069),
.B(n_951),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_948),
.A2(n_1072),
.B(n_1071),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1036),
.A2(n_1031),
.B1(n_1030),
.B2(n_979),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1049),
.B(n_1004),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_951),
.A2(n_1053),
.B(n_1035),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1054),
.A2(n_1051),
.B(n_961),
.C(n_950),
.Y(n_1116)
);

NAND3xp33_ASAP7_75t_L g1117 ( 
.A(n_1040),
.B(n_973),
.C(n_1006),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_950),
.A2(n_1033),
.B(n_1066),
.C(n_1059),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1018),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_1020),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1063),
.A2(n_971),
.B(n_1033),
.Y(n_1121)
);

BUFx2_ASAP7_75t_SL g1122 ( 
.A(n_1018),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_985),
.A2(n_1065),
.B(n_962),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1045),
.B(n_1022),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1041),
.A2(n_1037),
.B(n_1060),
.C(n_1048),
.Y(n_1125)
);

OA21x2_ASAP7_75t_L g1126 ( 
.A1(n_987),
.A2(n_995),
.B(n_967),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_960),
.A2(n_977),
.B(n_1015),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_994),
.A2(n_1001),
.B1(n_1007),
.B2(n_1058),
.Y(n_1128)
);

CKINVDCx8_ASAP7_75t_R g1129 ( 
.A(n_970),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_971),
.A2(n_987),
.B(n_981),
.Y(n_1130)
);

AOI211x1_ASAP7_75t_L g1131 ( 
.A1(n_1037),
.A2(n_1044),
.B(n_947),
.C(n_953),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1074),
.A2(n_965),
.B(n_999),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1018),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_992),
.Y(n_1134)
);

CKINVDCx6p67_ASAP7_75t_R g1135 ( 
.A(n_955),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_946),
.A2(n_956),
.B(n_1079),
.Y(n_1136)
);

OA21x2_ASAP7_75t_L g1137 ( 
.A1(n_995),
.A2(n_1028),
.B(n_1032),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_1028),
.A2(n_1032),
.B(n_1012),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1075),
.B(n_964),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1042),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_963),
.A2(n_978),
.B(n_969),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1043),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1017),
.A2(n_1023),
.B(n_1024),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_SL g1144 ( 
.A(n_1055),
.B(n_1068),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1064),
.A2(n_1050),
.B(n_1014),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_964),
.B(n_1004),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_996),
.B(n_993),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1025),
.A2(n_1029),
.B(n_976),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_996),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1011),
.A2(n_1016),
.A3(n_1052),
.B(n_1046),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1026),
.A2(n_1039),
.B1(n_997),
.B2(n_1070),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1011),
.A2(n_1024),
.A3(n_1023),
.B(n_1017),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_983),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1076),
.A2(n_1077),
.B(n_1034),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_952),
.A2(n_1026),
.B(n_983),
.Y(n_1155)
);

INVxp67_ASAP7_75t_SL g1156 ( 
.A(n_1013),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1026),
.B(n_1013),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1027),
.A2(n_1056),
.B1(n_988),
.B2(n_980),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1056),
.A2(n_1027),
.B(n_988),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_SL g1161 ( 
.A1(n_984),
.A2(n_688),
.B(n_1003),
.C(n_975),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1005),
.B(n_662),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_975),
.A2(n_885),
.B(n_631),
.C(n_864),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_998),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_968),
.B(n_1018),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_975),
.B(n_631),
.C(n_885),
.Y(n_1170)
);

BUFx2_ASAP7_75t_R g1171 ( 
.A(n_970),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_975),
.A2(n_853),
.B(n_885),
.C(n_631),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_975),
.A2(n_631),
.B1(n_885),
.B2(n_849),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1005),
.B(n_662),
.Y(n_1174)
);

INVxp67_ASAP7_75t_L g1175 ( 
.A(n_982),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1005),
.B(n_662),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_975),
.A2(n_885),
.B1(n_631),
.B2(n_917),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_975),
.B(n_715),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_998),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_968),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1005),
.B(n_662),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_998),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_975),
.A2(n_853),
.B(n_885),
.C(n_631),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1005),
.B(n_662),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_958),
.B(n_775),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_975),
.B(n_715),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_998),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_968),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_998),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_968),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1005),
.B(n_662),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_SL g1197 ( 
.A1(n_984),
.A2(n_688),
.B(n_1003),
.C(n_975),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_968),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_SL g1200 ( 
.A(n_975),
.B(n_470),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_SL g1201 ( 
.A1(n_975),
.A2(n_885),
.B(n_631),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1005),
.B(n_662),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1049),
.B(n_918),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_SL g1206 ( 
.A1(n_975),
.A2(n_700),
.B1(n_702),
.B2(n_917),
.C(n_650),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_982),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_958),
.B(n_775),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_975),
.B(n_631),
.C(n_885),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_975),
.A2(n_885),
.B(n_631),
.C(n_864),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_954),
.A2(n_764),
.B(n_1057),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_975),
.A2(n_917),
.B1(n_509),
.B2(n_885),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1002),
.A2(n_1061),
.B(n_1063),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_975),
.A2(n_885),
.B(n_631),
.C(n_864),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_998),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_SL g1217 ( 
.A1(n_1037),
.A2(n_1041),
.B(n_1035),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_975),
.B(n_662),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1005),
.A2(n_631),
.B1(n_609),
.B2(n_764),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1124),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1192),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_1085),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1194),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1170),
.A2(n_1210),
.B1(n_1173),
.B2(n_1177),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1201),
.A2(n_1177),
.B(n_1163),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1083),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1119),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1170),
.A2(n_1210),
.B1(n_1200),
.B2(n_1218),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1213),
.A2(n_1117),
.B1(n_1115),
.B2(n_1219),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1129),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1162),
.B(n_1174),
.Y(n_1231)
);

OAI22xp33_ASAP7_75t_R g1232 ( 
.A1(n_1207),
.A2(n_1084),
.B1(n_1182),
.B2(n_1094),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_SL g1233 ( 
.A1(n_1200),
.A2(n_1111),
.B1(n_1202),
.B2(n_1195),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1199),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1176),
.A2(n_1183),
.B1(n_1186),
.B2(n_1117),
.Y(n_1235)
);

OAI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1201),
.A2(n_1128),
.B1(n_1113),
.B2(n_1139),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_1135),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1113),
.A2(n_1217),
.B1(n_1128),
.B2(n_1189),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1171),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1087),
.Y(n_1240)
);

BUFx12f_ASAP7_75t_L g1241 ( 
.A(n_1120),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1178),
.A2(n_1104),
.B1(n_1151),
.B2(n_1112),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1119),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1134),
.A2(n_1146),
.B1(n_1089),
.B2(n_1147),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1107),
.Y(n_1245)
);

INVxp67_ASAP7_75t_SL g1246 ( 
.A(n_1160),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1211),
.A2(n_1215),
.B(n_1185),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1133),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1172),
.A2(n_1114),
.B1(n_1149),
.B2(n_1142),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1165),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1133),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1110),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1181),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1114),
.A2(n_1188),
.B1(n_1208),
.B2(n_1090),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1133),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1207),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1175),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1083),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1205),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1190),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1205),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1193),
.Y(n_1262)
);

INVx6_ASAP7_75t_L g1263 ( 
.A(n_1083),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1091),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1091),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1091),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1136),
.A2(n_1140),
.B1(n_1216),
.B2(n_1108),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1134),
.B(n_1157),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1166),
.A2(n_1196),
.B1(n_1203),
.B2(n_1212),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1169),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1082),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1158),
.A2(n_1206),
.B1(n_1179),
.B2(n_1187),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1082),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1106),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1158),
.A2(n_1125),
.B1(n_1191),
.B2(n_1118),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1116),
.A2(n_1103),
.B1(n_1155),
.B2(n_1145),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1153),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1082),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1206),
.A2(n_1088),
.B1(n_1086),
.B2(n_1122),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1096),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1127),
.A2(n_1088),
.B1(n_1109),
.B2(n_1148),
.Y(n_1281)
);

CKINVDCx6p67_ASAP7_75t_R g1282 ( 
.A(n_1144),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1137),
.A2(n_1138),
.B1(n_1126),
.B2(n_1154),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1137),
.A2(n_1138),
.B1(n_1126),
.B2(n_1132),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1105),
.A2(n_1156),
.B1(n_1143),
.B2(n_1123),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1096),
.A2(n_1081),
.B1(n_1092),
.B2(n_1159),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1161),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1092),
.A2(n_1081),
.B1(n_1197),
.B2(n_1121),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1131),
.B(n_1150),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1152),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1141),
.A2(n_1080),
.B1(n_1214),
.B2(n_1168),
.Y(n_1291)
);

BUFx4f_ASAP7_75t_L g1292 ( 
.A(n_1131),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1097),
.Y(n_1293)
);

INVx3_ASAP7_75t_SL g1294 ( 
.A(n_1080),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1080),
.A2(n_1209),
.B1(n_1164),
.B2(n_1204),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1167),
.A2(n_1198),
.B1(n_1180),
.B2(n_1130),
.Y(n_1296)
);

OAI21xp33_ASAP7_75t_L g1297 ( 
.A1(n_1098),
.A2(n_1101),
.B(n_1093),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1100),
.B(n_1095),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1099),
.Y(n_1299)
);

INVx6_ASAP7_75t_L g1300 ( 
.A(n_1102),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1177),
.A2(n_1173),
.B1(n_1210),
.B2(n_1170),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1213),
.A2(n_1210),
.B1(n_1170),
.B2(n_1173),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1188),
.B(n_1208),
.Y(n_1303)
);

BUFx4f_ASAP7_75t_SL g1304 ( 
.A(n_1135),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1177),
.A2(n_1173),
.B1(n_1210),
.B2(n_1170),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1188),
.B(n_1208),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1218),
.B(n_1162),
.Y(n_1307)
);

CKINVDCx11_ASAP7_75t_R g1308 ( 
.A(n_1129),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1184),
.Y(n_1309)
);

INVx6_ASAP7_75t_L g1310 ( 
.A(n_1083),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1085),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1188),
.B(n_1208),
.Y(n_1312)
);

OAI21xp33_ASAP7_75t_L g1313 ( 
.A1(n_1177),
.A2(n_1173),
.B(n_885),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1184),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1085),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_1119),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1213),
.A2(n_1210),
.B1(n_1170),
.B2(n_1173),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1213),
.A2(n_1210),
.B1(n_1170),
.B2(n_1173),
.Y(n_1318)
);

CKINVDCx6p67_ASAP7_75t_R g1319 ( 
.A(n_1192),
.Y(n_1319)
);

INVx6_ASAP7_75t_L g1320 ( 
.A(n_1083),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1213),
.A2(n_1210),
.B1(n_1170),
.B2(n_1173),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1170),
.A2(n_1210),
.B1(n_975),
.B2(n_1200),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1218),
.B(n_1162),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1085),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1170),
.A2(n_1210),
.B1(n_1173),
.B2(n_1177),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1184),
.Y(n_1326)
);

BUFx2_ASAP7_75t_SL g1327 ( 
.A(n_1192),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1192),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1201),
.A2(n_1177),
.B1(n_1210),
.B2(n_1170),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1177),
.A2(n_1173),
.B1(n_1210),
.B2(n_1170),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1129),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1119),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1213),
.A2(n_1210),
.B1(n_1170),
.B2(n_1173),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1184),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1129),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1129),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1129),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1170),
.A2(n_1210),
.B1(n_975),
.B2(n_1200),
.Y(n_1338)
);

BUFx4_ASAP7_75t_SL g1339 ( 
.A(n_1192),
.Y(n_1339)
);

BUFx12f_ASAP7_75t_L g1340 ( 
.A(n_1085),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1290),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1268),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1289),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1299),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1292),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1292),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1313),
.A2(n_1247),
.B(n_1301),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1293),
.Y(n_1348)
);

BUFx4f_ASAP7_75t_SL g1349 ( 
.A(n_1230),
.Y(n_1349)
);

AND2x2_ASAP7_75t_SL g1350 ( 
.A(n_1224),
.B(n_1325),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1246),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1287),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1246),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1240),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1294),
.B(n_1329),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1245),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1252),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1286),
.B(n_1253),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1250),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1298),
.B(n_1249),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1307),
.B(n_1323),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1300),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1262),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1294),
.Y(n_1364)
);

OAI211xp5_ASAP7_75t_L g1365 ( 
.A1(n_1302),
.A2(n_1318),
.B(n_1317),
.C(n_1333),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1297),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1229),
.B(n_1302),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1300),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1231),
.B(n_1235),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1275),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1260),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1276),
.A2(n_1269),
.B(n_1284),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1273),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1277),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1272),
.A2(n_1225),
.B(n_1305),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1309),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1272),
.A2(n_1330),
.B(n_1236),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1314),
.Y(n_1378)
);

OAI21xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1229),
.A2(n_1317),
.B(n_1318),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1236),
.A2(n_1238),
.B1(n_1228),
.B2(n_1333),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1326),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1334),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1321),
.B(n_1233),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1271),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1273),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1295),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1295),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1220),
.B(n_1257),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1269),
.A2(n_1283),
.B(n_1285),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1244),
.A2(n_1296),
.B(n_1291),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1321),
.B(n_1233),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1220),
.B(n_1303),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1288),
.A2(n_1281),
.B(n_1267),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1235),
.B(n_1244),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1306),
.B(n_1312),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1267),
.B(n_1242),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1291),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1288),
.A2(n_1281),
.B(n_1242),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1273),
.Y(n_1399)
);

INVxp67_ASAP7_75t_L g1400 ( 
.A(n_1324),
.Y(n_1400)
);

INVxp67_ASAP7_75t_R g1401 ( 
.A(n_1339),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1271),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1279),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1279),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1238),
.A2(n_1296),
.B(n_1254),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1228),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1322),
.A2(n_1338),
.B(n_1232),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1322),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1338),
.A2(n_1256),
.B1(n_1278),
.B2(n_1259),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1280),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1261),
.B(n_1223),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1270),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1222),
.A2(n_1340),
.B1(n_1315),
.B2(n_1311),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1316),
.B(n_1255),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1227),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1248),
.B(n_1255),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1380),
.A2(n_1274),
.B(n_1327),
.C(n_1332),
.Y(n_1417)
);

NOR4xp25_ASAP7_75t_SL g1418 ( 
.A(n_1366),
.B(n_1239),
.C(n_1264),
.D(n_1234),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1282),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1342),
.B(n_1221),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1342),
.B(n_1265),
.Y(n_1421)
);

AOI211xp5_ASAP7_75t_L g1422 ( 
.A1(n_1347),
.A2(n_1409),
.B(n_1365),
.C(n_1379),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1349),
.Y(n_1423)
);

OAI21xp33_ASAP7_75t_L g1424 ( 
.A1(n_1347),
.A2(n_1328),
.B(n_1237),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1380),
.A2(n_1251),
.B(n_1255),
.C(n_1332),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1355),
.B(n_1332),
.Y(n_1426)
);

AND2x2_ASAP7_75t_SL g1427 ( 
.A(n_1350),
.B(n_1243),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1351),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1395),
.B(n_1251),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1379),
.A2(n_1337),
.B(n_1336),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1361),
.B(n_1319),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1369),
.B(n_1251),
.Y(n_1432)
);

OAI21xp33_ASAP7_75t_L g1433 ( 
.A1(n_1350),
.A2(n_1255),
.B(n_1335),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1373),
.B(n_1258),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1350),
.A2(n_1304),
.B1(n_1241),
.B2(n_1263),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1392),
.B(n_1226),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1398),
.A2(n_1226),
.B(n_1263),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_SL g1438 ( 
.A1(n_1365),
.A2(n_1266),
.B(n_1308),
.C(n_1331),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1406),
.B(n_1383),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1406),
.B(n_1310),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1394),
.A2(n_1310),
.B(n_1320),
.C(n_1383),
.Y(n_1441)
);

AND2x6_ASAP7_75t_L g1442 ( 
.A(n_1345),
.B(n_1310),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1391),
.B(n_1320),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1394),
.A2(n_1346),
.B1(n_1345),
.B2(n_1352),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1398),
.A2(n_1372),
.B(n_1389),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1391),
.B(n_1408),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1367),
.B(n_1366),
.C(n_1408),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1364),
.B(n_1354),
.Y(n_1448)
);

AOI211xp5_ASAP7_75t_L g1449 ( 
.A1(n_1370),
.A2(n_1346),
.B(n_1396),
.C(n_1403),
.Y(n_1449)
);

INVxp33_ASAP7_75t_L g1450 ( 
.A(n_1411),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1407),
.A2(n_1377),
.B1(n_1375),
.B2(n_1396),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1376),
.B(n_1378),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1381),
.B(n_1410),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1407),
.B(n_1370),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1352),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1351),
.A2(n_1353),
.B(n_1377),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1362),
.B(n_1368),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_SL g1458 ( 
.A(n_1407),
.B(n_1375),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1364),
.B(n_1356),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1407),
.B(n_1403),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1410),
.B(n_1414),
.Y(n_1461)
);

AOI211xp5_ASAP7_75t_L g1462 ( 
.A1(n_1404),
.A2(n_1388),
.B(n_1400),
.C(n_1352),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1414),
.B(n_1375),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1359),
.Y(n_1464)
);

AND2x2_ASAP7_75t_SL g1465 ( 
.A(n_1393),
.B(n_1353),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1389),
.A2(n_1405),
.B(n_1387),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1362),
.B(n_1368),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1352),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1360),
.B(n_1358),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1377),
.A2(n_1404),
.B1(n_1360),
.B2(n_1352),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1374),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_SL g1472 ( 
.A(n_1352),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1377),
.B(n_1348),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1401),
.A2(n_1413),
.B1(n_1412),
.B2(n_1357),
.Y(n_1474)
);

AO32x1_ASAP7_75t_L g1475 ( 
.A1(n_1386),
.A2(n_1387),
.A3(n_1397),
.B1(n_1348),
.B2(n_1341),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1402),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1471),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1471),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1428),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1454),
.B(n_1343),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1466),
.B(n_1448),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1466),
.B(n_1397),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1424),
.A2(n_1393),
.B1(n_1358),
.B2(n_1390),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1465),
.B(n_1390),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1464),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1442),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1465),
.B(n_1390),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1466),
.B(n_1463),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1475),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1475),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1475),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1428),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1445),
.B(n_1390),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1459),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1433),
.A2(n_1393),
.B1(n_1358),
.B2(n_1371),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1445),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1419),
.B(n_1363),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1473),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1452),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1475),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1453),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1447),
.A2(n_1393),
.B1(n_1358),
.B2(n_1382),
.Y(n_1502)
);

INVx5_ASAP7_75t_L g1503 ( 
.A(n_1469),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1437),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1473),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1457),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1467),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1454),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1460),
.B(n_1451),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1486),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1503),
.B(n_1467),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1508),
.B(n_1498),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1503),
.B(n_1469),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1492),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1492),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1478),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1497),
.B(n_1460),
.Y(n_1517)
);

NAND4xp25_ASAP7_75t_L g1518 ( 
.A(n_1509),
.B(n_1422),
.C(n_1449),
.D(n_1462),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1496),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1508),
.B(n_1456),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1509),
.B(n_1470),
.C(n_1419),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1507),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1494),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1461),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1482),
.B(n_1432),
.Y(n_1525)
);

AND2x4_ASAP7_75t_SL g1526 ( 
.A(n_1494),
.B(n_1469),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1482),
.B(n_1344),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1504),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1482),
.B(n_1344),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1506),
.B(n_1458),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1479),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1497),
.B(n_1446),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1477),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1477),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1484),
.A2(n_1427),
.B1(n_1444),
.B2(n_1474),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1499),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1483),
.A2(n_1427),
.B1(n_1468),
.B2(n_1455),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1479),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1426),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1485),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1485),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1484),
.A2(n_1435),
.B1(n_1430),
.B2(n_1439),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1485),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1520),
.B(n_1505),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1541),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1540),
.B(n_1484),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1540),
.B(n_1487),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1525),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1511),
.B(n_1487),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1510),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1541),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1542),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1512),
.B(n_1505),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1542),
.Y(n_1555)
);

AOI33xp33_ASAP7_75t_L g1556 ( 
.A1(n_1535),
.A2(n_1487),
.A3(n_1483),
.B1(n_1493),
.B2(n_1502),
.B3(n_1488),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1511),
.B(n_1488),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1450),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1511),
.B(n_1488),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1518),
.B(n_1486),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1525),
.B(n_1481),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1516),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1512),
.B(n_1481),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1522),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1516),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1544),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1521),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1523),
.B(n_1481),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1511),
.B(n_1506),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1510),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1516),
.Y(n_1572)
);

AND2x2_ASAP7_75t_SL g1573 ( 
.A(n_1543),
.B(n_1502),
.Y(n_1573)
);

NAND2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1510),
.B(n_1503),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1544),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1533),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1527),
.B(n_1480),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1527),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1533),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1534),
.Y(n_1580)
);

INVx4_ASAP7_75t_L g1581 ( 
.A(n_1510),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1530),
.B(n_1506),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1522),
.B(n_1493),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1568),
.A2(n_1521),
.B1(n_1537),
.B2(n_1513),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1554),
.B(n_1549),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1513),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1568),
.B(n_1532),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1546),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1550),
.B(n_1536),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1550),
.B(n_1513),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1549),
.B(n_1529),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1567),
.B(n_1499),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1513),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1567),
.B(n_1524),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1546),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1551),
.B(n_1526),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1551),
.B(n_1503),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1552),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1545),
.B(n_1529),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1552),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1553),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1573),
.A2(n_1537),
.B1(n_1503),
.B2(n_1438),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1554),
.B(n_1524),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1562),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1553),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1564),
.B(n_1526),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1555),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1564),
.B(n_1526),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1555),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1571),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1566),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1562),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1566),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1575),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1545),
.B(n_1501),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1558),
.B(n_1450),
.Y(n_1616)
);

NAND2x1p5_ASAP7_75t_L g1617 ( 
.A(n_1581),
.B(n_1503),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1575),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1576),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1562),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1564),
.B(n_1514),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1565),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1576),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1563),
.B(n_1501),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1573),
.A2(n_1493),
.B(n_1441),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1588),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1606),
.B(n_1571),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1596),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1595),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1606),
.B(n_1557),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1598),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1610),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1608),
.B(n_1557),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1608),
.B(n_1590),
.Y(n_1635)
);

OAI321xp33_ASAP7_75t_L g1636 ( 
.A1(n_1584),
.A2(n_1574),
.A3(n_1558),
.B1(n_1563),
.B2(n_1556),
.C(n_1573),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1604),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1585),
.B(n_1569),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1596),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1600),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1625),
.A2(n_1438),
.B1(n_1578),
.B2(n_1581),
.C(n_1583),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1596),
.B(n_1586),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1601),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1599),
.B(n_1577),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1616),
.B(n_1560),
.Y(n_1646)
);

OAI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1616),
.A2(n_1560),
.B(n_1441),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1587),
.B(n_1423),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1605),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1594),
.B(n_1547),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1590),
.B(n_1559),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1589),
.B(n_1559),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1589),
.B(n_1581),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1586),
.B(n_1581),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1548),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_SL g1657 ( 
.A(n_1597),
.B(n_1472),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1607),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1621),
.B(n_1548),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1615),
.B(n_1577),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1632),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1639),
.B(n_1628),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1599),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1632),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1647),
.B(n_1591),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1646),
.A2(n_1468),
.B1(n_1455),
.B2(n_1586),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1647),
.B(n_1591),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1642),
.A2(n_1602),
.B1(n_1593),
.B2(n_1574),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_SL g1669 ( 
.A1(n_1648),
.A2(n_1472),
.B1(n_1636),
.B2(n_1423),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1626),
.A2(n_1593),
.B1(n_1623),
.B2(n_1619),
.C(n_1609),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1657),
.A2(n_1617),
.B(n_1597),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1627),
.B(n_1593),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1657),
.A2(n_1617),
.B1(n_1574),
.B2(n_1611),
.C(n_1618),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1643),
.A2(n_1434),
.B(n_1495),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1638),
.B(n_1624),
.Y(n_1676)
);

AOI211xp5_ASAP7_75t_L g1677 ( 
.A1(n_1655),
.A2(n_1401),
.B(n_1417),
.C(n_1434),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1627),
.B(n_1635),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1643),
.A2(n_1635),
.B(n_1654),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1626),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1629),
.A2(n_1613),
.B1(n_1614),
.B2(n_1620),
.C(n_1622),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1629),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1631),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1643),
.B(n_1431),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1630),
.B(n_1578),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1666),
.B(n_1643),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1661),
.B(n_1633),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1669),
.A2(n_1633),
.B1(n_1654),
.B2(n_1417),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1670),
.A2(n_1665),
.B1(n_1667),
.B2(n_1664),
.C(n_1662),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1674),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1678),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1679),
.A2(n_1655),
.B1(n_1630),
.B2(n_1634),
.Y(n_1692)
);

NAND4xp25_ASAP7_75t_L g1693 ( 
.A(n_1668),
.B(n_1631),
.C(n_1658),
.D(n_1644),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1685),
.B(n_1634),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1661),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1675),
.A2(n_1671),
.B1(n_1677),
.B2(n_1673),
.C(n_1672),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1674),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1685),
.B(n_1651),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1663),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1680),
.B(n_1640),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1684),
.B(n_1651),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1682),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1683),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_1638),
.Y(n_1704)
);

O2A1O1Ixp5_ASAP7_75t_L g1705 ( 
.A1(n_1688),
.A2(n_1686),
.B(n_1687),
.C(n_1699),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1689),
.A2(n_1693),
.B1(n_1695),
.B2(n_1696),
.C(n_1691),
.Y(n_1706)
);

NOR3x1_ASAP7_75t_L g1707 ( 
.A(n_1687),
.B(n_1688),
.C(n_1700),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1704),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1690),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1697),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1700),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1702),
.B(n_1681),
.Y(n_1712)
);

OAI31xp33_ASAP7_75t_L g1713 ( 
.A1(n_1694),
.A2(n_1684),
.A3(n_1640),
.B(n_1658),
.Y(n_1713)
);

AOI211x1_ASAP7_75t_L g1714 ( 
.A1(n_1701),
.A2(n_1644),
.B(n_1649),
.C(n_1656),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1698),
.B(n_1650),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1692),
.A2(n_1703),
.B(n_1649),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_L g1717 ( 
.A(n_1706),
.B(n_1641),
.C(n_1637),
.Y(n_1717)
);

NOR4xp25_ASAP7_75t_SL g1718 ( 
.A(n_1710),
.B(n_1531),
.C(n_1579),
.D(n_1580),
.Y(n_1718)
);

NOR3x1_ASAP7_75t_L g1719 ( 
.A(n_1708),
.B(n_1641),
.C(n_1659),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1705),
.A2(n_1637),
.B(n_1653),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1645),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_L g1722 ( 
.A(n_1712),
.B(n_1637),
.C(n_1660),
.Y(n_1722)
);

NOR2xp67_ASAP7_75t_SL g1723 ( 
.A(n_1711),
.B(n_1645),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1709),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1713),
.B(n_1652),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1712),
.B(n_1652),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1723),
.B(n_1716),
.Y(n_1727)
);

AOI211x1_ASAP7_75t_SL g1728 ( 
.A1(n_1720),
.A2(n_1707),
.B(n_1714),
.C(n_1604),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1717),
.A2(n_1622),
.B1(n_1620),
.B2(n_1612),
.C(n_1583),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1724),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1725),
.B(n_1726),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1730),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1727),
.A2(n_1722),
.B1(n_1721),
.B2(n_1719),
.C(n_1718),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_R g1734 ( 
.A(n_1731),
.B(n_1420),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1729),
.A2(n_1561),
.B1(n_1612),
.B2(n_1425),
.C(n_1583),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1728),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1727),
.A2(n_1539),
.B1(n_1514),
.B2(n_1515),
.C(n_1580),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1732),
.B(n_1579),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1734),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1736),
.Y(n_1740)
);

NAND4xp75_ASAP7_75t_L g1741 ( 
.A(n_1733),
.B(n_1539),
.C(n_1436),
.D(n_1515),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1735),
.Y(n_1742)
);

OAI321xp33_ASAP7_75t_L g1743 ( 
.A1(n_1740),
.A2(n_1737),
.A3(n_1561),
.B1(n_1443),
.B2(n_1440),
.C(n_1416),
.Y(n_1743)
);

AND4x1_ASAP7_75t_L g1744 ( 
.A(n_1739),
.B(n_1425),
.C(n_1418),
.D(n_1421),
.Y(n_1744)
);

OAI321xp33_ASAP7_75t_L g1745 ( 
.A1(n_1742),
.A2(n_1416),
.A3(n_1500),
.B1(n_1489),
.B2(n_1491),
.C(n_1490),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1743),
.Y(n_1746)
);

AO22x2_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1741),
.B1(n_1738),
.B2(n_1744),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_SL g1748 ( 
.A1(n_1747),
.A2(n_1745),
.B(n_1565),
.Y(n_1748)
);

AOI22x1_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1572),
.B1(n_1565),
.B2(n_1476),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1749),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1572),
.B1(n_1570),
.B2(n_1582),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1429),
.B(n_1415),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1752),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1528),
.B1(n_1538),
.B2(n_1519),
.Y(n_1754)
);

AOI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1385),
.B(n_1399),
.C(n_1384),
.Y(n_1755)
);


endmodule