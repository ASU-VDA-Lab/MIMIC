module fake_jpeg_29115_n_274 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_274);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_14),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_62),
.Y(n_80)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_9),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_69),
.Y(n_88)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_11),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_25),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_24),
.B1(n_20),
.B2(n_28),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_100),
.B1(n_81),
.B2(n_74),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_24),
.B1(n_22),
.B2(n_39),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_20),
.B1(n_69),
.B2(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_41),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_41),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_101),
.Y(n_143)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_111),
.B1(n_119),
.B2(n_128),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_109),
.Y(n_145)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_107),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_20),
.B(n_29),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_72),
.B1(n_67),
.B2(n_61),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_120),
.B1(n_127),
.B2(n_129),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_57),
.B1(n_64),
.B2(n_47),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_116),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_54),
.C(n_39),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_123),
.CI(n_43),
.CON(n_137),
.SN(n_137)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_49),
.B1(n_50),
.B2(n_28),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_124),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_34),
.B(n_31),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_89),
.B(n_85),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

AO22x2_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_42),
.B1(n_38),
.B2(n_27),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_26),
.B1(n_42),
.B2(n_38),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_27),
.B1(n_50),
.B2(n_3),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_77),
.B1(n_26),
.B2(n_28),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_119),
.B1(n_136),
.B2(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_128),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_117),
.B(n_115),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_166),
.B(n_15),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_144),
.B(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_131),
.B1(n_141),
.B2(n_135),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_128),
.B1(n_114),
.B2(n_112),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_134),
.B1(n_141),
.B2(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_111),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_163),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_124),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_164),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_144),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_17),
.B(n_18),
.C(n_16),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_174),
.B1(n_160),
.B2(n_132),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_162),
.B1(n_151),
.B2(n_159),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_116),
.B1(n_113),
.B2(n_102),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_184),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_147),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_196),
.B1(n_200),
.B2(n_174),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_150),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_180),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_197),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_151),
.B1(n_161),
.B2(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_166),
.B1(n_132),
.B2(n_142),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_147),
.B(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_146),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_183),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_132),
.B1(n_139),
.B2(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_175),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_208),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_179),
.C(n_177),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_206),
.C(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_179),
.C(n_182),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_210),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_190),
.B1(n_195),
.B2(n_181),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_183),
.C(n_106),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_186),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_196),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_187),
.B1(n_193),
.B2(n_200),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_223),
.B1(n_219),
.B2(n_225),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_195),
.C(n_121),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_209),
.C(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_173),
.B(n_169),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_0),
.B(n_1),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_212),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_215),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_230),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_235),
.C(n_1),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_214),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_169),
.C(n_139),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_122),
.C(n_107),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_15),
.C(n_14),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_216),
.B(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_223),
.C(n_13),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_0),
.B(n_1),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_43),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_235),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_236),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_254),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_240),
.C(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_233),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_242),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_258),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_4),
.C(n_6),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_7),
.C(n_8),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_250),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_265),
.B(n_263),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_267),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_7),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_270),
.C(n_8),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_8),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_273),
.A2(n_43),
.B(n_216),
.Y(n_274)
);


endmodule