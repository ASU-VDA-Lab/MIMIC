module real_jpeg_2394_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_0),
.B(n_29),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_0),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_0),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_0),
.B(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_0),
.B(n_134),
.Y(n_221)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_29),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_2),
.B(n_36),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_2),
.B(n_47),
.Y(n_192)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_2),
.B(n_59),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_2),
.B(n_79),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_3),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_3),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_3),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_3),
.B(n_24),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_5),
.B(n_59),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_5),
.B(n_110),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_5),
.B(n_79),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_134),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_5),
.B(n_24),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_6),
.B(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_6),
.B(n_29),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_6),
.B(n_47),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_6),
.B(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_6),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_11),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_11),
.B(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_11),
.B(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_11),
.B(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_11),
.B(n_110),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_11),
.B(n_79),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_36),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_12),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_12),
.B(n_29),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_12),
.B(n_47),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_12),
.B(n_59),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_14),
.B(n_29),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_14),
.B(n_47),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_14),
.B(n_59),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_14),
.B(n_36),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_14),
.B(n_79),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_14),
.B(n_110),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_14),
.B(n_134),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_14),
.B(n_24),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_88),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_87),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_62),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_62),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_48),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_41),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_73),
.C(n_74),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_23),
.A2(n_39),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_24),
.Y(n_159)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_38),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_32),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_42),
.C(n_45),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_28),
.A2(n_52),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_28),
.B(n_331),
.C(n_332),
.Y(n_343)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_29),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_32),
.A2(n_33),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_33),
.B(n_109),
.C(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_35),
.B(n_167),
.Y(n_315)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_42),
.A2(n_43),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_43),
.B(n_101),
.C(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_45),
.A2(n_46),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_55),
.C(n_57),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_46),
.B(n_102),
.C(n_211),
.Y(n_316)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_47),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.C(n_54),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_54),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_56),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_58),
.B1(n_77),
.B2(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_57),
.A2(n_58),
.B1(n_121),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_77),
.C(n_80),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_58),
.B(n_121),
.C(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_59),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_84),
.C(n_85),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_64),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_76),
.C(n_81),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_66),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_71),
.C(n_72),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_68),
.A2(n_69),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_68),
.A2(n_69),
.B1(n_135),
.B2(n_373),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_69),
.B(n_131),
.C(n_135),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_69),
.B(n_345),
.C(n_348),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_73),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_73),
.A2(n_128),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_73),
.B(n_311),
.C(n_315),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_81),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_106),
.C(n_108),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_78),
.B1(n_108),
.B2(n_109),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_77),
.A2(n_78),
.B1(n_182),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_78),
.B(n_182),
.C(n_183),
.Y(n_181)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_84),
.B(n_85),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_139),
.B(n_403),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_136),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_91),
.B(n_136),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_113),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_96),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_97),
.A2(n_98),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_100),
.B(n_105),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_101),
.A2(n_102),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_107),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_108),
.A2(n_109),
.B1(n_221),
.B2(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_108),
.A2(n_109),
.B1(n_133),
.B2(n_245),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_111),
.B(n_226),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_113),
.B(n_388),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_126),
.C(n_130),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_114),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.C(n_123),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_115),
.A2(n_116),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_119),
.B(n_123),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.C(n_122),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_120),
.B(n_122),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_121),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_121),
.A2(n_161),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_126),
.B(n_130),
.Y(n_392)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_131),
.A2(n_132),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_133),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_133),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_133),
.A2(n_149),
.B1(n_179),
.B2(n_245),
.Y(n_318)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_134),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_135),
.Y(n_373)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_385),
.B(n_400),
.Y(n_139)
);

OAI31xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_335),
.A3(n_374),
.B(n_379),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_303),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_227),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_195),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_144),
.B(n_195),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_162),
.C(n_185),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_145),
.B(n_300),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_145),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_152),
.CI(n_156),
.CON(n_145),
.SN(n_145)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_146),
.B(n_152),
.C(n_156),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_147),
.A2(n_148),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_148),
.A2(n_179),
.B(n_245),
.C(n_319),
.Y(n_357)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_176),
.B1(n_179),
.B2(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_150),
.B(n_151),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_155),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_155),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_158),
.B(n_177),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_158),
.B(n_206),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_159),
.B(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_162),
.B(n_185),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_173),
.B2(n_184),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_174),
.C(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_170),
.C(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_180),
.B2(n_181),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_178),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_193),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_186),
.B(n_189),
.CI(n_193),
.CON(n_290),
.SN(n_290)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.C(n_192),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_192),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_238),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g412 ( 
.A(n_195),
.Y(n_412)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_213),
.CI(n_214),
.CON(n_195),
.SN(n_195)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_196),
.B(n_213),
.C(n_214),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_197),
.B(n_200),
.C(n_207),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_207),
.B2(n_208),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_201),
.B(n_203),
.C(n_205),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_211),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_216),
.B(n_217),
.C(n_219),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_221),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_221),
.B(n_223),
.C(n_225),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_298),
.B(n_302),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_286),
.B(n_297),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_258),
.B(n_285),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_249),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_249),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_241),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_235),
.CI(n_236),
.CON(n_250),
.SN(n_250)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_237),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_239),
.C(n_241),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_247),
.C(n_248),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.C(n_257),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_282),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_250),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_279),
.B(n_284),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_270),
.B(n_278),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_266),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_266),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_264),
.C(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_273),
.B(n_277),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_288),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_293),
.C(n_294),
.Y(n_301)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_290),
.Y(n_411)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_304),
.A2(n_381),
.B(n_382),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_334),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_305),
.B(n_334),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_306),
.B(n_308),
.C(n_321),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_320),
.B2(n_321),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g407 ( 
.A(n_309),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_316),
.CI(n_317),
.CON(n_309),
.SN(n_309)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_316),
.C(n_317),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_326),
.C(n_327),
.Y(n_350)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_332),
.B2(n_333),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g379 ( 
.A1(n_336),
.A2(n_375),
.B(n_380),
.C(n_383),
.D(n_384),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_361),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_337),
.B(n_361),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_350),
.C(n_351),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_338),
.A2(n_339),
.B1(n_351),
.B2(n_352),
.Y(n_377)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_349),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_343),
.C(n_344),
.Y(n_362)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_347),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_356),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_357),
.C(n_358),
.Y(n_368)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_359),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_364),
.C(n_367),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_367),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_369),
.CI(n_370),
.CON(n_367),
.SN(n_367)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_369),
.C(n_370),
.Y(n_396)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_378),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_397),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_386),
.A2(n_401),
.B(n_402),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_390),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.C(n_396),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g398 ( 
.A(n_391),
.B(n_393),
.CI(n_396),
.CON(n_398),
.SN(n_398)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_394),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_399),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_398),
.Y(n_410)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);


endmodule