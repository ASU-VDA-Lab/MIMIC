module fake_jpeg_13400_n_245 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_44),
.Y(n_80)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_16),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g103 ( 
.A(n_45),
.Y(n_103)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_51),
.Y(n_83)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_2),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_18),
.B(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_4),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_4),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_72),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_37),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_30),
.B(n_4),
.CON(n_72),
.SN(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_21),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_74),
.A2(n_76),
.B1(n_85),
.B2(n_92),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_27),
.B1(n_28),
.B2(n_26),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_95),
.B(n_93),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_33),
.B1(n_36),
.B2(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_8),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_21),
.B1(n_32),
.B2(n_31),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_104),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_43),
.A2(n_26),
.B1(n_6),
.B2(n_7),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_5),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_8),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_144),
.B1(n_124),
.B2(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_122),
.Y(n_156)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_72),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_74),
.B1(n_102),
.B2(n_60),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_129),
.B(n_53),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_100),
.B(n_111),
.C(n_87),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_136),
.B(n_119),
.C(n_138),
.Y(n_149)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_134),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_133),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_45),
.B(n_37),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_132),
.Y(n_168)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_8),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_12),
.A3(n_37),
.B1(n_100),
.B2(n_87),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_81),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_146),
.Y(n_158)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_113),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_86),
.B1(n_98),
.B2(n_90),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_94),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_167),
.B(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_126),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_120),
.C(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_164),
.C(n_158),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_161),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_115),
.B1(n_121),
.B2(n_130),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_170),
.B1(n_154),
.B2(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_123),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_165),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_137),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_145),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_113),
.B1(n_122),
.B2(n_127),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_168),
.B(n_164),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_161),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_162),
.B(n_147),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_149),
.B(n_151),
.C(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_183),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_186),
.B(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_156),
.B(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_185),
.B(n_188),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_147),
.Y(n_191)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_169),
.C(n_166),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_169),
.C(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_157),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_182),
.C(n_172),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_208),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_172),
.C(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_178),
.B1(n_179),
.B2(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_176),
.B1(n_186),
.B2(n_189),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_213),
.A2(n_204),
.B1(n_208),
.B2(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_215),
.Y(n_219)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_222),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_198),
.B1(n_193),
.B2(n_174),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_224),
.B1(n_216),
.B2(n_205),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_192),
.B(n_175),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_206),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_205),
.B1(n_194),
.B2(n_177),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_227),
.Y(n_235)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_206),
.C(n_188),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_230),
.B(n_218),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_212),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_229),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_221),
.B1(n_220),
.B2(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_228),
.Y(n_236)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_222),
.B(n_221),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_234),
.B(n_173),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_237),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_230),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_241),
.B(n_235),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_240),
.B(n_241),
.CI(n_238),
.CON(n_242),
.SN(n_242)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_243),
.B(n_196),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_242),
.A3(n_215),
.B1(n_157),
.B2(n_190),
.C1(n_184),
.C2(n_170),
.Y(n_245)
);


endmodule