module fake_jpeg_424_n_431 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_50),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_8),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_68),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_8),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_79),
.Y(n_107)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_40),
.B1(n_36),
.B2(n_27),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_83),
.A2(n_92),
.B1(n_120),
.B2(n_71),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_33),
.B1(n_38),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_84),
.A2(n_88),
.B1(n_112),
.B2(n_124),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_38),
.B1(n_28),
.B2(n_16),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_33),
.B1(n_18),
.B2(n_16),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_78),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_43),
.A2(n_27),
.B1(n_64),
.B2(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_45),
.B(n_67),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_46),
.B(n_18),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_66),
.A2(n_24),
.B1(n_19),
.B2(n_29),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_43),
.A2(n_48),
.B1(n_76),
.B2(n_75),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_42),
.B1(n_60),
.B2(n_24),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_144),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_89),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_148),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_151),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_98),
.B1(n_86),
.B2(n_104),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_135),
.A2(n_136),
.B(n_111),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_41),
.A3(n_54),
.B1(n_65),
.B2(n_70),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_74),
.C(n_80),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_153),
.C(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_62),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_92),
.B(n_19),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_163),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_87),
.B(n_44),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_112),
.B1(n_115),
.B2(n_109),
.Y(n_173)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_146),
.Y(n_206)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_149),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_84),
.B(n_0),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_91),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_121),
.B(n_60),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_0),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_157),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_72),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_0),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_161),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_1),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_167),
.Y(n_188)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_99),
.A2(n_47),
.B1(n_52),
.B2(n_59),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_155),
.B1(n_135),
.B2(n_166),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_95),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_61),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_69),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_42),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_1),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_53),
.C(n_37),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_35),
.C(n_29),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_179),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_101),
.B1(n_93),
.B2(n_116),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_101),
.B1(n_93),
.B2(n_116),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_123),
.B1(n_111),
.B2(n_37),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_136),
.B1(n_131),
.B2(n_154),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_180),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_123),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_1),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_2),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_197),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_37),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_144),
.C(n_128),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_2),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_131),
.A2(n_35),
.B1(n_29),
.B2(n_5),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_132),
.A2(n_35),
.B1(n_4),
.B2(n_6),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_127),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_209),
.B(n_230),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_212),
.B(n_214),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_225),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_168),
.B(n_139),
.C(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_147),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_217),
.B(n_227),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_153),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_171),
.C(n_186),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_159),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_224),
.Y(n_248)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_220),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_138),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_171),
.C(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_188),
.B(n_137),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_144),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_231),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_202),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_169),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_193),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_232),
.B(n_233),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_240),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_186),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_156),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_184),
.B(n_161),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_183),
.A2(n_150),
.B1(n_133),
.B2(n_141),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_174),
.B1(n_175),
.B2(n_179),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_142),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_197),
.A2(n_158),
.B(n_146),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_182),
.B(n_178),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_148),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_158),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_199),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_245),
.A2(n_186),
.B1(n_187),
.B2(n_173),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_247),
.A2(n_261),
.B(n_269),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_254),
.B1(n_257),
.B2(n_276),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_218),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_268),
.C(n_273),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_210),
.A2(n_187),
.B1(n_204),
.B2(n_177),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_210),
.A2(n_187),
.B1(n_191),
.B2(n_198),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_221),
.A2(n_203),
.B1(n_200),
.B2(n_192),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_201),
.B1(n_195),
.B2(n_176),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_263),
.A2(n_265),
.B1(n_275),
.B2(n_242),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_221),
.A2(n_176),
.B1(n_192),
.B2(n_196),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_225),
.B(n_178),
.C(n_196),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_234),
.A2(n_182),
.B1(n_126),
.B2(n_7),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_270),
.A2(n_238),
.B1(n_230),
.B2(n_222),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_182),
.C(n_126),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_126),
.B1(n_6),
.B2(n_7),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_226),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_4),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_9),
.C(n_10),
.Y(n_304)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_211),
.Y(n_283)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_290),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_239),
.B1(n_219),
.B2(n_215),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_287),
.A2(n_294),
.B1(n_302),
.B2(n_305),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_253),
.A2(n_217),
.B1(n_236),
.B2(n_245),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_250),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_292),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_216),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_293),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_301),
.C(n_251),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_261),
.A2(n_227),
.B1(n_216),
.B2(n_228),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_272),
.B1(n_271),
.B2(n_246),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_237),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_297),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_214),
.B(n_213),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_298),
.A2(n_303),
.B(n_270),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_222),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_262),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_235),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_256),
.A2(n_211),
.B1(n_238),
.B2(n_220),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_280),
.A2(n_9),
.B(n_10),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_308),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_256),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_280),
.B1(n_275),
.B2(n_260),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_307),
.B1(n_305),
.B2(n_289),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_260),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_11),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_11),
.Y(n_309)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_311),
.A2(n_331),
.B1(n_333),
.B2(n_292),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_315),
.Y(n_346)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_252),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_317),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_329),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_299),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_265),
.B(n_250),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_323),
.B(n_282),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_293),
.A2(n_271),
.B1(n_264),
.B2(n_266),
.Y(n_325)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_287),
.A2(n_268),
.B1(n_273),
.B2(n_264),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_297),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_297),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_284),
.A2(n_259),
.B1(n_267),
.B2(n_258),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_281),
.A2(n_262),
.B(n_259),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_294),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_285),
.C(n_295),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_345),
.C(n_357),
.Y(n_360)
);

AOI21xp33_ASAP7_75t_L g340 ( 
.A1(n_322),
.A2(n_298),
.B(n_291),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_340),
.A2(n_319),
.B(n_328),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_348),
.Y(n_375)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_344),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_285),
.C(n_283),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_290),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_353),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_311),
.B(n_290),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_350),
.B(n_351),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_296),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_351),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g363 ( 
.A1(n_352),
.A2(n_327),
.B(n_335),
.C(n_321),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_302),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_329),
.C(n_310),
.Y(n_366)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_330),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_312),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_286),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_306),
.C(n_286),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_338),
.C(n_346),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_368),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_337),
.A2(n_314),
.B1(n_334),
.B2(n_312),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_366),
.Y(n_384)
);

AOI221xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_328),
.B1(n_332),
.B2(n_319),
.C(n_325),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_369),
.C(n_366),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_327),
.B1(n_316),
.B2(n_310),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_342),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_318),
.C(n_333),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_352),
.C(n_357),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_339),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_324),
.C(n_326),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_350),
.C(n_341),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_307),
.Y(n_383)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_361),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_381),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_352),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_380),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_387),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_317),
.B(n_371),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_339),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_373),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_304),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_336),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_288),
.C(n_309),
.Y(n_400)
);

FAx1_ASAP7_75t_SL g390 ( 
.A(n_384),
.B(n_370),
.CI(n_363),
.CON(n_390),
.SN(n_390)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_394),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_385),
.A2(n_336),
.B1(n_363),
.B2(n_369),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_392),
.B(n_11),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_385),
.A2(n_372),
.B1(n_355),
.B2(n_347),
.Y(n_395)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_363),
.B(n_347),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_399),
.B(n_401),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_382),
.A2(n_326),
.B1(n_288),
.B2(n_258),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_400),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_382),
.A2(n_380),
.B(n_379),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_378),
.C(n_389),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_404),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_381),
.C(n_303),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_402),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_390),
.Y(n_419)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_407),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_393),
.B(n_14),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_408),
.B(n_400),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_396),
.A2(n_14),
.B1(n_394),
.B2(n_398),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_411),
.B(n_390),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_410),
.B(n_397),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_413),
.B(n_415),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_412),
.A2(n_401),
.B(n_392),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_414),
.A2(n_419),
.B(n_420),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_417),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_410),
.B(n_409),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_418),
.A2(n_405),
.B(n_403),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_425),
.C(n_405),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_417),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_426),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_411),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_428),
.A2(n_421),
.B(n_427),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_422),
.C(n_404),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_416),
.Y(n_431)
);


endmodule