module fake_jpeg_3111_n_657 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_657);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_657;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_58),
.B(n_62),
.Y(n_145)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_20),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_64),
.B(n_78),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_65),
.Y(n_186)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_28),
.A2(n_0),
.B(n_2),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_67),
.A2(n_42),
.B(n_38),
.Y(n_220)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_71),
.Y(n_193)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_74),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_20),
.B(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_75),
.B(n_76),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_2),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_3),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_79),
.Y(n_233)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_80),
.Y(n_183)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_81),
.Y(n_225)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_23),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_84),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_85),
.Y(n_177)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_88),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_89),
.Y(n_205)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_91),
.Y(n_218)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_97),
.Y(n_187)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_112),
.Y(n_154)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_110),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_21),
.Y(n_111)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_25),
.B(n_3),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_115),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_25),
.B(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_22),
.Y(n_119)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_121),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_22),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_124),
.Y(n_180)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_130),
.Y(n_190)
);

CKINVDCx9p33_ASAP7_75t_R g126 ( 
.A(n_54),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_49),
.Y(n_167)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_127),
.Y(n_196)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_26),
.Y(n_128)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_26),
.Y(n_129)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_129),
.Y(n_234)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_31),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_36),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_36),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_132),
.B(n_49),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_56),
.B1(n_51),
.B2(n_50),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_133),
.A2(n_225),
.B1(n_233),
.B2(n_142),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_56),
.C(n_51),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_134),
.B(n_197),
.C(n_213),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_137),
.B(n_150),
.Y(n_237)
);

CKINVDCx12_ASAP7_75t_R g138 ( 
.A(n_80),
.Y(n_138)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_138),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_56),
.B1(n_51),
.B2(n_50),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_176),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_60),
.A2(n_53),
.B1(n_52),
.B2(n_31),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_45),
.B1(n_52),
.B2(n_39),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_102),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_78),
.A2(n_36),
.B(n_50),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_157),
.A2(n_13),
.B(n_14),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_111),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_165),
.B(n_168),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_53),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_166),
.B(n_178),
.Y(n_257)
);

INVx4_ASAP7_75t_SL g303 ( 
.A(n_167),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_39),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_65),
.A2(n_48),
.B1(n_46),
.B2(n_45),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_48),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_181),
.B(n_185),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_123),
.B(n_46),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_132),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_199),
.B(n_201),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_101),
.B(n_49),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_203),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_74),
.A2(n_91),
.B1(n_79),
.B2(n_83),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_204),
.A2(n_206),
.B1(n_208),
.B2(n_219),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_68),
.A2(n_81),
.B1(n_69),
.B2(n_94),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_85),
.A2(n_44),
.B1(n_42),
.B2(n_38),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_100),
.B(n_44),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_220),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_89),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_212),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_115),
.B(n_44),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_222),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_98),
.A2(n_42),
.B1(n_38),
.B2(n_5),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_90),
.B(n_3),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_116),
.B(n_18),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_228),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_117),
.A2(n_122),
.B1(n_124),
.B2(n_120),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_224),
.A2(n_226),
.B1(n_231),
.B2(n_177),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_127),
.A2(n_18),
.B1(n_6),
.B2(n_7),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_58),
.B(n_4),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_15),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_62),
.B(n_6),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_129),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_16),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_62),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_230),
.B(n_152),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_92),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_157),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_235),
.A2(n_250),
.B1(n_173),
.B2(n_186),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_148),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_236),
.B(n_242),
.Y(n_335)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_158),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_239),
.Y(n_367)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_240),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_190),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_243),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_190),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_244),
.B(n_245),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_156),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_246),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_247),
.Y(n_354)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_164),
.Y(n_248)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_156),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_249),
.B(n_274),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g346 ( 
.A1(n_251),
.A2(n_261),
.B(n_311),
.Y(n_346)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_252),
.Y(n_384)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_153),
.Y(n_254)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_254),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_140),
.A2(n_231),
.B1(n_219),
.B2(n_172),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_255),
.A2(n_283),
.B1(n_291),
.B2(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_256),
.Y(n_350)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_259),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_199),
.A2(n_14),
.B(n_15),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_260),
.A2(n_292),
.B(n_189),
.Y(n_349)
);

BUFx12f_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_263),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_182),
.A2(n_180),
.B1(n_175),
.B2(n_183),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_SL g362 ( 
.A1(n_268),
.A2(n_271),
.B(n_277),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_147),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_269),
.Y(n_376)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_182),
.Y(n_270)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_270),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_175),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_272),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_273),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_156),
.Y(n_274)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_164),
.Y(n_276)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_276),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_180),
.A2(n_183),
.B1(n_167),
.B2(n_194),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_161),
.A2(n_179),
.B1(n_134),
.B2(n_163),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_278),
.Y(n_385)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_136),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_279),
.B(n_281),
.Y(n_365)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_133),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_282),
.B(n_285),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_228),
.A2(n_230),
.B1(n_145),
.B2(n_139),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_147),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_284),
.Y(n_328)
);

INVx3_ASAP7_75t_SL g285 ( 
.A(n_162),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_290),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_162),
.A2(n_214),
.B1(n_146),
.B2(n_221),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_287),
.A2(n_299),
.B1(n_313),
.B2(n_314),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_154),
.B(n_139),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_289),
.Y(n_338)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_136),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_149),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_SL g292 ( 
.A(n_160),
.B(n_214),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_159),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_297),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_225),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_295),
.Y(n_340)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_198),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_298),
.Y(n_364)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_159),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_215),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_152),
.A2(n_202),
.B1(n_209),
.B2(n_171),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_143),
.A2(n_188),
.B1(n_197),
.B2(n_171),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_301),
.A2(n_323),
.B1(n_237),
.B2(n_282),
.Y(n_357)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_147),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_302),
.Y(n_341)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_198),
.B(n_170),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_170),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_306),
.B(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_195),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_155),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_308),
.Y(n_353)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_143),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_312),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_202),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_310),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_196),
.B(n_209),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_188),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_193),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_316),
.Y(n_366)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_169),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_169),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_317),
.B(n_321),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_323),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_172),
.A2(n_205),
.B1(n_177),
.B2(n_218),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_155),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_174),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_322),
.A2(n_270),
.B1(n_285),
.B2(n_284),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_173),
.B(n_233),
.C(n_213),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_324),
.B(n_342),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_241),
.B(n_193),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_337),
.C(n_373),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_281),
.A2(n_207),
.B(n_151),
.C(n_200),
.Y(n_327)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_327),
.A2(n_345),
.B(n_365),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_241),
.A2(n_218),
.B1(n_205),
.B2(n_200),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_330),
.A2(n_342),
.B1(n_345),
.B2(n_358),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_207),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_291),
.A2(n_186),
.B1(n_174),
.B2(n_184),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_303),
.A2(n_184),
.B1(n_189),
.B2(n_151),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_349),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_184),
.B1(n_300),
.B2(n_283),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_355),
.A2(n_356),
.B1(n_385),
.B2(n_378),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_303),
.A2(n_255),
.B1(n_311),
.B2(n_266),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g412 ( 
.A1(n_357),
.A2(n_262),
.B1(n_240),
.B2(n_269),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_280),
.A2(n_257),
.B1(n_265),
.B2(n_264),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_320),
.A2(n_311),
.B1(n_239),
.B2(n_301),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_363),
.B1(n_375),
.B2(n_321),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_267),
.A2(n_260),
.B1(n_251),
.B2(n_304),
.Y(n_363)
);

AOI32xp33_ASAP7_75t_L g371 ( 
.A1(n_292),
.A2(n_261),
.A3(n_258),
.B1(n_279),
.B2(n_304),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_247),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_238),
.B(n_254),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_309),
.A2(n_314),
.B1(n_307),
.B2(n_290),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_379),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_373),
.B(n_297),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_386),
.B(n_391),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_336),
.B(n_306),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_417),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_336),
.B(n_286),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_256),
.C(n_293),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_392),
.B(n_415),
.C(n_420),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_SL g393 ( 
.A(n_371),
.B(n_243),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_393),
.A2(n_328),
.B(n_333),
.Y(n_448)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_381),
.Y(n_398)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_355),
.A2(n_246),
.B1(n_317),
.B2(n_316),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_400),
.A2(n_406),
.B1(n_411),
.B2(n_419),
.Y(n_446)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_298),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_402),
.B(n_421),
.Y(n_467)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_403),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_428),
.C(n_376),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_296),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_405),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_348),
.A2(n_295),
.B1(n_322),
.B2(n_308),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_408),
.Y(n_435)
);

AOI32xp33_ASAP7_75t_L g408 ( 
.A1(n_385),
.A2(n_302),
.A3(n_263),
.B1(n_252),
.B2(n_253),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_335),
.B(n_289),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_409),
.B(n_410),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_358),
.B(n_259),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_348),
.A2(n_272),
.B1(n_248),
.B2(n_276),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_422),
.B1(n_367),
.B2(n_353),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_413),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_382),
.Y(n_414)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_275),
.C(n_262),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_332),
.B(n_275),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_416),
.B(n_418),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_351),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_334),
.B(n_370),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_356),
.B(n_363),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_326),
.B(n_347),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_357),
.A2(n_359),
.B1(n_330),
.B2(n_365),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_341),
.B(n_366),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_429),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_362),
.B(n_346),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_354),
.Y(n_447)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_425),
.Y(n_461)
);

OA22x2_ASAP7_75t_L g426 ( 
.A1(n_327),
.A2(n_365),
.B1(n_349),
.B2(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_431),
.Y(n_465)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_427),
.Y(n_462)
);

AOI21xp33_ASAP7_75t_L g428 ( 
.A1(n_372),
.A2(n_366),
.B(n_351),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_340),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_333),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_430),
.B(n_380),
.Y(n_475)
);

OA22x2_ASAP7_75t_L g431 ( 
.A1(n_379),
.A2(n_350),
.B1(n_333),
.B2(n_374),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_329),
.B(n_339),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_433),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_367),
.A2(n_329),
.B1(n_339),
.B2(n_350),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_434),
.B(n_457),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_328),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_436),
.B(n_426),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_388),
.B(n_369),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_440),
.B(n_445),
.Y(n_507)
);

BUFx12_ASAP7_75t_L g443 ( 
.A(n_430),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_443),
.Y(n_486)
);

XOR2x1_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_375),
.Y(n_445)
);

XNOR2x1_ASAP7_75t_SL g481 ( 
.A(n_447),
.B(n_392),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_448),
.A2(n_463),
.B(n_474),
.Y(n_491)
);

NAND3xp33_ASAP7_75t_L g497 ( 
.A(n_450),
.B(n_468),
.C(n_470),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_422),
.A2(n_353),
.B1(n_344),
.B2(n_368),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_451),
.A2(n_390),
.B1(n_425),
.B2(n_413),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_388),
.B(n_368),
.C(n_369),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_456),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_391),
.B(n_343),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_421),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_395),
.B(n_383),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_389),
.A2(n_376),
.B(n_352),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_383),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_387),
.B(n_343),
.C(n_374),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_414),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_417),
.B(n_361),
.Y(n_470)
);

NOR4xp25_ASAP7_75t_SL g474 ( 
.A(n_424),
.B(n_361),
.C(n_380),
.D(n_352),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_475),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_477),
.Y(n_515)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_449),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_478),
.Y(n_548)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_479),
.B(n_480),
.Y(n_536)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_481),
.B(n_492),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_464),
.B(n_394),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_482),
.B(n_499),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_483),
.A2(n_490),
.B1(n_458),
.B2(n_469),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_460),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_484),
.B(n_493),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_439),
.A2(n_396),
.B1(n_398),
.B2(n_390),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_487),
.A2(n_434),
.B1(n_446),
.B2(n_400),
.Y(n_517)
);

A2O1A1O1Ixp25_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_432),
.B(n_389),
.C(n_415),
.D(n_433),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_489),
.A2(n_495),
.B(n_498),
.Y(n_538)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_441),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_454),
.A2(n_419),
.B(n_399),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_494),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_439),
.A2(n_397),
.B1(n_411),
.B2(n_406),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_467),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_496),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_435),
.A2(n_444),
.B1(n_461),
.B2(n_465),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_466),
.B(n_402),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_441),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_500),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_457),
.B(n_386),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_501),
.B(n_504),
.Y(n_525)
);

A2O1A1O1Ixp25_ASAP7_75t_L g502 ( 
.A1(n_472),
.A2(n_426),
.B(n_427),
.C(n_401),
.D(n_425),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_502),
.A2(n_408),
.B(n_452),
.Y(n_540)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_503),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_407),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_467),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_506),
.B(n_512),
.Y(n_521)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_451),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_508),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_466),
.B(n_426),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_509),
.B(n_511),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g510 ( 
.A1(n_465),
.A2(n_431),
.B(n_413),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_SL g518 ( 
.A1(n_510),
.A2(n_445),
.B(n_436),
.C(n_474),
.Y(n_518)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_438),
.B(n_360),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_513),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_438),
.B(n_431),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_514),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_498),
.A2(n_461),
.B1(n_446),
.B2(n_448),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_516),
.A2(n_522),
.B1(n_532),
.B2(n_533),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_517),
.A2(n_527),
.B1(n_495),
.B2(n_476),
.Y(n_570)
);

A2O1A1Ixp33_ASAP7_75t_L g571 ( 
.A1(n_518),
.A2(n_546),
.B(n_497),
.C(n_486),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_514),
.A2(n_505),
.B1(n_508),
.B2(n_509),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_437),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_523),
.B(n_481),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_485),
.B(n_440),
.C(n_437),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_524),
.B(n_526),
.C(n_535),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_453),
.C(n_447),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_487),
.A2(n_413),
.B1(n_455),
.B2(n_397),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_491),
.A2(n_463),
.B(n_471),
.Y(n_530)
);

AO21x1_ASAP7_75t_L g560 ( 
.A1(n_530),
.A2(n_540),
.B(n_541),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_505),
.A2(n_458),
.B1(n_431),
.B2(n_473),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_507),
.B(n_456),
.C(n_452),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_491),
.A2(n_443),
.B(n_360),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_504),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_542),
.B(n_477),
.Y(n_574)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_513),
.Y(n_545)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_545),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_510),
.A2(n_443),
.B(n_384),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_496),
.B(n_384),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_547),
.B(n_501),
.Y(n_566)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_528),
.Y(n_550)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_550),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_546),
.B(n_510),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_551),
.B(n_558),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_533),
.A2(n_505),
.B1(n_511),
.B2(n_486),
.Y(n_552)
);

INVx11_ASAP7_75t_L g580 ( 
.A(n_552),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_529),
.B(n_488),
.Y(n_554)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_554),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_529),
.B(n_503),
.Y(n_555)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_555),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_520),
.B(n_492),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_556),
.B(n_568),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_557),
.B(n_577),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_521),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_536),
.Y(n_559)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_559),
.Y(n_599)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_549),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_562),
.Y(n_587)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_539),
.Y(n_562)
);

BUFx5_ASAP7_75t_L g563 ( 
.A(n_537),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_563),
.B(n_566),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_543),
.B(n_493),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_564),
.B(n_565),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_543),
.B(n_500),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_523),
.B(n_489),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g569 ( 
.A(n_520),
.B(n_502),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_525),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_570),
.A2(n_516),
.B1(n_541),
.B2(n_534),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_571),
.A2(n_518),
.B(n_545),
.Y(n_602)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_572),
.B(n_573),
.Y(n_600)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_548),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_574),
.B(n_558),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_544),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_576),
.A2(n_578),
.B1(n_517),
.B2(n_515),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_525),
.B(n_403),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_544),
.A2(n_344),
.B1(n_443),
.B2(n_522),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_582),
.A2(n_585),
.B1(n_570),
.B2(n_578),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_SL g618 ( 
.A(n_583),
.B(n_518),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_553),
.A2(n_531),
.B1(n_534),
.B2(n_527),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_575),
.B(n_524),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_588),
.B(n_591),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_575),
.B(n_538),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_568),
.B(n_526),
.C(n_535),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_592),
.B(n_597),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_569),
.B(n_538),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_594),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_556),
.B(n_530),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_595),
.B(n_560),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_596),
.A2(n_551),
.B1(n_518),
.B2(n_576),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_557),
.B(n_540),
.C(n_519),
.Y(n_597)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_601),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_602),
.Y(n_610)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_606),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_593),
.B(n_554),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_608),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_553),
.C(n_571),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_609),
.A2(n_611),
.B1(n_616),
.B2(n_602),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_591),
.B(n_551),
.C(n_555),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_614),
.C(n_590),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_613),
.B(n_618),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_597),
.B(n_564),
.C(n_565),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_581),
.A2(n_560),
.B(n_577),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_596),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_585),
.A2(n_518),
.B1(n_567),
.B2(n_563),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_599),
.B(n_567),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_617),
.B(n_619),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_586),
.B(n_581),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_600),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_620),
.B(n_589),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_622),
.B(n_624),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_623),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_604),
.B(n_592),
.C(n_584),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_625),
.B(n_626),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_605),
.B(n_582),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_629),
.B(n_630),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_614),
.B(n_584),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_603),
.B(n_598),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_633),
.B(n_612),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_610),
.B(n_598),
.Y(n_634)
);

AOI21xp33_ASAP7_75t_L g635 ( 
.A1(n_634),
.A2(n_610),
.B(n_616),
.Y(n_635)
);

AOI21xp33_ASAP7_75t_L g647 ( 
.A1(n_635),
.A2(n_640),
.B(n_636),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_634),
.A2(n_608),
.B(n_583),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_639),
.A2(n_638),
.B1(n_626),
.B2(n_623),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_627),
.A2(n_604),
.B(n_609),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_641),
.B(n_642),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_611),
.Y(n_642)
);

FAx1_ASAP7_75t_SL g644 ( 
.A(n_639),
.B(n_624),
.CI(n_621),
.CON(n_644),
.SN(n_644)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_644),
.A2(n_580),
.B(n_631),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_645),
.A2(n_646),
.B(n_647),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_SL g646 ( 
.A(n_637),
.B(n_625),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_SL g649 ( 
.A(n_643),
.B(n_579),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_649),
.B(n_632),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_650),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_652),
.A2(n_648),
.B(n_644),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_653),
.A2(n_651),
.B(n_613),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_655),
.B(n_654),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_656),
.B(n_632),
.Y(n_657)
);


endmodule