module real_aes_1420_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_20;
wire n_18;
wire n_10;
HB1xp67_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
OAI221xp5_ASAP7_75t_L g16 ( .A1(n_1), .A2(n_4), .B1(n_14), .B2(n_17), .C(n_18), .Y(n_16) );
OAI211xp5_ASAP7_75t_L g12 ( .A1(n_2), .A2(n_10), .B(n_13), .C(n_14), .Y(n_12) );
INVx3_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
AOI321xp33_ASAP7_75t_L g9 ( .A1(n_6), .A2(n_7), .A3(n_10), .B1(n_11), .B2(n_12), .C(n_15), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_10), .B(n_16), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_11), .Y(n_14) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
endmodule