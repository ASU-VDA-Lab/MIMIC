module fake_jpeg_27697_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVxp67_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_12),
.B1(n_0),
.B2(n_19),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_8),
.B(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_8),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_19),
.C(n_18),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_19),
.C(n_20),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_21),
.B1(n_9),
.B2(n_15),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_31),
.B1(n_37),
.B2(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_32),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_14),
.B1(n_13),
.B2(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

OR2x6_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_20),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_0),
.B(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_35),
.B1(n_43),
.B2(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_51),
.C(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_45),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_55),
.C(n_48),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_6),
.Y(n_59)
);


endmodule