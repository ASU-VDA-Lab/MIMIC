module fake_jpeg_20526_n_26 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_4),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

AOI22xp33_ASAP7_75t_SL g9 ( 
.A1(n_3),
.A2(n_6),
.B1(n_5),
.B2(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_0),
.B(n_6),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

AO22x1_ASAP7_75t_SL g15 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_19),
.C(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_17),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_11),
.B(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_12),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_8),
.Y(n_21)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_12),
.B1(n_9),
.B2(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_22),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_19),
.Y(n_25)
);

AOI332xp33_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_10),
.A3(n_14),
.B1(n_15),
.B2(n_20),
.B3(n_23),
.C1(n_24),
.C2(n_22),
.Y(n_26)
);


endmodule