module fake_jpeg_30070_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_7),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_19),
.Y(n_69)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_25),
.B1(n_32),
.B2(n_29),
.Y(n_60)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_24),
.B1(n_17),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_59),
.B1(n_74),
.B2(n_75),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_92),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_36),
.C(n_26),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_82),
.Y(n_130)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_35),
.B1(n_24),
.B2(n_36),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_35),
.B1(n_24),
.B2(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_35),
.B1(n_37),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_77),
.B1(n_80),
.B2(n_84),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_29),
.B1(n_19),
.B2(n_33),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_34),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_19),
.B1(n_32),
.B2(n_28),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_37),
.B1(n_22),
.B2(n_23),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_35),
.B1(n_37),
.B2(n_30),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_88),
.B1(n_55),
.B2(n_67),
.Y(n_126)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_26),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_51),
.B(n_23),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_101),
.B(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_104),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_54),
.A3(n_50),
.B1(n_34),
.B2(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_50),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_18),
.B1(n_34),
.B2(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_109),
.A2(n_131),
.B1(n_56),
.B2(n_79),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_62),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_114),
.Y(n_146)
);

CKINVDCx10_ASAP7_75t_R g111 ( 
.A(n_65),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_9),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_1),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_122),
.Y(n_137)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_34),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_34),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_66),
.B1(n_79),
.B2(n_56),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_63),
.B(n_34),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_129),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

CKINVDCx12_ASAP7_75t_R g132 ( 
.A(n_128),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_63),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_18),
.B1(n_3),
.B2(n_2),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_130),
.A2(n_71),
.B(n_57),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_89),
.C(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_70),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_144),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_86),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_94),
.B(n_98),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_156),
.B(n_111),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_95),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_70),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_93),
.B(n_66),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_116),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_124),
.B1(n_125),
.B2(n_97),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_65),
.B(n_90),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_131),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_2),
.CI(n_3),
.CON(n_163),
.SN(n_163)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_163),
.B(n_12),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_113),
.B1(n_95),
.B2(n_93),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_164),
.A2(n_170),
.B1(n_178),
.B2(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_109),
.B1(n_108),
.B2(n_110),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_155),
.B1(n_157),
.B2(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_136),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_175),
.B(n_179),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_102),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_181),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_109),
.B(n_131),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_187),
.B(n_195),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_102),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_109),
.B1(n_131),
.B2(n_116),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_142),
.B(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_96),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_186),
.B(n_188),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_134),
.B(n_140),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_189),
.B(n_192),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_119),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_196),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_96),
.B1(n_120),
.B2(n_118),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_107),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_163),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_120),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_134),
.B(n_128),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_144),
.B(n_8),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_141),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_209),
.B(n_191),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_203),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_137),
.C(n_142),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_226),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_175),
.B(n_163),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_204),
.B(n_210),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_152),
.A3(n_137),
.B1(n_135),
.B2(n_132),
.C1(n_147),
.C2(n_159),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_132),
.B(n_151),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_152),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_174),
.A2(n_151),
.B(n_153),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_152),
.C(n_158),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_147),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_158),
.C(n_153),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_159),
.C(n_160),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_4),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_231),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_206),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_250),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_222),
.A2(n_182),
.B1(n_170),
.B2(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_166),
.Y(n_236)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_217),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_191),
.C(n_169),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_243),
.C(n_226),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_221),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_214),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_248),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_169),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_215),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_199),
.A2(n_178),
.B1(n_192),
.B2(n_181),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_217),
.B1(n_211),
.B2(n_213),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_178),
.B1(n_228),
.B2(n_164),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_253),
.B1(n_213),
.B2(n_218),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_222),
.A2(n_185),
.B1(n_180),
.B2(n_168),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_260),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_254),
.A2(n_211),
.B1(n_209),
.B2(n_205),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_263),
.B1(n_269),
.B2(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_261),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_254),
.A2(n_212),
.B1(n_208),
.B2(n_201),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_232),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_264),
.B(n_273),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_219),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_272),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_236),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_268),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_240),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_233),
.A2(n_204),
.B(n_227),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_229),
.C(n_239),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_241),
.C(n_210),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_238),
.B(n_234),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_237),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_288),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_229),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_260),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_267),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_283),
.Y(n_293)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

A2O1A1O1Ixp25_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_246),
.B(n_235),
.C(n_247),
.D(n_220),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_290),
.B1(n_255),
.B2(n_261),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_245),
.B1(n_252),
.B2(n_216),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_278),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_292),
.B(n_302),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_272),
.C(n_270),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_297),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_303),
.Y(n_308)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_258),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_245),
.B1(n_270),
.B2(n_266),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_300),
.B1(n_167),
.B2(n_230),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_276),
.A2(n_253),
.B1(n_250),
.B2(n_249),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_241),
.C(n_240),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_284),
.C(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_305),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_279),
.C(n_280),
.Y(n_305)
);

OAI221xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_288),
.B1(n_286),
.B2(n_257),
.C(n_285),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_306),
.Y(n_321)
);

OAI221xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_285),
.B1(n_283),
.B2(n_242),
.C(n_165),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_301),
.B(n_297),
.Y(n_315)
);

AO22x1_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_230),
.B1(n_242),
.B2(n_225),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_5),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_167),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_314),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_322),
.B(n_6),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_301),
.B1(n_311),
.B2(n_313),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_316),
.A2(n_321),
.B1(n_318),
.B2(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_303),
.C(n_160),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_304),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_5),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_327),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_326),
.B1(n_308),
.B2(n_14),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_320),
.A2(n_308),
.B1(n_8),
.B2(n_9),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_7),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_14),
.C2(n_16),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_324),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_324),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_332),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_16),
.Y(n_336)
);


endmodule