module fake_netlist_6_1562_n_1996 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1996);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1996;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_170),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_91),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_99),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_0),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_10),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_20),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_112),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

BUFx2_ASAP7_75t_SL g219 ( 
.A(n_1),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_80),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_36),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_44),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_32),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_110),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_73),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_54),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_25),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_65),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_0),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_172),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_68),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_70),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_51),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_145),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_117),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_88),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_125),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_59),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_106),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_142),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_21),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_21),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_45),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_75),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_78),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_13),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_151),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_19),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_79),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_132),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_121),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_105),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_53),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_50),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_155),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_61),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_183),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_84),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_38),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_139),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_169),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_89),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_72),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_164),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_77),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_2),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_200),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_137),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_101),
.Y(n_284)
);

BUFx8_ASAP7_75t_SL g285 ( 
.A(n_150),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_58),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_124),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_178),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_51),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_188),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_100),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_46),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_8),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_32),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_49),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_71),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_53),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_143),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_140),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_160),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_25),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_87),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_159),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_41),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_90),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_93),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_66),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_54),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_34),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_45),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_108),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_156),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_36),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_31),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_1),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_196),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_98),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_192),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_180),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_92),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_177),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_14),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_131),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_39),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_9),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_26),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_5),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_203),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_115),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_44),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_14),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_171),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_9),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_122),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_49),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_149),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_46),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_138),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_181),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_2),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_12),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_47),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_168),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_133),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_95),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_176),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_38),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_109),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_83),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_86),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_186),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_185),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_58),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_52),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_147),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_11),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_116),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_153),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_6),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_8),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_19),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_205),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_146),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_103),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_47),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_26),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_59),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_126),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_129),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_63),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_175),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_40),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_20),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_199),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_41),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_107),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_5),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_62),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_165),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_30),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_119),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_4),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_17),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_204),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_182),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_190),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_64),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_67),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_18),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_114),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_206),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_22),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_28),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_193),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_187),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_7),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_113),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_96),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_3),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_118),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_173),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_18),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_57),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_16),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_104),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_3),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_123),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_39),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_7),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_82),
.Y(n_414)
);

BUFx8_ASAP7_75t_SL g415 ( 
.A(n_81),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_166),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_293),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_403),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_316),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_344),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_251),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_231),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_408),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_359),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_257),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_265),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_318),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_247),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_255),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_260),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_268),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_289),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_254),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_272),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_264),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_280),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_232),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_309),
.Y(n_446)
);

INVxp33_ASAP7_75t_SL g447 ( 
.A(n_214),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_279),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_307),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_321),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_368),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_292),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_374),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_351),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_296),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_306),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_302),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_315),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_254),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_378),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_214),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_215),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_317),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_388),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_281),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_332),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_343),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_362),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_366),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_369),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_371),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_254),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_318),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_361),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_286),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_285),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_386),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_361),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_294),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_404),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_212),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_213),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_230),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_233),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_215),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_239),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_240),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_216),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_242),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_245),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_246),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g495 ( 
.A(n_415),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_248),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_269),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_252),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_270),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_218),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_295),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_253),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_249),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_249),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_266),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_266),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_298),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_355),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_216),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_254),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_267),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_275),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_277),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_355),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_276),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_276),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_221),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_254),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_354),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_310),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_354),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_367),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_261),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_474),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_480),
.B(n_218),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_457),
.B(n_235),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_510),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_267),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_478),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_218),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_460),
.B(n_263),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_440),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_510),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_440),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_497),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_518),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_484),
.B(n_267),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_518),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_455),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_485),
.B(n_367),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_486),
.B(n_209),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_426),
.B(n_375),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_476),
.B(n_314),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_462),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_499),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_440),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_515),
.A2(n_383),
.B(n_271),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_437),
.A2(n_376),
.B1(n_324),
.B2(n_384),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_463),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_440),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_488),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_454),
.B(n_446),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_425),
.A2(n_396),
.B1(n_413),
.B2(n_412),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_512),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_429),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_459),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_459),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_433),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_444),
.B(n_500),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_459),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_515),
.B(n_291),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_516),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_513),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_516),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_461),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_442),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_487),
.B(n_209),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_500),
.B(n_431),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_519),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_521),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_431),
.B(n_221),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_489),
.B(n_383),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_521),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_522),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_490),
.B(n_211),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_450),
.B(n_314),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_522),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_492),
.B(n_262),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_481),
.B(n_314),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_483),
.B(n_222),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_493),
.B(n_273),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_417),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_435),
.Y(n_593)
);

OA21x2_ASAP7_75t_L g594 ( 
.A1(n_494),
.A2(n_284),
.B(n_274),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_433),
.B(n_211),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_441),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_496),
.B(n_287),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_435),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_417),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_430),
.B(n_217),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_418),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_498),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_418),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_421),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_441),
.B(n_210),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_436),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_436),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_421),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_590),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_595),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_566),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_550),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_565),
.Y(n_613)
);

INVx6_ASAP7_75t_L g614 ( 
.A(n_588),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_550),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_595),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_600),
.B(n_430),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_529),
.B(n_502),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_524),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_524),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_544),
.B(n_443),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_529),
.A2(n_445),
.B1(n_439),
.B2(n_523),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_524),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_550),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_527),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_536),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_529),
.A2(n_445),
.B1(n_439),
.B2(n_461),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_527),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_447),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_560),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_590),
.B(n_458),
.C(n_456),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_575),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_593),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_528),
.Y(n_635)
);

OAI21xp33_ASAP7_75t_SL g636 ( 
.A1(n_525),
.A2(n_434),
.B(n_432),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_526),
.B(n_447),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_593),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_529),
.B(n_443),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_596),
.B(n_419),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_548),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_528),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_532),
.B(n_545),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_534),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_525),
.B(n_465),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_577),
.B(n_427),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_598),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_559),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_571),
.Y(n_649)
);

AO21x2_ASAP7_75t_L g650 ( 
.A1(n_544),
.A2(n_297),
.B(n_288),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_565),
.B(n_465),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_530),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_531),
.B(n_432),
.Y(n_653)
);

AND3x2_ASAP7_75t_L g654 ( 
.A(n_574),
.B(n_398),
.C(n_479),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_606),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_534),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_533),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_565),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_576),
.B(n_477),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_581),
.B(n_509),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_SL g662 ( 
.A(n_586),
.B(n_420),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_537),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_606),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_607),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_607),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_537),
.Y(n_667)
);

INVxp33_ASAP7_75t_L g668 ( 
.A(n_574),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_538),
.B(n_588),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_533),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_570),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_576),
.B(n_477),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_533),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_539),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_531),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_592),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_592),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_SL g680 ( 
.A(n_551),
.B(n_448),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_592),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_592),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_570),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_546),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_572),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_592),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_572),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_592),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_579),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_580),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_585),
.B(n_482),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_557),
.B(n_219),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_546),
.B(n_434),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_580),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_578),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_578),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_580),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_583),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_579),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_589),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_583),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_533),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_533),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_584),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_583),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_587),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_589),
.B(n_422),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_547),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_602),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_535),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_547),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_588),
.B(n_482),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_602),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_555),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_588),
.B(n_501),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_585),
.B(n_449),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_591),
.A2(n_517),
.B1(n_509),
.B2(n_473),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_591),
.B(n_501),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_538),
.B(n_423),
.Y(n_720)
);

AO22x2_ASAP7_75t_L g721 ( 
.A1(n_551),
.A2(n_234),
.B1(n_303),
.B2(n_326),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_535),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_602),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_568),
.B(n_520),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_587),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_535),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_579),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_579),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_535),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_579),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_549),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_579),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_535),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_543),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_587),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_543),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_535),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_604),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_591),
.B(n_507),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_555),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_556),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_543),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_556),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_591),
.B(n_507),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_543),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_604),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_597),
.B(n_520),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_604),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_597),
.B(n_278),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_573),
.B(n_420),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_556),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_556),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_556),
.Y(n_753)
);

AND2x2_ASAP7_75t_SL g754 ( 
.A(n_594),
.B(n_291),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_573),
.Y(n_755)
);

INVxp33_ASAP7_75t_L g756 ( 
.A(n_558),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_582),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_558),
.A2(n_410),
.B1(n_356),
.B2(n_397),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_556),
.Y(n_759)
);

OAI22x1_ASAP7_75t_L g760 ( 
.A1(n_597),
.A2(n_517),
.B1(n_413),
.B2(n_412),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_563),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_643),
.B(n_597),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_610),
.B(n_616),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_657),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_634),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_657),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_657),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_634),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_671),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_613),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_611),
.B(n_637),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_641),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_709),
.B(n_424),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_610),
.B(n_291),
.Y(n_774)
);

AOI221xp5_ASAP7_75t_L g775 ( 
.A1(n_721),
.A2(n_382),
.B1(n_364),
.B2(n_381),
.C(n_363),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_616),
.A2(n_451),
.B1(n_453),
.B2(n_464),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_754),
.B(n_291),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_623),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_638),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_623),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_754),
.B(n_291),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_630),
.B(n_495),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_677),
.B(n_503),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_710),
.B(n_538),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_710),
.B(n_538),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_709),
.B(n_503),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_714),
.B(n_594),
.Y(n_787)
);

AND2x2_ASAP7_75t_SL g788 ( 
.A(n_680),
.B(n_385),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_750),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_714),
.B(n_594),
.Y(n_790)
);

INVxp33_ASAP7_75t_L g791 ( 
.A(n_668),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_723),
.B(n_594),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_723),
.B(n_604),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_638),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_663),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_609),
.B(n_582),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_653),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_645),
.B(n_217),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_639),
.A2(n_360),
.B1(n_330),
.B2(n_334),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_609),
.B(n_582),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_647),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_734),
.B(n_582),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_660),
.B(n_220),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_684),
.A2(n_282),
.B1(n_283),
.B2(n_290),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_647),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_734),
.B(n_540),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_754),
.B(n_385),
.Y(n_807)
);

INVxp67_ASAP7_75t_L g808 ( 
.A(n_715),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_655),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_736),
.B(n_540),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_663),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_663),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_736),
.B(n_540),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_655),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_656),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_742),
.B(n_553),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_656),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_715),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_742),
.B(n_745),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_653),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_745),
.B(n_553),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_757),
.B(n_553),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_664),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_684),
.B(n_385),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_613),
.B(n_466),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_693),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_701),
.B(n_385),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_674),
.B(n_220),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_757),
.B(n_564),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_740),
.B(n_755),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_650),
.A2(n_385),
.B1(n_336),
.B2(n_341),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_664),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_618),
.B(n_564),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_671),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_614),
.A2(n_347),
.B1(n_322),
.B2(n_350),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_667),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_636),
.A2(n_621),
.B(n_617),
.C(n_691),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_613),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_701),
.B(n_665),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_671),
.B(n_305),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_740),
.B(n_693),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_671),
.B(n_313),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_661),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_758),
.A2(n_370),
.B1(n_377),
.B2(n_379),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_665),
.B(n_564),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_666),
.B(n_567),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_628),
.B(n_468),
.Y(n_847)
);

BUFx2_ASAP7_75t_R g848 ( 
.A(n_626),
.Y(n_848)
);

AND2x6_ASAP7_75t_SL g849 ( 
.A(n_692),
.B(n_469),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_666),
.B(n_567),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_673),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_622),
.B(n_471),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_650),
.A2(n_319),
.B1(n_345),
.B2(n_389),
.Y(n_853)
);

INVx8_ASAP7_75t_L g854 ( 
.A(n_692),
.Y(n_854)
);

INVxp33_ASAP7_75t_SL g855 ( 
.A(n_648),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_636),
.B(n_223),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_673),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_708),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_659),
.B(n_472),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_617),
.A2(n_470),
.B(n_452),
.C(n_438),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_713),
.B(n_391),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_716),
.A2(n_304),
.B1(n_299),
.B2(n_300),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_683),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_708),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_683),
.B(n_567),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_685),
.B(n_394),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_667),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_685),
.B(n_599),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_669),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_718),
.B(n_720),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_669),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_687),
.B(n_599),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_614),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_687),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_739),
.A2(n_308),
.B1(n_301),
.B2(n_320),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_695),
.B(n_599),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_695),
.B(n_601),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_744),
.B(n_323),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_703),
.A2(n_563),
.B(n_561),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_696),
.B(n_601),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_696),
.B(n_601),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_747),
.B(n_325),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_700),
.B(n_603),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_705),
.B(n_603),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_669),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_705),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_676),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_720),
.B(n_650),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_738),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_738),
.Y(n_890)
);

AND2x6_ASAP7_75t_SL g891 ( 
.A(n_692),
.B(n_438),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_746),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_L g893 ( 
.A(n_749),
.B(n_331),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_746),
.B(n_338),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_614),
.B(n_603),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_614),
.A2(n_340),
.B1(n_346),
.B2(n_348),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_748),
.B(n_608),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_748),
.B(n_608),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_649),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_670),
.B(n_608),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_635),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_635),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_719),
.A2(n_241),
.B1(n_223),
.B2(n_414),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_642),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_651),
.B(n_312),
.C(n_311),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_717),
.B(n_352),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_642),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_646),
.B(n_225),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_640),
.B(n_692),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_679),
.B(n_416),
.Y(n_910)
);

AOI221xp5_ASAP7_75t_L g911 ( 
.A1(n_721),
.A2(n_238),
.B1(n_228),
.B2(n_227),
.C(n_224),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_670),
.B(n_563),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_724),
.B(n_452),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_670),
.B(n_675),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_679),
.B(n_225),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_644),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_644),
.Y(n_917)
);

INVxp33_ASAP7_75t_L g918 ( 
.A(n_721),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_670),
.B(n_563),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_675),
.B(n_563),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_676),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_692),
.B(n_721),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_681),
.B(n_226),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_675),
.B(n_704),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_758),
.B(n_504),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_612),
.A2(n_470),
.B(n_562),
.C(n_554),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_690),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_631),
.B(n_504),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_675),
.B(n_563),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_690),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_735),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_788),
.A2(n_662),
.B1(n_760),
.B2(n_756),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_764),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_788),
.A2(n_760),
.B1(n_712),
.B2(n_681),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_901),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_SL g936 ( 
.A(n_771),
.B(n_632),
.C(n_229),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_830),
.B(n_633),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_771),
.B(n_652),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_843),
.B(n_632),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_899),
.B(n_612),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_762),
.B(n_694),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_796),
.B(n_694),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_841),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_853),
.A2(n_624),
.B1(n_615),
.B2(n_698),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_769),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_766),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_853),
.A2(n_624),
.B1(n_615),
.B2(n_698),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_766),
.Y(n_948)
);

NOR2x1p5_ASAP7_75t_L g949 ( 
.A(n_847),
.B(n_224),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_800),
.B(n_697),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_769),
.A2(n_688),
.B1(n_686),
.B2(n_682),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_928),
.B(n_505),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_765),
.B(n_697),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_834),
.A2(n_682),
.B1(n_686),
.B2(n_688),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_808),
.B(n_226),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_797),
.B(n_229),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_768),
.B(n_779),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_794),
.B(n_702),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_L g959 ( 
.A(n_770),
.B(n_831),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_767),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_854),
.B(n_505),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_820),
.B(n_826),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_888),
.A2(n_725),
.B1(n_702),
.B2(n_706),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_SL g964 ( 
.A(n_803),
.B(n_237),
.C(n_236),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_795),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_791),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_902),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_772),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_795),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_801),
.B(n_706),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_811),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_805),
.B(n_707),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_904),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_809),
.B(n_707),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_814),
.B(n_725),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_854),
.B(n_506),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_783),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_770),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_789),
.B(n_654),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_782),
.B(n_236),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_858),
.B(n_237),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_812),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_907),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_855),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_815),
.B(n_735),
.Y(n_985)
);

AO22x1_ASAP7_75t_L g986 ( 
.A1(n_918),
.A2(n_258),
.B1(n_256),
.B2(n_250),
.Y(n_986)
);

AND2x2_ASAP7_75t_SL g987 ( 
.A(n_909),
.B(n_506),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_916),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_817),
.B(n_823),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_917),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_763),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_782),
.B(n_798),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_798),
.B(n_241),
.Y(n_993)
);

NOR2x1p5_ASAP7_75t_L g994 ( 
.A(n_852),
.B(n_227),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_864),
.B(n_244),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_859),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_860),
.A2(n_735),
.B(n_629),
.C(n_625),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_832),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_825),
.B(n_731),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_851),
.B(n_678),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_770),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_834),
.B(n_731),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_825),
.B(n_731),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_857),
.B(n_678),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_863),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_770),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_786),
.B(n_508),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_874),
.B(n_678),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_SL g1009 ( 
.A1(n_922),
.A2(n_854),
.B1(n_925),
.B2(n_803),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_873),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_837),
.A2(n_730),
.B(n_727),
.C(n_728),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_SL g1012 ( 
.A(n_848),
.B(n_244),
.Y(n_1012)
);

AOI22x1_ASAP7_75t_L g1013 ( 
.A1(n_886),
.A2(n_761),
.B1(n_759),
.B2(n_753),
.Y(n_1013)
);

AND2x4_ASAP7_75t_SL g1014 ( 
.A(n_773),
.B(n_386),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_889),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_873),
.B(n_689),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_819),
.B(n_727),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_839),
.B(n_259),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_870),
.B(n_727),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_859),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_828),
.B(n_259),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_828),
.B(n_353),
.Y(n_1022)
);

CKINVDCx11_ASAP7_75t_R g1023 ( 
.A(n_849),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_776),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_838),
.B(n_541),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_773),
.B(n_508),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_836),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_818),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_836),
.B(n_728),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_773),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_891),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_867),
.B(n_728),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_818),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_838),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_890),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_908),
.B(n_353),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_861),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_867),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_844),
.B(n_238),
.C(n_228),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_905),
.B(n_541),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_869),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_861),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_913),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_908),
.B(n_357),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_892),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_840),
.A2(n_732),
.B1(n_689),
.B2(n_699),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_871),
.B(n_732),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_860),
.B(n_514),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_840),
.B(n_514),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_866),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_885),
.B(n_732),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_885),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_887),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_887),
.Y(n_1054)
);

AND2x6_ASAP7_75t_L g1055 ( 
.A(n_787),
.B(n_743),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_842),
.A2(n_699),
.B1(n_689),
.B2(n_711),
.Y(n_1056)
);

NOR2x2_ASAP7_75t_L g1057 ( 
.A(n_844),
.B(n_386),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_878),
.B(n_357),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_856),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_921),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_921),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_845),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_862),
.B(n_358),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_875),
.B(n_358),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_856),
.B(n_743),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_878),
.B(n_243),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_L g1067 ( 
.A(n_906),
.B(n_743),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_846),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_777),
.B(n_759),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_894),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_842),
.B(n_689),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_850),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_777),
.B(n_753),
.Y(n_1073)
);

OR2x2_ASAP7_75t_SL g1074 ( 
.A(n_775),
.B(n_428),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_781),
.A2(n_629),
.B1(n_625),
.B2(n_620),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_931),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_807),
.B(n_753),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_778),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_784),
.B(n_751),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_927),
.B(n_930),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_865),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_894),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_L g1083 ( 
.A(n_913),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_915),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_882),
.B(n_542),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_882),
.B(n_542),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_906),
.B(n_243),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_785),
.B(n_552),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_793),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_790),
.A2(n_792),
.B(n_833),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_806),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_780),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_810),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_804),
.B(n_365),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_802),
.A2(n_620),
.B1(n_619),
.B2(n_627),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_915),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_896),
.B(n_365),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_911),
.B(n_552),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_903),
.B(n_372),
.Y(n_1099)
);

NAND2x1p5_ASAP7_75t_L g1100 ( 
.A(n_910),
.B(n_699),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_L g1101 ( 
.A(n_923),
.B(n_751),
.Y(n_1101)
);

OAI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_799),
.A2(n_372),
.B1(n_373),
.B2(n_380),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_914),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_813),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_923),
.B(n_554),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_774),
.A2(n_619),
.B1(n_623),
.B2(n_627),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_SL g1107 ( 
.A(n_774),
.B(n_373),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_868),
.B(n_751),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_910),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_872),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_824),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1076),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_966),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_937),
.Y(n_1114)
);

NOR2x1p5_ASAP7_75t_L g1115 ( 
.A(n_984),
.B(n_250),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_978),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_959),
.A2(n_941),
.B(n_1090),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_992),
.A2(n_926),
.B(n_824),
.C(n_827),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_962),
.B(n_895),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1043),
.A2(n_827),
.B1(n_884),
.B2(n_883),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_978),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_941),
.A2(n_924),
.B(n_822),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1021),
.A2(n_881),
.B(n_876),
.C(n_877),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_977),
.B(n_880),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_939),
.B(n_835),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_978),
.B(n_699),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1001),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_980),
.B(n_893),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_991),
.B(n_816),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1059),
.A2(n_821),
.B1(n_829),
.B2(n_897),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_993),
.A2(n_900),
.B(n_898),
.C(n_919),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_968),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_1011),
.A2(n_929),
.A3(n_920),
.B(n_912),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1076),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_938),
.B(n_327),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1043),
.A2(n_256),
.B1(n_258),
.B2(n_407),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1030),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1090),
.A2(n_722),
.B(n_658),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1028),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_SL g1140 ( 
.A(n_994),
.B(n_380),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_SL g1141 ( 
.A(n_1024),
.B(n_363),
.C(n_381),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_991),
.B(n_328),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_964),
.A2(n_562),
.B(n_569),
.C(n_627),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_1023),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1001),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_998),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1058),
.A2(n_752),
.B(n_711),
.C(n_741),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_936),
.A2(n_401),
.B1(n_390),
.B2(n_402),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_942),
.A2(n_658),
.B(n_672),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1005),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1099),
.A2(n_752),
.B(n_711),
.C(n_741),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_987),
.B(n_390),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_950),
.A2(n_658),
.B(n_672),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_943),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1001),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_943),
.B(n_569),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1037),
.A2(n_752),
.B(n_704),
.C(n_741),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1050),
.B(n_329),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_953),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_953),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_SL g1161 ( 
.A(n_1083),
.B(n_392),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1091),
.B(n_704),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_962),
.B(n_392),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1017),
.A2(n_722),
.B(n_737),
.Y(n_1164)
);

OAI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_952),
.A2(n_370),
.B(n_397),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1013),
.A2(n_879),
.B(n_741),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_1034),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_996),
.B(n_428),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_932),
.B(n_1042),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1087),
.B(n_335),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1079),
.A2(n_1065),
.B(n_1108),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_964),
.A2(n_729),
.B(n_726),
.C(n_711),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_1012),
.Y(n_1173)
);

O2A1O1Ixp5_ASAP7_75t_L g1174 ( 
.A1(n_1022),
.A2(n_704),
.B(n_726),
.C(n_729),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_1034),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_934),
.B(n_337),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1009),
.B(n_395),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1093),
.B(n_726),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1009),
.A2(n_405),
.B1(n_395),
.B2(n_411),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1070),
.A2(n_726),
.B(n_729),
.C(n_399),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_958),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_933),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1079),
.A2(n_737),
.B(n_733),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1020),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1104),
.B(n_729),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1066),
.B(n_364),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1026),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_946),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1026),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1082),
.A2(n_401),
.B(n_402),
.C(n_414),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1036),
.B(n_339),
.Y(n_1191)
);

INVx6_ASAP7_75t_L g1192 ( 
.A(n_1026),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_999),
.B(n_69),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1108),
.A2(n_733),
.B(n_722),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1019),
.B(n_722),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1019),
.B(n_733),
.Y(n_1196)
);

NOR3xp33_ASAP7_75t_L g1197 ( 
.A(n_1044),
.B(n_979),
.C(n_986),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_958),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1033),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1062),
.B(n_405),
.Y(n_1200)
);

AOI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1067),
.A2(n_733),
.B(n_549),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_961),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1025),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_970),
.Y(n_1204)
);

BUFx4f_ASAP7_75t_SL g1205 ( 
.A(n_1031),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1069),
.A2(n_568),
.B(n_409),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1025),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_999),
.Y(n_1208)
);

BUFx4f_ASAP7_75t_L g1209 ( 
.A(n_961),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1069),
.A2(n_733),
.B(n_561),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_948),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1073),
.A2(n_561),
.B(n_411),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1014),
.A2(n_382),
.B1(n_407),
.B2(n_396),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_970),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_949),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1073),
.A2(n_561),
.B(n_409),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_940),
.B(n_342),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1077),
.A2(n_561),
.B(n_549),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1084),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1003),
.B(n_201),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1003),
.B(n_194),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_961),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1077),
.A2(n_349),
.B(n_379),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1039),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1096),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_972),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_936),
.A2(n_377),
.B(n_6),
.C(n_10),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1068),
.B(n_568),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_944),
.A2(n_561),
.B(n_549),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_955),
.B(n_4),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1102),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_947),
.A2(n_549),
.B1(n_16),
.B2(n_17),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_976),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1006),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1072),
.B(n_1081),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1109),
.A2(n_15),
.B(n_23),
.C(n_24),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1101),
.A2(n_568),
.B(n_561),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1000),
.A2(n_568),
.A3(n_27),
.B(n_28),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_976),
.B(n_76),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1110),
.B(n_568),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_972),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1071),
.A2(n_568),
.B(n_74),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_974),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_974),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1018),
.A2(n_24),
.B(n_27),
.C(n_29),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_957),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_957),
.B(n_97),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1000),
.A2(n_568),
.A3(n_34),
.B(n_35),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_976),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_956),
.B(n_33),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_981),
.B(n_995),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1071),
.A2(n_102),
.B(n_189),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1006),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1063),
.A2(n_35),
.B(n_37),
.C(n_40),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1085),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_1255)
);

AO32x1_ASAP7_75t_L g1256 ( 
.A1(n_1111),
.A2(n_42),
.A3(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_SL g1257 ( 
.A(n_1039),
.B(n_1064),
.C(n_1094),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_989),
.B(n_1088),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_997),
.A2(n_141),
.B(n_184),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_L g1260 ( 
.A(n_1007),
.B(n_134),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1040),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1040),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1088),
.B(n_128),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1049),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1117),
.A2(n_1053),
.B(n_1100),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1201),
.A2(n_997),
.B(n_1047),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1135),
.A2(n_1097),
.B(n_1098),
.C(n_1049),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1146),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1235),
.B(n_1129),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1114),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1235),
.A2(n_1010),
.B1(n_945),
.B2(n_1053),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1128),
.A2(n_1010),
.B1(n_945),
.B2(n_1053),
.Y(n_1272)
);

NOR2x1_ASAP7_75t_L g1273 ( 
.A(n_1199),
.B(n_935),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1258),
.B(n_1105),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1138),
.A2(n_1051),
.B(n_1029),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1258),
.B(n_1105),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1150),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1166),
.A2(n_1051),
.B(n_1047),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1171),
.A2(n_1008),
.B(n_1004),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1122),
.A2(n_1053),
.B(n_1100),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1114),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1169),
.A2(n_1085),
.B1(n_1086),
.B2(n_1049),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1118),
.A2(n_963),
.B(n_1032),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1159),
.B(n_1086),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1262),
.B(n_967),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1160),
.B(n_1089),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1156),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1151),
.A2(n_985),
.A3(n_975),
.B(n_1060),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1259),
.A2(n_1046),
.B(n_954),
.Y(n_1289)
);

OAI22x1_ASAP7_75t_L g1290 ( 
.A1(n_1176),
.A2(n_1057),
.B1(n_988),
.B2(n_973),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1181),
.B(n_1089),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1113),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1194),
.A2(n_1183),
.B(n_1164),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1191),
.A2(n_1107),
.B(n_983),
.C(n_990),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1259),
.A2(n_975),
.B(n_985),
.Y(n_1295)
);

BUFx2_ASAP7_75t_SL g1296 ( 
.A(n_1132),
.Y(n_1296)
);

OAI22x1_ASAP7_75t_L g1297 ( 
.A1(n_1224),
.A2(n_1080),
.B1(n_1015),
.B2(n_1035),
.Y(n_1297)
);

AOI211x1_ASAP7_75t_L g1298 ( 
.A1(n_1232),
.A2(n_1045),
.B(n_1054),
.C(n_1074),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1198),
.B(n_1204),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1250),
.A2(n_1048),
.B1(n_1055),
.B2(n_1089),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1123),
.A2(n_1016),
.B(n_1002),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1147),
.A2(n_1157),
.B(n_1174),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1170),
.A2(n_1251),
.B(n_1230),
.C(n_1125),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1149),
.A2(n_1103),
.B(n_1002),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1131),
.A2(n_1016),
.B(n_1078),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1120),
.A2(n_965),
.A3(n_969),
.B(n_971),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1214),
.B(n_960),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1142),
.B(n_1048),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1226),
.B(n_1241),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1243),
.B(n_1052),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1195),
.A2(n_1078),
.B(n_1056),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1180),
.A2(n_1061),
.A3(n_982),
.B(n_1041),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_1116),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_R g1315 ( 
.A(n_1139),
.B(n_1092),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1195),
.A2(n_1078),
.B(n_1095),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1244),
.B(n_1038),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1188),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1200),
.B(n_1027),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1208),
.B(n_951),
.Y(n_1320)
);

OAI21xp33_ASAP7_75t_L g1321 ( 
.A1(n_1148),
.A2(n_1255),
.B(n_1158),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1192),
.B(n_1048),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1196),
.A2(n_1078),
.B(n_1075),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1206),
.A2(n_1055),
.B(n_1106),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1173),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1193),
.A2(n_1221),
.B(n_1220),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1119),
.B(n_1055),
.Y(n_1327)
);

BUFx12f_ASAP7_75t_L g1328 ( 
.A(n_1144),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1153),
.A2(n_1055),
.A3(n_55),
.B(n_56),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1119),
.B(n_1261),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1210),
.A2(n_111),
.B(n_163),
.Y(n_1331)
);

OA21x2_ASAP7_75t_L g1332 ( 
.A1(n_1196),
.A2(n_94),
.B(n_161),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1116),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1116),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1211),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1263),
.A2(n_1162),
.B(n_1260),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1154),
.B(n_1197),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1218),
.A2(n_85),
.B(n_158),
.Y(n_1338)
);

OAI22x1_ASAP7_75t_L g1339 ( 
.A1(n_1177),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1206),
.A2(n_191),
.B(n_148),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1152),
.B(n_1219),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1213),
.B(n_57),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_SL g1343 ( 
.A1(n_1246),
.A2(n_60),
.B(n_62),
.C(n_154),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1112),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1130),
.A2(n_157),
.B(n_60),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1227),
.B(n_1254),
.C(n_1231),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1203),
.B(n_1225),
.Y(n_1347)
);

AOI221x1_ASAP7_75t_L g1348 ( 
.A1(n_1232),
.A2(n_1246),
.B1(n_1257),
.B2(n_1236),
.C(n_1252),
.Y(n_1348)
);

BUFx10_ASAP7_75t_L g1349 ( 
.A(n_1115),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1237),
.A2(n_1172),
.B(n_1162),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1263),
.A2(n_1178),
.B(n_1185),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1167),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1134),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1229),
.A2(n_1126),
.B(n_1242),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1124),
.A2(n_1228),
.B(n_1240),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1208),
.B(n_1193),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1208),
.B(n_1221),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1212),
.A2(n_1216),
.A3(n_1190),
.B(n_1133),
.Y(n_1358)
);

NOR2x1_ASAP7_75t_SL g1359 ( 
.A(n_1167),
.B(n_1175),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1220),
.B(n_1207),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1187),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1175),
.A2(n_1209),
.B1(n_1192),
.B2(n_1179),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1189),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1133),
.A2(n_1136),
.A3(n_1256),
.B(n_1223),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1161),
.B(n_1264),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1239),
.A2(n_1145),
.B(n_1127),
.Y(n_1366)
);

AO32x2_ASAP7_75t_L g1367 ( 
.A1(n_1136),
.A2(n_1256),
.A3(n_1133),
.B1(n_1223),
.B2(n_1238),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1143),
.A2(n_1121),
.B(n_1155),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1217),
.A2(n_1239),
.B(n_1209),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1165),
.B(n_1186),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_R g1371 ( 
.A(n_1140),
.B(n_1205),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1168),
.B(n_1137),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1168),
.B(n_1163),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1245),
.A2(n_1141),
.B(n_1233),
.C(n_1222),
.Y(n_1374)
);

BUFx10_ASAP7_75t_L g1375 ( 
.A(n_1127),
.Y(n_1375)
);

NAND3x1_ASAP7_75t_L g1376 ( 
.A(n_1121),
.B(n_1155),
.C(n_1215),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1202),
.A2(n_1249),
.B(n_1184),
.C(n_1234),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1234),
.B(n_1253),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1234),
.B(n_1253),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1253),
.A2(n_1127),
.B(n_1145),
.C(n_1256),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1145),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1238),
.B(n_1248),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1238),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1248),
.B(n_992),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1248),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1117),
.A2(n_959),
.B(n_1171),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1262),
.B(n_1208),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1116),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1117),
.A2(n_959),
.B(n_1171),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1235),
.B(n_992),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1235),
.B(n_992),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1128),
.A2(n_992),
.B(n_1021),
.C(n_993),
.Y(n_1392)
);

AOI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1176),
.A2(n_992),
.B1(n_771),
.B2(n_844),
.C(n_637),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1192),
.B(n_1239),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1117),
.A2(n_959),
.B(n_1171),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1235),
.B(n_992),
.Y(n_1396)
);

NOR2xp67_ASAP7_75t_L g1397 ( 
.A(n_1261),
.B(n_1070),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_SL g1398 ( 
.A1(n_1118),
.A2(n_1247),
.B(n_1259),
.C(n_1263),
.Y(n_1398)
);

AOI221x1_ASAP7_75t_L g1399 ( 
.A1(n_1259),
.A2(n_992),
.B1(n_1021),
.B2(n_993),
.C(n_1232),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1114),
.B(n_631),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1235),
.B(n_992),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1201),
.A2(n_1138),
.B(n_1166),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1235),
.B(n_992),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1117),
.A2(n_1171),
.B(n_992),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1117),
.A2(n_959),
.B(n_1171),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1135),
.B(n_992),
.C(n_1021),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1235),
.B(n_992),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1114),
.Y(n_1408)
);

BUFx8_ASAP7_75t_SL g1409 ( 
.A(n_1144),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1113),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1117),
.A2(n_959),
.B(n_1171),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1135),
.B(n_992),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1117),
.A2(n_959),
.B(n_1171),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1235),
.B(n_992),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1139),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1114),
.B(n_830),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1146),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1235),
.B(n_992),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1146),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1235),
.B(n_992),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1116),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1113),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1114),
.B(n_631),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1393),
.A2(n_1412),
.B1(n_1406),
.B2(n_1321),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1406),
.B(n_1392),
.C(n_1303),
.Y(n_1426)
);

BUFx2_ASAP7_75t_SL g1427 ( 
.A(n_1325),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1399),
.A2(n_1414),
.B1(n_1401),
.B2(n_1420),
.Y(n_1429)
);

INVx3_ASAP7_75t_SL g1430 ( 
.A(n_1415),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1417),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1267),
.A2(n_1346),
.B(n_1336),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1293),
.A2(n_1304),
.B(n_1265),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1410),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1386),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1340),
.A2(n_1345),
.B(n_1321),
.C(n_1407),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1352),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1396),
.A2(n_1403),
.B1(n_1418),
.B2(n_1282),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1269),
.B(n_1416),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1395),
.A2(n_1411),
.B(n_1405),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1268),
.Y(n_1441)
);

OAI22x1_ASAP7_75t_L g1442 ( 
.A1(n_1282),
.A2(n_1300),
.B1(n_1346),
.B2(n_1342),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1404),
.A2(n_1413),
.B(n_1383),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1398),
.A2(n_1280),
.B(n_1301),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1277),
.Y(n_1445)
);

AOI22x1_ASAP7_75t_L g1446 ( 
.A1(n_1297),
.A2(n_1290),
.B1(n_1345),
.B2(n_1340),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1354),
.A2(n_1266),
.B(n_1350),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1309),
.B(n_1270),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1449)
);

AOI221x1_ASAP7_75t_L g1450 ( 
.A1(n_1339),
.A2(n_1380),
.B1(n_1384),
.B2(n_1294),
.C(n_1337),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1400),
.B(n_1423),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1307),
.Y(n_1452)
);

BUFx10_ASAP7_75t_L g1453 ( 
.A(n_1341),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1270),
.B(n_1281),
.Y(n_1454)
);

BUFx2_ASAP7_75t_SL g1455 ( 
.A(n_1333),
.Y(n_1455)
);

AO31x2_ASAP7_75t_L g1456 ( 
.A1(n_1348),
.A2(n_1312),
.A3(n_1305),
.B(n_1316),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1292),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1370),
.A2(n_1373),
.B1(n_1374),
.B2(n_1369),
.C(n_1365),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1322),
.B(n_1394),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1283),
.A2(n_1295),
.B(n_1351),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1274),
.B(n_1276),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1281),
.Y(n_1462)
);

AO31x2_ASAP7_75t_L g1463 ( 
.A1(n_1323),
.A2(n_1272),
.A3(n_1271),
.B(n_1355),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1382),
.A2(n_1283),
.B(n_1338),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1326),
.B(n_1394),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1333),
.B(n_1352),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1419),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1308),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1333),
.B(n_1273),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1331),
.A2(n_1368),
.B(n_1327),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1289),
.A2(n_1394),
.B1(n_1362),
.B2(n_1315),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1320),
.B(n_1300),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1311),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1377),
.A2(n_1372),
.B(n_1284),
.C(n_1330),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1302),
.A2(n_1332),
.B(n_1317),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1288),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1322),
.A2(n_1287),
.B1(n_1397),
.B2(n_1422),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1332),
.A2(n_1291),
.B(n_1286),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1343),
.A2(n_1319),
.B(n_1335),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1322),
.B(n_1320),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1289),
.A2(n_1318),
.B1(n_1361),
.B2(n_1363),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1306),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1296),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_SL g1484 ( 
.A1(n_1356),
.A2(n_1357),
.B(n_1379),
.C(n_1378),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1288),
.Y(n_1485)
);

AOI22x1_ASAP7_75t_L g1486 ( 
.A1(n_1385),
.A2(n_1285),
.B1(n_1353),
.B2(n_1344),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1285),
.A2(n_1324),
.B1(n_1347),
.B2(n_1397),
.Y(n_1487)
);

OAI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1360),
.A2(n_1366),
.B1(n_1381),
.B2(n_1421),
.C(n_1349),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1288),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1314),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1387),
.B(n_1375),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1387),
.B(n_1375),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1421),
.B(n_1388),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1279),
.A2(n_1349),
.B1(n_1371),
.B2(n_1328),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1314),
.B(n_1388),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1314),
.B(n_1334),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1298),
.A2(n_1376),
.B1(n_1388),
.B2(n_1334),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1313),
.A2(n_1358),
.B(n_1367),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1367),
.A2(n_1364),
.B(n_1329),
.C(n_1358),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1364),
.A2(n_1329),
.B(n_1358),
.C(n_1359),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1329),
.Y(n_1501)
);

O2A1O1Ixp33_ASAP7_75t_SL g1502 ( 
.A1(n_1364),
.A2(n_1392),
.B(n_1303),
.C(n_1340),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1409),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1417),
.Y(n_1504)
);

INVx4_ASAP7_75t_L g1505 ( 
.A(n_1333),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_SL g1508 ( 
.A1(n_1345),
.A2(n_1369),
.B(n_1259),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1404),
.A2(n_1392),
.B(n_1389),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1393),
.A2(n_1412),
.B1(n_1406),
.B2(n_992),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1511)
);

AOI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1393),
.A2(n_1412),
.B1(n_992),
.B2(n_771),
.C(n_1406),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1392),
.A2(n_1412),
.B(n_1303),
.C(n_992),
.Y(n_1513)
);

AOI21xp33_ASAP7_75t_L g1514 ( 
.A1(n_1412),
.A2(n_1406),
.B(n_992),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1410),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1412),
.B(n_1390),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1412),
.A2(n_1406),
.B1(n_1393),
.B2(n_1392),
.Y(n_1517)
);

AO31x2_ASAP7_75t_L g1518 ( 
.A1(n_1399),
.A2(n_1383),
.A3(n_1380),
.B(n_1386),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1416),
.B(n_1114),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1410),
.Y(n_1520)
);

BUFx4_ASAP7_75t_SL g1521 ( 
.A(n_1415),
.Y(n_1521)
);

AOI21xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1412),
.A2(n_855),
.B(n_548),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1417),
.Y(n_1523)
);

NOR2xp67_ASAP7_75t_L g1524 ( 
.A(n_1415),
.B(n_899),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1410),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1386),
.A2(n_1395),
.B(n_1389),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1410),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1417),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1412),
.A2(n_1393),
.B1(n_1406),
.B2(n_992),
.Y(n_1529)
);

AO21x1_ASAP7_75t_L g1530 ( 
.A1(n_1412),
.A2(n_992),
.B(n_1345),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1416),
.B(n_1114),
.Y(n_1531)
);

AO32x2_ASAP7_75t_L g1532 ( 
.A1(n_1272),
.A2(n_1246),
.A3(n_1232),
.B1(n_1367),
.B2(n_1271),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1386),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1406),
.A2(n_1392),
.B(n_1412),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1315),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1406),
.A2(n_1392),
.B(n_1412),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1393),
.A2(n_1412),
.B1(n_1406),
.B2(n_992),
.Y(n_1537)
);

NOR2xp67_ASAP7_75t_L g1538 ( 
.A(n_1415),
.B(n_899),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1408),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1417),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1417),
.Y(n_1542)
);

AO21x2_ASAP7_75t_L g1543 ( 
.A1(n_1386),
.A2(n_1395),
.B(n_1389),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1417),
.Y(n_1544)
);

AO22x1_ASAP7_75t_L g1545 ( 
.A1(n_1412),
.A2(n_992),
.B1(n_1021),
.B2(n_1135),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1333),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1412),
.B(n_1390),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1549)
);

AO22x2_ASAP7_75t_L g1550 ( 
.A1(n_1399),
.A2(n_1406),
.B1(n_1348),
.B2(n_1346),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1333),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1393),
.A2(n_1412),
.B1(n_1406),
.B2(n_992),
.Y(n_1553)
);

NAND2x1p5_ASAP7_75t_L g1554 ( 
.A(n_1333),
.B(n_1352),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1328),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1415),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1417),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1404),
.A2(n_1389),
.B(n_1386),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_SL g1560 ( 
.A1(n_1345),
.A2(n_1369),
.B(n_1259),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1417),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1402),
.A2(n_1275),
.B(n_1278),
.Y(n_1562)
);

OAI222xp33_ASAP7_75t_L g1563 ( 
.A1(n_1412),
.A2(n_1255),
.B1(n_1282),
.B2(n_992),
.C1(n_1342),
.C2(n_932),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1412),
.A2(n_1393),
.B1(n_1406),
.B2(n_992),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1406),
.A2(n_1392),
.B(n_1412),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1412),
.A2(n_1406),
.B1(n_1393),
.B2(n_1392),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1417),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1410),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1417),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1510),
.A2(n_1537),
.B1(n_1553),
.B2(n_1564),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1510),
.A2(n_1537),
.B1(n_1553),
.B2(n_1529),
.Y(n_1571)
);

NOR2x1_ASAP7_75t_SL g1572 ( 
.A(n_1465),
.B(n_1455),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1424),
.A2(n_1517),
.B1(n_1566),
.B2(n_1536),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1462),
.B(n_1439),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1461),
.B(n_1548),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1555),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1441),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_SL g1578 ( 
.A(n_1465),
.B(n_1426),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1513),
.A2(n_1512),
.B(n_1514),
.C(n_1565),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1500),
.A2(n_1432),
.B(n_1460),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1462),
.B(n_1448),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1424),
.A2(n_1436),
.B1(n_1428),
.B2(n_1449),
.Y(n_1582)
);

AOI21x1_ASAP7_75t_SL g1583 ( 
.A1(n_1459),
.A2(n_1545),
.B(n_1485),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1445),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1534),
.A2(n_1471),
.B1(n_1458),
.B2(n_1494),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1480),
.B(n_1465),
.Y(n_1586)
);

AOI21x1_ASAP7_75t_SL g1587 ( 
.A1(n_1476),
.A2(n_1489),
.B(n_1485),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1429),
.B(n_1461),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1519),
.B(n_1531),
.Y(n_1589)
);

O2A1O1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1563),
.A2(n_1436),
.B(n_1508),
.C(n_1560),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1550),
.A2(n_1502),
.B1(n_1438),
.B2(n_1530),
.C(n_1429),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1474),
.A2(n_1552),
.B(n_1547),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1556),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1499),
.A2(n_1498),
.B(n_1450),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1467),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1550),
.A2(n_1438),
.B1(n_1471),
.B2(n_1451),
.Y(n_1597)
);

O2A1O1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1502),
.A2(n_1477),
.B(n_1522),
.C(n_1484),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1550),
.A2(n_1442),
.B1(n_1457),
.B2(n_1539),
.C(n_1481),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1539),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1484),
.A2(n_1497),
.B(n_1457),
.C(n_1488),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1435),
.A2(n_1558),
.B(n_1533),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1468),
.B(n_1473),
.Y(n_1603)
);

AOI21x1_ASAP7_75t_SL g1604 ( 
.A1(n_1476),
.A2(n_1489),
.B(n_1496),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1547),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1494),
.A2(n_1481),
.B(n_1487),
.C(n_1479),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1446),
.A2(n_1472),
.B1(n_1504),
.B2(n_1544),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1472),
.A2(n_1569),
.B1(n_1567),
.B2(n_1561),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1525),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1431),
.A2(n_1523),
.B1(n_1557),
.B2(n_1528),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1435),
.A2(n_1558),
.B(n_1533),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1520),
.B(n_1527),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1568),
.B(n_1542),
.Y(n_1613)
);

AOI21x1_ASAP7_75t_SL g1614 ( 
.A1(n_1491),
.A2(n_1492),
.B(n_1452),
.Y(n_1614)
);

O2A1O1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1535),
.A2(n_1483),
.B(n_1541),
.C(n_1515),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1475),
.A2(n_1425),
.B(n_1559),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1437),
.B(n_1493),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1427),
.B(n_1482),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1453),
.B(n_1490),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1490),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1521),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1487),
.A2(n_1469),
.B1(n_1501),
.B2(n_1552),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1478),
.B(n_1518),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1506),
.A2(n_1562),
.B(n_1549),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1469),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1552),
.A2(n_1486),
.B1(n_1554),
.B2(n_1466),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1518),
.B(n_1443),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1518),
.B(n_1443),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1507),
.A2(n_1540),
.B(n_1546),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1443),
.B(n_1456),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1430),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1453),
.B(n_1495),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1466),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1505),
.B(n_1495),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1505),
.A2(n_1554),
.B(n_1524),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1538),
.B(n_1430),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1470),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1556),
.B(n_1526),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1503),
.B(n_1555),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1526),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1464),
.A2(n_1503),
.B1(n_1532),
.B2(n_1521),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1543),
.A2(n_1440),
.B(n_1433),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1464),
.A2(n_1532),
.B1(n_1463),
.B2(n_1447),
.Y(n_1643)
);

OA22x2_ASAP7_75t_L g1644 ( 
.A1(n_1511),
.A2(n_1564),
.B1(n_1529),
.B2(n_1536),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1551),
.A2(n_1392),
.B(n_1412),
.C(n_1303),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1461),
.B(n_1516),
.Y(n_1646)
);

OA21x2_ASAP7_75t_L g1647 ( 
.A1(n_1500),
.A2(n_1432),
.B(n_1460),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1517),
.A2(n_1392),
.B(n_1412),
.C(n_1303),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1461),
.B(n_1516),
.Y(n_1649)
);

O2A1O1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1517),
.A2(n_1392),
.B(n_1412),
.C(n_1303),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1434),
.Y(n_1651)
);

O2A1O1Ixp5_ASAP7_75t_L g1652 ( 
.A1(n_1545),
.A2(n_1530),
.B(n_1392),
.C(n_1432),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1510),
.A2(n_1553),
.B1(n_1537),
.B2(n_1412),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1429),
.B(n_1461),
.Y(n_1654)
);

O2A1O1Ixp5_ASAP7_75t_L g1655 ( 
.A1(n_1545),
.A2(n_1530),
.B(n_1392),
.C(n_1432),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1429),
.B(n_1461),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1510),
.A2(n_1553),
.B1(n_1537),
.B2(n_1412),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1448),
.B(n_1519),
.Y(n_1658)
);

A2O1A1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1513),
.A2(n_1412),
.B(n_992),
.C(n_1406),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1448),
.B(n_1519),
.Y(n_1660)
);

BUFx4f_ASAP7_75t_L g1661 ( 
.A(n_1430),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1444),
.A2(n_1392),
.B(n_1509),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1500),
.A2(n_1432),
.B(n_1460),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1461),
.B(n_1516),
.Y(n_1664)
);

O2A1O1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1517),
.A2(n_1392),
.B(n_1412),
.C(n_1303),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1448),
.B(n_1519),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1441),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1545),
.B(n_938),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1451),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1638),
.B(n_1593),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1662),
.B(n_1622),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1577),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1632),
.Y(n_1673)
);

AO21x2_ASAP7_75t_L g1674 ( 
.A1(n_1642),
.A2(n_1611),
.B(n_1602),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1584),
.Y(n_1675)
);

AOI33xp33_ASAP7_75t_L g1676 ( 
.A1(n_1648),
.A2(n_1665),
.A3(n_1650),
.B1(n_1591),
.B2(n_1599),
.B3(n_1600),
.Y(n_1676)
);

INVxp33_ASAP7_75t_L g1677 ( 
.A(n_1589),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1622),
.B(n_1590),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1641),
.B(n_1596),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1667),
.B(n_1595),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1573),
.A2(n_1570),
.B1(n_1571),
.B2(n_1653),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1579),
.A2(n_1659),
.B(n_1652),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1595),
.B(n_1580),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1655),
.A2(n_1657),
.B(n_1653),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1651),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1616),
.Y(n_1686)
);

OR2x6_ASAP7_75t_L g1687 ( 
.A(n_1580),
.B(n_1647),
.Y(n_1687)
);

OR2x6_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1663),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_R g1689 ( 
.A(n_1621),
.B(n_1594),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1586),
.B(n_1637),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1610),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1657),
.A2(n_1570),
.B(n_1571),
.Y(n_1692)
);

AOI33xp33_ASAP7_75t_L g1693 ( 
.A1(n_1600),
.A2(n_1615),
.A3(n_1645),
.B1(n_1660),
.B2(n_1658),
.B3(n_1666),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1663),
.B(n_1644),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1623),
.A2(n_1630),
.B(n_1628),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1644),
.B(n_1581),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1610),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1574),
.Y(n_1698)
);

OR2x6_ASAP7_75t_L g1699 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1627),
.B(n_1588),
.Y(n_1700)
);

BUFx6f_ASAP7_75t_L g1701 ( 
.A(n_1634),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1585),
.A2(n_1582),
.B(n_1668),
.Y(n_1702)
);

BUFx2_ASAP7_75t_L g1703 ( 
.A(n_1608),
.Y(n_1703)
);

OR2x6_ASAP7_75t_L g1704 ( 
.A(n_1608),
.B(n_1598),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1588),
.B(n_1656),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1603),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1654),
.B(n_1656),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1613),
.Y(n_1708)
);

AO21x2_ASAP7_75t_L g1709 ( 
.A1(n_1643),
.A2(n_1654),
.B(n_1597),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1607),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1643),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1597),
.A2(n_1582),
.B(n_1587),
.Y(n_1712)
);

AO21x2_ASAP7_75t_L g1713 ( 
.A1(n_1578),
.A2(n_1626),
.B(n_1601),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1624),
.Y(n_1714)
);

AO21x2_ASAP7_75t_L g1715 ( 
.A1(n_1626),
.A2(n_1572),
.B(n_1633),
.Y(n_1715)
);

AO21x2_ASAP7_75t_L g1716 ( 
.A1(n_1624),
.A2(n_1629),
.B(n_1604),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1629),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1618),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1692),
.A2(n_1649),
.B1(n_1575),
.B2(n_1664),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1683),
.B(n_1687),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1672),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1635),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1672),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1700),
.B(n_1705),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1683),
.B(n_1669),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1711),
.B(n_1592),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1686),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1675),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1711),
.B(n_1612),
.Y(n_1729)
);

NOR4xp25_ASAP7_75t_SL g1730 ( 
.A(n_1703),
.B(n_1625),
.C(n_1620),
.D(n_1583),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1700),
.B(n_1646),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1681),
.A2(n_1609),
.B1(n_1661),
.B2(n_1631),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1714),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1715),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1687),
.B(n_1619),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1687),
.B(n_1688),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1715),
.Y(n_1737)
);

CKINVDCx11_ASAP7_75t_R g1738 ( 
.A(n_1673),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1694),
.B(n_1631),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1690),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1680),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1717),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1705),
.B(n_1605),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1694),
.B(n_1631),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1695),
.B(n_1617),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1684),
.A2(n_1636),
.B(n_1661),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1695),
.B(n_1639),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1690),
.B(n_1614),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1745),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1741),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1739),
.B(n_1698),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1738),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1721),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1719),
.A2(n_1702),
.B1(n_1682),
.B2(n_1678),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1724),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1740),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1721),
.Y(n_1757)
);

AOI31xp33_ASAP7_75t_L g1758 ( 
.A1(n_1746),
.A2(n_1670),
.A3(n_1707),
.B(n_1677),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1739),
.B(n_1679),
.Y(n_1759)
);

NOR3xp33_ASAP7_75t_L g1760 ( 
.A(n_1719),
.B(n_1676),
.C(n_1670),
.Y(n_1760)
);

AND2x2_ASAP7_75t_SL g1761 ( 
.A(n_1748),
.B(n_1712),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1723),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1732),
.A2(n_1678),
.B1(n_1671),
.B2(n_1704),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1723),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1746),
.A2(n_1678),
.B1(n_1671),
.B2(n_1704),
.Y(n_1765)
);

AO21x2_ASAP7_75t_L g1766 ( 
.A1(n_1727),
.A2(n_1716),
.B(n_1674),
.Y(n_1766)
);

OAI31xp33_ASAP7_75t_L g1767 ( 
.A1(n_1747),
.A2(n_1710),
.A3(n_1696),
.B(n_1718),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1728),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1724),
.B(n_1708),
.Y(n_1769)
);

AO21x2_ASAP7_75t_L g1770 ( 
.A1(n_1736),
.A2(n_1716),
.B(n_1674),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1738),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1744),
.B(n_1747),
.Y(n_1772)
);

OAI321xp33_ASAP7_75t_L g1773 ( 
.A1(n_1747),
.A2(n_1678),
.A3(n_1699),
.B1(n_1691),
.B2(n_1697),
.C(n_1696),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1731),
.B(n_1718),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1743),
.B(n_1693),
.C(n_1712),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1728),
.Y(n_1776)
);

AO21x2_ASAP7_75t_L g1777 ( 
.A1(n_1736),
.A2(n_1674),
.B(n_1709),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1744),
.B(n_1679),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1748),
.B(n_1685),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1748),
.B(n_1685),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1722),
.A2(n_1712),
.B1(n_1743),
.B2(n_1729),
.C(n_1706),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1748),
.B(n_1701),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1725),
.B(n_1735),
.Y(n_1783)
);

INVx5_ASAP7_75t_L g1784 ( 
.A(n_1722),
.Y(n_1784)
);

NOR2x1_ASAP7_75t_L g1785 ( 
.A(n_1734),
.B(n_1713),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1750),
.Y(n_1786)
);

INVxp67_ASAP7_75t_SL g1787 ( 
.A(n_1750),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1753),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1757),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1762),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1785),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1764),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1768),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1758),
.A2(n_1713),
.B(n_1730),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1771),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1784),
.B(n_1736),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1749),
.B(n_1720),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1773),
.A2(n_1733),
.B(n_1742),
.Y(n_1798)
);

NOR2x1p5_ASAP7_75t_L g1799 ( 
.A(n_1752),
.B(n_1734),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1776),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1761),
.B(n_1720),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1769),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1760),
.B(n_1748),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1766),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1770),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1783),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1783),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1752),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1774),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1755),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1761),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1759),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1808),
.B(n_1771),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1800),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1800),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1812),
.B(n_1767),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1788),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1811),
.B(n_1772),
.Y(n_1818)
);

AOI221x1_ASAP7_75t_L g1819 ( 
.A1(n_1794),
.A2(n_1771),
.B1(n_1775),
.B2(n_1765),
.C(n_1763),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1811),
.B(n_1756),
.Y(n_1820)
);

AND2x2_ASAP7_75t_SL g1821 ( 
.A(n_1798),
.B(n_1754),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1795),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1801),
.B(n_1756),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1810),
.B(n_1759),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1801),
.B(n_1756),
.Y(n_1825)
);

INVx5_ASAP7_75t_L g1826 ( 
.A(n_1791),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1801),
.B(n_1777),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1797),
.B(n_1778),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_SL g1829 ( 
.A(n_1803),
.B(n_1782),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1802),
.B(n_1726),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1788),
.Y(n_1831)
);

BUFx3_ASAP7_75t_L g1832 ( 
.A(n_1795),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1778),
.Y(n_1833)
);

INVx6_ASAP7_75t_L g1834 ( 
.A(n_1799),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1808),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1796),
.B(n_1784),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1798),
.B(n_1782),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1798),
.B(n_1734),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1786),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1789),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1786),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1810),
.B(n_1751),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1789),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1798),
.B(n_1734),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1798),
.B(n_1737),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1795),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1799),
.B(n_1779),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1817),
.Y(n_1848)
);

NAND2x1p5_ASAP7_75t_L g1849 ( 
.A(n_1826),
.B(n_1803),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1840),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1832),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1830),
.B(n_1802),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1840),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1822),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1829),
.B(n_1796),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1819),
.A2(n_1794),
.B(n_1754),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1835),
.B(n_1809),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1835),
.B(n_1846),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1817),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1824),
.B(n_1806),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1846),
.B(n_1813),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1829),
.B(n_1796),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1828),
.B(n_1796),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1824),
.B(n_1806),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1832),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1839),
.B(n_1807),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1832),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1821),
.B(n_1795),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1828),
.B(n_1796),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1828),
.B(n_1796),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1821),
.B(n_1807),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1821),
.B(n_1790),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1822),
.B(n_1792),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1843),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1841),
.B(n_1787),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1833),
.B(n_1787),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1822),
.B(n_1792),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1842),
.B(n_1793),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1833),
.B(n_1791),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1842),
.B(n_1793),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1831),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1826),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1833),
.B(n_1791),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1849),
.Y(n_1884)
);

INVx1_ASAP7_75t_SL g1885 ( 
.A(n_1858),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1848),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1865),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1865),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1867),
.B(n_1818),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1868),
.Y(n_1890)
);

OAI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1849),
.A2(n_1837),
.B(n_1819),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1861),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1848),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1875),
.B(n_1866),
.Y(n_1894)
);

OAI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1856),
.A2(n_1834),
.B1(n_1816),
.B2(n_1837),
.C(n_1827),
.Y(n_1895)
);

AOI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1849),
.A2(n_1709),
.B1(n_1781),
.B2(n_1834),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1855),
.B(n_1847),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1851),
.B(n_1847),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1855),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1859),
.Y(n_1900)
);

BUFx2_ASAP7_75t_L g1901 ( 
.A(n_1854),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1851),
.B(n_1818),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1862),
.B(n_1834),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1859),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1876),
.B(n_1872),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1854),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1862),
.B(n_1876),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1875),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1857),
.B(n_1863),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1881),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1879),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1901),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1895),
.A2(n_1871),
.B(n_1836),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1891),
.A2(n_1837),
.B(n_1838),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1901),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1888),
.B(n_1863),
.Y(n_1916)
);

O2A1O1Ixp33_ASAP7_75t_SL g1917 ( 
.A1(n_1887),
.A2(n_1882),
.B(n_1873),
.C(n_1877),
.Y(n_1917)
);

AOI22x1_ASAP7_75t_L g1918 ( 
.A1(n_1884),
.A2(n_1882),
.B1(n_1771),
.B2(n_1836),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1906),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1906),
.Y(n_1920)
);

NOR3xp33_ASAP7_75t_SL g1921 ( 
.A(n_1889),
.B(n_1576),
.C(n_1850),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1894),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1908),
.B(n_1892),
.Y(n_1923)
);

OAI211xp5_ASAP7_75t_L g1924 ( 
.A1(n_1896),
.A2(n_1826),
.B(n_1827),
.C(n_1838),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1888),
.Y(n_1925)
);

OAI31xp33_ASAP7_75t_L g1926 ( 
.A1(n_1885),
.A2(n_1827),
.A3(n_1845),
.B(n_1844),
.Y(n_1926)
);

NOR2x1_ASAP7_75t_L g1927 ( 
.A(n_1884),
.B(n_1853),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1894),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1886),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1886),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1898),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1907),
.B(n_1869),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1890),
.B(n_1834),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1897),
.A2(n_1911),
.B1(n_1903),
.B2(n_1907),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1931),
.B(n_1899),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1912),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1916),
.B(n_1903),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1915),
.Y(n_1938)
);

INVxp67_ASAP7_75t_SL g1939 ( 
.A(n_1927),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1919),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1934),
.B(n_1898),
.Y(n_1941)
);

OAI31xp33_ASAP7_75t_SL g1942 ( 
.A1(n_1924),
.A2(n_1891),
.A3(n_1897),
.B(n_1898),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1920),
.B(n_1884),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1925),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1916),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1925),
.B(n_1905),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1923),
.B(n_1909),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1939),
.A2(n_1917),
.B(n_1914),
.Y(n_1948)
);

NOR3xp33_ASAP7_75t_L g1949 ( 
.A(n_1939),
.B(n_1933),
.C(n_1913),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1937),
.A2(n_1921),
.B1(n_1933),
.B2(n_1932),
.Y(n_1950)
);

NOR3xp33_ASAP7_75t_L g1951 ( 
.A(n_1941),
.B(n_1928),
.C(n_1922),
.Y(n_1951)
);

NOR3xp33_ASAP7_75t_L g1952 ( 
.A(n_1935),
.B(n_1917),
.C(n_1929),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1945),
.Y(n_1953)
);

OAI211xp5_ASAP7_75t_L g1954 ( 
.A1(n_1942),
.A2(n_1918),
.B(n_1921),
.C(n_1926),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1946),
.A2(n_1896),
.B1(n_1930),
.B2(n_1902),
.C(n_1904),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1946),
.A2(n_1910),
.B1(n_1904),
.B2(n_1900),
.C(n_1893),
.Y(n_1956)
);

AOI221x1_ASAP7_75t_L g1957 ( 
.A1(n_1944),
.A2(n_1910),
.B1(n_1900),
.B2(n_1893),
.C(n_1874),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1945),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1952),
.A2(n_1834),
.B1(n_1947),
.B2(n_1943),
.Y(n_1959)
);

OAI222xp33_ASAP7_75t_L g1960 ( 
.A1(n_1948),
.A2(n_1940),
.B1(n_1938),
.B2(n_1936),
.C1(n_1826),
.C2(n_1943),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1953),
.Y(n_1961)
);

AND3x4_ASAP7_75t_L g1962 ( 
.A(n_1949),
.B(n_1836),
.C(n_1780),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1958),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1954),
.A2(n_1950),
.B1(n_1955),
.B2(n_1951),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1957),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1963),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_SL g1967 ( 
.A(n_1960),
.B(n_1826),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1961),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1959),
.B(n_1826),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1964),
.B(n_1852),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1965),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1962),
.B(n_1869),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1959),
.B(n_1870),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1972),
.A2(n_1956),
.B1(n_1836),
.B2(n_1879),
.Y(n_1974)
);

INVx5_ASAP7_75t_L g1975 ( 
.A(n_1973),
.Y(n_1975)
);

OAI211xp5_ASAP7_75t_L g1976 ( 
.A1(n_1971),
.A2(n_1826),
.B(n_1689),
.C(n_1883),
.Y(n_1976)
);

OAI221xp5_ASAP7_75t_L g1977 ( 
.A1(n_1967),
.A2(n_1881),
.B1(n_1883),
.B2(n_1880),
.C(n_1878),
.Y(n_1977)
);

NAND2xp33_ASAP7_75t_L g1978 ( 
.A(n_1970),
.B(n_1866),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1966),
.B(n_1852),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1975),
.B(n_1969),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1975),
.B(n_1968),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1979),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1982),
.A2(n_1978),
.B1(n_1974),
.B2(n_1977),
.Y(n_1983)
);

OAI322xp33_ASAP7_75t_SL g1984 ( 
.A1(n_1983),
.A2(n_1981),
.A3(n_1980),
.B1(n_1976),
.B2(n_1967),
.C1(n_1814),
.C2(n_1815),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1984),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1984),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1986),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1985),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1987),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1988),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1989),
.A2(n_1870),
.B1(n_1836),
.B2(n_1814),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1991),
.A2(n_1990),
.B1(n_1815),
.B2(n_1820),
.Y(n_1992)
);

NAND2x2_ASAP7_75t_L g1993 ( 
.A(n_1992),
.B(n_1860),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1993),
.B(n_1860),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1820),
.B1(n_1823),
.B2(n_1825),
.Y(n_1995)
);

AOI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1995),
.A2(n_1864),
.B(n_1805),
.C(n_1804),
.Y(n_1996)
);


endmodule