module real_aes_4663_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_235;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_780;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_954;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_968;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g645 ( .A(n_0), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_1), .A2(n_13), .B1(n_159), .B2(n_568), .Y(n_575) );
INVx2_ASAP7_75t_L g555 ( .A(n_2), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_3), .A2(n_33), .B1(n_117), .B2(n_121), .Y(n_116) );
INVx1_ASAP7_75t_SL g611 ( .A(n_4), .Y(n_611) );
INVx1_ASAP7_75t_L g530 ( .A(n_5), .Y(n_530) );
INVx1_ASAP7_75t_L g902 ( .A(n_5), .Y(n_902) );
INVxp67_ASAP7_75t_L g924 ( .A(n_5), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_6), .A2(n_90), .B1(n_197), .B2(n_198), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_7), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_8), .B(n_169), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_9), .A2(n_34), .B1(n_157), .B2(n_158), .Y(n_156) );
INVx2_ASAP7_75t_L g304 ( .A(n_10), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_11), .A2(n_57), .B1(n_164), .B2(n_624), .Y(n_623) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_12), .A2(n_68), .B(n_142), .Y(n_141) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_12), .A2(n_68), .B(n_142), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_14), .B(n_238), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_15), .A2(n_905), .B1(n_906), .B2(n_910), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_15), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_16), .A2(n_81), .B1(n_122), .B2(n_163), .Y(n_550) );
INVx2_ASAP7_75t_L g571 ( .A(n_17), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_18), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_SL g302 ( .A(n_19), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_20), .B(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_21), .A2(n_25), .B1(n_197), .B2(n_198), .Y(n_576) );
BUFx3_ASAP7_75t_L g928 ( .A(n_22), .Y(n_928) );
BUFx8_ASAP7_75t_SL g965 ( .A(n_22), .Y(n_965) );
O2A1O1Ixp5_ASAP7_75t_L g566 ( .A1(n_23), .A2(n_117), .B(n_126), .C(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_24), .A2(n_63), .B1(n_118), .B2(n_553), .Y(n_552) );
O2A1O1Ixp5_ASAP7_75t_L g246 ( .A1(n_26), .A2(n_125), .B(n_247), .C(n_250), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_27), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_28), .B(n_131), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_29), .A2(n_95), .B1(n_943), .B2(n_944), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_29), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_30), .A2(n_82), .B1(n_254), .B2(n_299), .Y(n_629) );
INVx1_ASAP7_75t_L g534 ( .A(n_31), .Y(n_534) );
INVx1_ASAP7_75t_L g563 ( .A(n_32), .Y(n_563) );
AND2x2_ASAP7_75t_L g930 ( .A(n_35), .B(n_931), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_36), .B(n_233), .Y(n_641) );
INVx2_ASAP7_75t_L g569 ( .A(n_37), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_38), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_39), .A2(n_44), .B1(n_130), .B2(n_133), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_40), .A2(n_67), .B1(n_133), .B2(n_180), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_41), .B(n_122), .Y(n_231) );
INVx2_ASAP7_75t_L g173 ( .A(n_42), .Y(n_173) );
INVx2_ASAP7_75t_L g668 ( .A(n_43), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_45), .B(n_131), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_46), .B(n_167), .Y(n_203) );
INVx1_ASAP7_75t_SL g615 ( .A(n_47), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_48), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_49), .A2(n_136), .B(n_299), .C(n_300), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_50), .A2(n_94), .B1(n_908), .B2(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g909 ( .A(n_50), .Y(n_909) );
INVx1_ASAP7_75t_L g278 ( .A(n_51), .Y(n_278) );
INVx1_ASAP7_75t_L g596 ( .A(n_52), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_53), .A2(n_66), .B1(n_939), .B2(n_940), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_53), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_54), .B(n_952), .Y(n_951) );
INVx2_ASAP7_75t_L g257 ( .A(n_55), .Y(n_257) );
INVx1_ASAP7_75t_L g142 ( .A(n_56), .Y(n_142) );
AND2x4_ASAP7_75t_L g145 ( .A(n_58), .B(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g188 ( .A(n_58), .B(n_146), .Y(n_188) );
INVx2_ASAP7_75t_L g182 ( .A(n_59), .Y(n_182) );
INVx1_ASAP7_75t_L g619 ( .A(n_60), .Y(n_619) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_61), .Y(n_127) );
INVx1_ASAP7_75t_SL g251 ( .A(n_62), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_64), .B(n_613), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_65), .Y(n_186) );
INVx1_ASAP7_75t_L g940 ( .A(n_66), .Y(n_940) );
XOR2xp5_ASAP7_75t_L g906 ( .A(n_69), .B(n_907), .Y(n_906) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_70), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_71), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_72), .A2(n_117), .B(n_136), .C(n_185), .Y(n_184) );
OR2x6_ASAP7_75t_L g531 ( .A(n_73), .B(n_532), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_74), .Y(n_264) );
INVx1_ASAP7_75t_L g274 ( .A(n_75), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_76), .B(n_123), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_77), .B(n_157), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g295 ( .A(n_78), .B(n_296), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_79), .A2(n_177), .B(n_179), .C(n_183), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_79), .A2(n_177), .B(n_179), .C(n_183), .Y(n_215) );
INVx1_ASAP7_75t_L g533 ( .A(n_80), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g161 ( .A1(n_83), .A2(n_96), .B1(n_162), .B2(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g931 ( .A(n_84), .Y(n_931) );
INVx1_ASAP7_75t_L g120 ( .A(n_85), .Y(n_120) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
BUFx5_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_86), .B(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_87), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g671 ( .A(n_88), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_89), .Y(n_914) );
INVx1_ASAP7_75t_L g675 ( .A(n_91), .Y(n_675) );
INVx2_ASAP7_75t_L g603 ( .A(n_92), .Y(n_603) );
INVx2_ASAP7_75t_SL g146 ( .A(n_93), .Y(n_146) );
INVx1_ASAP7_75t_L g908 ( .A(n_94), .Y(n_908) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_95), .B(n_242), .Y(n_634) );
INVx1_ASAP7_75t_L g944 ( .A(n_95), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_97), .B(n_149), .Y(n_275) );
INVx1_ASAP7_75t_SL g150 ( .A(n_98), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_99), .B(n_189), .Y(n_260) );
AND2x2_ASAP7_75t_L g168 ( .A(n_100), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_SL g255 ( .A(n_101), .Y(n_255) );
AO32x2_ASAP7_75t_L g573 ( .A1(n_102), .A2(n_194), .A3(n_227), .B1(n_574), .B2(n_577), .Y(n_573) );
AO22x2_ASAP7_75t_L g694 ( .A1(n_102), .A2(n_226), .B1(n_574), .B2(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_918), .B1(n_932), .B2(n_954), .C(n_959), .Y(n_103) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_904), .B(n_911), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_526), .B1(n_535), .B2(n_897), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22xp33_ASAP7_75t_SL g912 ( .A1(n_108), .A2(n_526), .B1(n_538), .B2(n_898), .Y(n_912) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_108), .Y(n_936) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_416), .Y(n_108) );
NAND4xp25_ASAP7_75t_L g109 ( .A(n_110), .B(n_342), .C(n_376), .D(n_385), .Y(n_109) );
O2A1O1Ixp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_204), .B(n_220), .C(n_280), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_151), .Y(n_111) );
INVxp67_ASAP7_75t_L g350 ( .A(n_112), .Y(n_350) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g206 ( .A(n_113), .B(n_207), .Y(n_206) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_113), .B(n_219), .Y(n_365) );
NOR2x1_ASAP7_75t_L g374 ( .A(n_113), .B(n_211), .Y(n_374) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g313 ( .A(n_114), .Y(n_313) );
AOI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_128), .B(n_147), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_125), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_117), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g613 ( .A(n_119), .Y(n_613) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g198 ( .A(n_123), .Y(n_198) );
INVx1_ASAP7_75t_L g296 ( .A(n_123), .Y(n_296) );
INVx1_ASAP7_75t_L g624 ( .A(n_123), .Y(n_624) );
INVx1_ASAP7_75t_L g638 ( .A(n_123), .Y(n_638) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g159 ( .A(n_124), .Y(n_159) );
INVx2_ASAP7_75t_L g181 ( .A(n_124), .Y(n_181) );
INVx6_ASAP7_75t_L g238 ( .A(n_124), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_125), .B(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_125), .B(n_187), .Y(n_598) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_126), .A2(n_240), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_126), .A2(n_637), .B(n_639), .Y(n_636) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g136 ( .A(n_127), .Y(n_136) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_127), .Y(n_183) );
INVxp67_ASAP7_75t_L g200 ( .A(n_127), .Y(n_200) );
INVx4_ASAP7_75t_L g234 ( .A(n_127), .Y(n_234) );
INVx1_ASAP7_75t_L g631 ( .A(n_127), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_135), .B(n_137), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g157 ( .A(n_132), .Y(n_157) );
INVx2_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
INVx1_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
INVx2_ASAP7_75t_L g197 ( .A(n_132), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g293 ( .A(n_132), .B(n_294), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g591 ( .A(n_133), .B(n_592), .Y(n_591) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_133), .A2(n_183), .B(n_671), .C(n_672), .Y(n_670) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_135), .B(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_135), .A2(n_550), .B1(n_551), .B2(n_552), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_135), .B(n_187), .Y(n_593) );
NOR3xp33_ASAP7_75t_L g595 ( .A(n_135), .B(n_187), .C(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_136), .A2(n_157), .B(n_615), .C(n_616), .Y(n_614) );
A2O1A1Ixp33_ASAP7_75t_L g666 ( .A1(n_136), .A2(n_667), .B(n_668), .C(n_669), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
AOI21x1_ASAP7_75t_L g207 ( .A1(n_138), .A2(n_208), .B(n_209), .Y(n_207) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g290 ( .A(n_140), .Y(n_290) );
INVx4_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx3_ASAP7_75t_L g167 ( .A(n_141), .Y(n_167) );
INVx2_ASAP7_75t_L g228 ( .A(n_141), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_143), .A2(n_230), .B(n_235), .Y(n_229) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_144), .A2(n_226), .B(n_275), .Y(n_279) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g165 ( .A(n_145), .B(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
INVx1_ASAP7_75t_L g259 ( .A(n_145), .Y(n_259) );
AND2x2_ASAP7_75t_L g548 ( .A(n_145), .B(n_289), .Y(n_548) );
INVx3_ASAP7_75t_L g608 ( .A(n_145), .Y(n_608) );
AND2x2_ASAP7_75t_L g695 ( .A(n_145), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx3_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
INVx1_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
INVx1_ASAP7_75t_L g578 ( .A(n_149), .Y(n_578) );
INVx1_ASAP7_75t_L g618 ( .A(n_149), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g626 ( .A(n_149), .B(n_608), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_149), .B(n_608), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_149), .B(n_608), .Y(n_673) );
INVx1_ASAP7_75t_L g696 ( .A(n_149), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_151), .A2(n_361), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_151), .Y(n_423) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_170), .Y(n_151) );
INVx1_ASAP7_75t_L g333 ( .A(n_152), .Y(n_333) );
AND2x6_ASAP7_75t_SL g348 ( .A(n_152), .B(n_206), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_152), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_152), .B(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_153), .B(n_191), .Y(n_308) );
AND2x2_ASAP7_75t_L g453 ( .A(n_153), .B(n_171), .Y(n_453) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_SL g219 ( .A(n_154), .Y(n_219) );
AO31x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_160), .A3(n_165), .B(n_168), .Y(n_154) );
INVx1_ASAP7_75t_L g564 ( .A(n_158), .Y(n_564) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g256 ( .A(n_159), .Y(n_256) );
INVxp67_ASAP7_75t_SL g299 ( .A(n_159), .Y(n_299) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g272 ( .A(n_164), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_166), .B(n_194), .Y(n_212) );
AO21x2_ASAP7_75t_L g588 ( .A1(n_166), .A2(n_589), .B(n_602), .Y(n_588) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_167), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g468 ( .A(n_170), .Y(n_468) );
NOR2x1_ASAP7_75t_L g170 ( .A(n_171), .B(n_190), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_171), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g353 ( .A(n_171), .Y(n_353) );
AND2x4_ASAP7_75t_L g379 ( .A(n_171), .B(n_218), .Y(n_379) );
INVx1_ASAP7_75t_L g389 ( .A(n_171), .Y(n_389) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_175), .Y(n_171) );
INVxp67_ASAP7_75t_SL g217 ( .A(n_172), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx1_ASAP7_75t_L g192 ( .A(n_174), .Y(n_192) );
NOR4xp25_ASAP7_75t_L g175 ( .A(n_176), .B(n_184), .C(n_187), .D(n_189), .Y(n_175) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g642 ( .A(n_178), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_182), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_180), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g254 ( .A(n_180), .Y(n_254) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g269 ( .A(n_181), .Y(n_269) );
INVx2_ASAP7_75t_SL g202 ( .A(n_183), .Y(n_202) );
INVx1_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_183), .B(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_183), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g551 ( .A(n_183), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_183), .A2(n_610), .B(n_611), .C(n_612), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_183), .B(n_626), .Y(n_625) );
INVxp67_ASAP7_75t_SL g216 ( .A(n_184), .Y(n_216) );
NOR2x1_ASAP7_75t_SL g287 ( .A(n_187), .B(n_288), .Y(n_287) );
AOI221x1_ASAP7_75t_L g557 ( .A1(n_187), .A2(n_558), .B1(n_560), .B2(n_562), .C(n_564), .Y(n_557) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g332 ( .A(n_191), .B(n_319), .Y(n_332) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_191), .Y(n_341) );
INVx1_ASAP7_75t_L g508 ( .A(n_191), .Y(n_508) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_203), .Y(n_191) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_192), .A2(n_229), .B(n_241), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_199), .B1(n_201), .B2(n_202), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g599 ( .A1(n_197), .A2(n_249), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g610 ( .A(n_198), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g252 ( .A1(n_199), .A2(n_253), .B(n_258), .Y(n_252) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g209 ( .A(n_203), .Y(n_209) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_210), .Y(n_205) );
AND2x2_ASAP7_75t_L g439 ( .A(n_206), .B(n_358), .Y(n_439) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_206), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_206), .B(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g318 ( .A(n_207), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g410 ( .A(n_207), .Y(n_410) );
AND2x2_ASAP7_75t_L g339 ( .A(n_210), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g362 ( .A(n_210), .B(n_350), .Y(n_362) );
AND2x4_ASAP7_75t_L g525 ( .A(n_210), .B(n_378), .Y(n_525) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_218), .Y(n_210) );
AND2x4_ASAP7_75t_L g359 ( .A(n_211), .B(n_319), .Y(n_359) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_211), .Y(n_505) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_217), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g317 ( .A(n_218), .Y(n_317) );
BUFx2_ASAP7_75t_SL g358 ( .A(n_218), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_218), .B(n_410), .Y(n_490) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_220), .A2(n_359), .B1(n_377), .B2(n_380), .C(n_383), .Y(n_376) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_222), .B(n_243), .Y(n_221) );
INVx2_ASAP7_75t_L g382 ( .A(n_222), .Y(n_382) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g395 ( .A(n_223), .B(n_328), .Y(n_395) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_223), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_223), .B(n_261), .Y(n_437) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g356 ( .A(n_224), .B(n_262), .Y(n_356) );
AND2x2_ASAP7_75t_L g399 ( .A(n_224), .B(n_244), .Y(n_399) );
AND2x2_ASAP7_75t_L g474 ( .A(n_224), .B(n_338), .Y(n_474) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_229), .B(n_241), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AO31x2_ASAP7_75t_L g556 ( .A1(n_227), .A2(n_557), .A3(n_565), .B(n_570), .Y(n_556) );
BUFx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g242 ( .A(n_228), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_228), .B(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_228), .B(n_555), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_228), .B(n_571), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g560 ( .A(n_233), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g562 ( .A(n_233), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
O2A1O1Ixp5_ASAP7_75t_SL g263 ( .A1(n_234), .A2(n_264), .B(n_265), .C(n_268), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_234), .B(n_645), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_239), .B(n_240), .Y(n_235) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g249 ( .A(n_238), .Y(n_249) );
INVx1_ASAP7_75t_L g267 ( .A(n_238), .Y(n_267) );
INVx2_ASAP7_75t_L g301 ( .A(n_238), .Y(n_301) );
INVx1_ASAP7_75t_L g553 ( .A(n_238), .Y(n_553) );
INVx2_ASAP7_75t_SL g568 ( .A(n_238), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_240), .A2(n_292), .B(n_295), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_243), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_261), .Y(n_243) );
INVx2_ASAP7_75t_SL g323 ( .A(n_244), .Y(n_323) );
BUFx2_ASAP7_75t_L g502 ( .A(n_244), .Y(n_502) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g284 ( .A(n_245), .Y(n_284) );
INVx3_ASAP7_75t_L g331 ( .A(n_245), .Y(n_331) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_252), .B(n_260), .Y(n_245) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_249), .B(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B1(n_256), .B2(n_257), .Y(n_253) );
AND2x4_ASAP7_75t_L g285 ( .A(n_261), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g460 ( .A(n_261), .B(n_286), .Y(n_460) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g346 ( .A(n_262), .B(n_330), .Y(n_346) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_270), .B(n_279), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_263), .A2(n_270), .B(n_279), .Y(n_325) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_266), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g594 ( .A(n_269), .Y(n_594) );
NAND3x1_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .C(n_276), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OAI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_305), .B(n_314), .C(n_326), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g435 ( .A(n_283), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_283), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g459 ( .A(n_283), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_R g283 ( .A(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g404 ( .A(n_284), .Y(n_404) );
INVx2_ASAP7_75t_L g375 ( .A(n_285), .Y(n_375) );
AND2x2_ASAP7_75t_L g381 ( .A(n_285), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_285), .B(n_404), .Y(n_403) );
OAI322xp33_ASAP7_75t_L g431 ( .A1(n_285), .A2(n_361), .A3(n_432), .B1(n_434), .B2(n_438), .C1(n_440), .C2(n_446), .Y(n_431) );
AND2x2_ASAP7_75t_L g519 ( .A(n_285), .B(n_474), .Y(n_519) );
OR2x2_ASAP7_75t_L g324 ( .A(n_286), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g328 ( .A(n_286), .Y(n_328) );
INVx1_ASAP7_75t_L g336 ( .A(n_286), .Y(n_336) );
AND2x2_ASAP7_75t_L g510 ( .A(n_286), .B(n_325), .Y(n_510) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_286), .Y(n_522) );
AO31x2_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .A3(n_297), .B(n_303), .Y(n_286) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_290), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g559 ( .A(n_301), .Y(n_559) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g409 ( .A(n_312), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_312), .Y(n_415) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_312), .Y(n_514) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g319 ( .A(n_313), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_320), .Y(n_314) );
NOR3xp33_ASAP7_75t_L g347 ( .A(n_315), .B(n_348), .C(n_349), .Y(n_347) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g408 ( .A(n_317), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g478 ( .A(n_317), .Y(n_478) );
INVx2_ASAP7_75t_L g378 ( .A(n_318), .Y(n_378) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
AND2x2_ASAP7_75t_L g524 ( .A(n_322), .B(n_356), .Y(n_524) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g355 ( .A(n_323), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g380 ( .A(n_323), .B(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g430 ( .A(n_323), .B(n_324), .Y(n_430) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_323), .B(n_478), .C(n_505), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_324), .A2(n_419), .B(n_421), .Y(n_418) );
OAI31xp33_ASAP7_75t_L g422 ( .A1(n_324), .A2(n_423), .A3(n_424), .B(n_425), .Y(n_422) );
AOI32xp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_332), .A3(n_333), .B1(n_334), .B2(n_339), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g392 ( .A(n_328), .B(n_338), .Y(n_392) );
INVx1_ASAP7_75t_L g444 ( .A(n_328), .Y(n_444) );
INVx1_ASAP7_75t_L g456 ( .A(n_328), .Y(n_456) );
AND2x2_ASAP7_75t_L g469 ( .A(n_328), .B(n_356), .Y(n_469) );
INVx1_ASAP7_75t_L g473 ( .A(n_328), .Y(n_473) );
OR2x2_ASAP7_75t_L g476 ( .A(n_328), .B(n_442), .Y(n_476) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
INVx1_ASAP7_75t_L g497 ( .A(n_329), .Y(n_497) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g337 ( .A(n_330), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_331), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_331), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g401 ( .A(n_332), .Y(n_401) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g345 ( .A(n_336), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g496 ( .A(n_336), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_337), .Y(n_424) );
AND2x2_ASAP7_75t_L g394 ( .A(n_338), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g405 ( .A(n_339), .Y(n_405) );
INVx1_ASAP7_75t_L g452 ( .A(n_340), .Y(n_452) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g371 ( .A(n_341), .Y(n_371) );
NOR2x1p5_ASAP7_75t_L g428 ( .A(n_341), .B(n_365), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_341), .B(n_359), .Y(n_480) );
NOR2xp33_ASAP7_75t_SL g342 ( .A(n_343), .B(n_363), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B(n_354), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_345), .B(n_357), .Y(n_384) );
AND2x2_ASAP7_75t_L g391 ( .A(n_346), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g455 ( .A(n_346), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_346), .B(n_404), .Y(n_475) );
INVx1_ASAP7_75t_L g425 ( .A(n_348), .Y(n_425) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
NOR2xp33_ASAP7_75t_SL g506 ( .A(n_350), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_352), .B(n_442), .Y(n_445) );
INVx1_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
AND2x2_ASAP7_75t_L g433 ( .A(n_353), .B(n_415), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B1(n_360), .B2(n_362), .Y(n_354) );
OAI21xp5_ASAP7_75t_SL g393 ( .A1(n_355), .A2(n_394), .B(n_396), .Y(n_393) );
INVx2_ASAP7_75t_L g442 ( .A(n_356), .Y(n_442) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B(n_367), .C(n_375), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g467 ( .A(n_365), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g465 ( .A(n_366), .Y(n_465) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_369), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_369), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g463 ( .A(n_373), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_374), .A2(n_465), .B1(n_466), .B2(n_469), .Y(n_464) );
AND2x2_ASAP7_75t_L g488 ( .A(n_374), .B(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_379), .Y(n_396) );
INVx2_ASAP7_75t_SL g402 ( .A(n_379), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_379), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g513 ( .A(n_379), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI211xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_387), .B(n_397), .C(n_406), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_390), .B(n_393), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g413 ( .A(n_392), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_395), .A2(n_524), .B(n_525), .Y(n_523) );
OAI22xp33_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_400), .B1(n_403), .B2(n_405), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g420 ( .A(n_399), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_399), .B(n_516), .Y(n_515) );
NAND2x1_ASAP7_75t_SL g521 ( .A(n_399), .B(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_411), .B1(n_413), .B2(n_414), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g483 ( .A(n_409), .Y(n_483) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_413), .B(n_462), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_448), .C(n_491), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_422), .B1(n_426), .B2(n_429), .C(n_431), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_421), .A2(n_482), .B1(n_484), .B2(n_485), .C(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g493 ( .A(n_426), .Y(n_493) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_428), .Y(n_518) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g462 ( .A(n_436), .Y(n_462) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_439), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_445), .Y(n_440) );
INVx2_ASAP7_75t_SL g484 ( .A(n_441), .Y(n_484) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_470), .C(n_481), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_454), .B(n_457), .C(n_464), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g516 ( .A(n_456), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .B(n_463), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI31xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_475), .A3(n_476), .B(n_477), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_471), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_478), .Y(n_500) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g494 ( .A(n_488), .Y(n_494) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI211xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_495), .B(n_498), .C(n_511), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_501), .B(n_503), .C(n_509), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI211xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_515), .B(n_517), .C(n_523), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
INVx4_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx8_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
OR2x6_ASAP7_75t_L g917 ( .A(n_530), .B(n_531), .Y(n_917) );
INVx8_ASAP7_75t_L g903 ( .A(n_531), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_791), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_689), .C(n_743), .Y(n_539) );
AOI211xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_583), .B(n_657), .C(n_687), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_579), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_572), .Y(n_543) );
AND2x4_ASAP7_75t_L g749 ( .A(n_544), .B(n_713), .Y(n_749) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g692 ( .A(n_545), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_556), .Y(n_545) );
OR2x2_ASAP7_75t_L g581 ( .A(n_546), .B(n_556), .Y(n_581) );
AND2x2_ASAP7_75t_L g742 ( .A(n_546), .B(n_694), .Y(n_742) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g662 ( .A(n_547), .Y(n_662) );
INVx1_ASAP7_75t_L g718 ( .A(n_547), .Y(n_718) );
AOI21x1_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B(n_554), .Y(n_547) );
INVx1_ASAP7_75t_L g667 ( .A(n_553), .Y(n_667) );
INVx1_ASAP7_75t_L g676 ( .A(n_556), .Y(n_676) );
INVx2_ASAP7_75t_L g682 ( .A(n_556), .Y(n_682) );
AND2x2_ASAP7_75t_L g703 ( .A(n_556), .B(n_697), .Y(n_703) );
AND2x2_ASAP7_75t_L g712 ( .A(n_556), .B(n_664), .Y(n_712) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g582 ( .A(n_572), .Y(n_582) );
AND2x2_ASAP7_75t_L g702 ( .A(n_572), .B(n_703), .Y(n_702) );
OR2x2_ASAP7_75t_L g736 ( .A(n_572), .B(n_737), .Y(n_736) );
AND2x4_ASAP7_75t_L g814 ( .A(n_572), .B(n_717), .Y(n_814) );
AND2x2_ASAP7_75t_L g867 ( .A(n_572), .B(n_712), .Y(n_867) );
AND2x2_ASAP7_75t_SL g883 ( .A(n_572), .B(n_663), .Y(n_883) );
BUFx3_ASAP7_75t_L g893 ( .A(n_572), .Y(n_893) );
BUFx8_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g680 ( .A(n_573), .Y(n_680) );
AND2x2_ASAP7_75t_L g783 ( .A(n_573), .B(n_784), .Y(n_783) );
INVxp67_ASAP7_75t_L g656 ( .A(n_577), .Y(n_656) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_578), .B(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND3xp33_ASAP7_75t_SL g878 ( .A(n_580), .B(n_879), .C(n_882), .Y(n_878) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g757 ( .A(n_581), .Y(n_757) );
NAND2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_647), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_584), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_620), .Y(n_585) );
INVx1_ASAP7_75t_L g704 ( .A(n_586), .Y(n_704) );
AND2x2_ASAP7_75t_L g834 ( .A(n_586), .B(n_835), .Y(n_834) );
AND2x2_ASAP7_75t_L g872 ( .A(n_586), .B(n_725), .Y(n_872) );
AND2x4_ASAP7_75t_L g586 ( .A(n_587), .B(n_604), .Y(n_586) );
OR2x2_ASAP7_75t_L g739 ( .A(n_587), .B(n_654), .Y(n_739) );
AND2x2_ASAP7_75t_L g826 ( .A(n_587), .B(n_700), .Y(n_826) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g727 ( .A(n_588), .B(n_686), .Y(n_727) );
BUFx2_ASAP7_75t_L g731 ( .A(n_588), .Y(n_731) );
OR2x2_ASAP7_75t_L g748 ( .A(n_588), .B(n_606), .Y(n_748) );
AO21x2_ASAP7_75t_L g655 ( .A1(n_589), .A2(n_602), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_597), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .B1(n_594), .B2(n_595), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g778 ( .A(n_605), .B(n_633), .Y(n_778) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g652 ( .A(n_606), .Y(n_652) );
INVx2_ASAP7_75t_L g686 ( .A(n_606), .Y(n_686) );
AND2x2_ASAP7_75t_L g759 ( .A(n_606), .B(n_655), .Y(n_759) );
INVx1_ASAP7_75t_L g811 ( .A(n_606), .Y(n_811) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_606), .Y(n_845) );
AO31x2_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .A3(n_614), .B(n_617), .Y(n_606) );
NOR2xp33_ASAP7_75t_SL g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_618), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_620), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g763 ( .A(n_620), .B(n_759), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_620), .B(n_731), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_620), .B(n_730), .Y(n_894) );
NAND2xp67_ASAP7_75t_L g895 ( .A(n_620), .B(n_896), .Y(n_895) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_632), .Y(n_620) );
INVx1_ASAP7_75t_L g650 ( .A(n_621), .Y(n_650) );
INVx2_ASAP7_75t_L g700 ( .A(n_621), .Y(n_700) );
INVx1_ASAP7_75t_L g708 ( .A(n_621), .Y(n_708) );
AND2x2_ASAP7_75t_L g770 ( .A(n_621), .B(n_633), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g621 ( .A(n_622), .B(n_628), .Y(n_621) );
AND2x2_ASAP7_75t_SL g807 ( .A(n_622), .B(n_628), .Y(n_807) );
OA21x2_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B(n_627), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_626), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
OR2x2_ASAP7_75t_L g710 ( .A(n_632), .B(n_655), .Y(n_710) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g654 ( .A(n_633), .Y(n_654) );
INVx1_ASAP7_75t_L g734 ( .A(n_633), .Y(n_734) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_633), .Y(n_802) );
AND2x4_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_640), .B(n_646), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_643), .Y(n_640) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_648), .A2(n_840), .B1(n_842), .B2(n_844), .Y(n_839) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
BUFx3_ASAP7_75t_L g754 ( .A(n_650), .Y(n_754) );
AND2x2_ASAP7_75t_L g801 ( .A(n_651), .B(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
AND2x2_ASAP7_75t_L g810 ( .A(n_654), .B(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g699 ( .A(n_655), .B(n_700), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_677), .B(n_683), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_658), .A2(n_780), .B(n_781), .Y(n_779) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
AND2x4_ASAP7_75t_L g678 ( .A(n_660), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_660), .B(n_693), .Y(n_812) );
INVx4_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g768 ( .A(n_661), .B(n_663), .Y(n_768) );
INVx2_ASAP7_75t_L g819 ( .A(n_661), .Y(n_819) );
NAND2xp5_ASAP7_75t_SL g873 ( .A(n_661), .B(n_703), .Y(n_873) );
BUFx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g784 ( .A(n_662), .Y(n_784) );
INVx2_ASAP7_75t_L g688 ( .A(n_663), .Y(n_688) );
INVx2_ASAP7_75t_L g737 ( .A(n_663), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_663), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_663), .B(n_727), .Y(n_830) );
AND2x4_ASAP7_75t_L g663 ( .A(n_664), .B(n_676), .Y(n_663) );
INVx2_ASAP7_75t_L g697 ( .A(n_664), .Y(n_697) );
INVx1_ASAP7_75t_L g720 ( .A(n_664), .Y(n_720) );
BUFx3_ASAP7_75t_L g751 ( .A(n_664), .Y(n_751) );
AND2x4_ASAP7_75t_L g821 ( .A(n_664), .B(n_680), .Y(n_821) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AO31x2_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .A3(n_673), .B(n_674), .Y(n_665) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g767 ( .A(n_679), .Y(n_767) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_680), .B(n_784), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_681), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g717 ( .A(n_682), .B(n_718), .Y(n_717) );
BUFx3_ASAP7_75t_L g761 ( .A(n_682), .Y(n_761) );
INVx1_ASAP7_75t_L g843 ( .A(n_682), .Y(n_843) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g773 ( .A(n_685), .B(n_739), .Y(n_773) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g789 ( .A(n_686), .B(n_776), .Y(n_789) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_686), .Y(n_889) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_705), .C(n_714), .Y(n_689) );
OAI22xp33_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_698), .B1(n_701), .B2(n_704), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx2_ASAP7_75t_L g864 ( .A(n_692), .Y(n_864) );
AND2x4_ASAP7_75t_L g756 ( .A(n_693), .B(n_757), .Y(n_756) );
INVx4_ASAP7_75t_L g772 ( .A(n_693), .Y(n_772) );
AND2x4_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g713 ( .A(n_694), .Y(n_713) );
INVx1_ASAP7_75t_L g721 ( .A(n_694), .Y(n_721) );
AND2x4_ASAP7_75t_L g750 ( .A(n_694), .B(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g762 ( .A(n_697), .B(n_718), .Y(n_762) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g809 ( .A(n_699), .B(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g862 ( .A(n_699), .B(n_778), .Y(n_862) );
BUFx2_ASAP7_75t_L g725 ( .A(n_700), .Y(n_725) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_700), .Y(n_851) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR2x1_ASAP7_75t_L g715 ( .A(n_702), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g782 ( .A(n_703), .B(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g822 ( .A(n_703), .B(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g857 ( .A(n_703), .B(n_776), .Y(n_857) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_711), .Y(n_705) );
INVx3_ASAP7_75t_L g780 ( .A(n_706), .Y(n_780) );
AND2x4_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
AND2x2_ASAP7_75t_L g804 ( .A(n_707), .B(n_759), .Y(n_804) );
INVx1_ASAP7_75t_L g886 ( .A(n_707), .Y(n_886) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g777 ( .A(n_708), .B(n_778), .Y(n_777) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g787 ( .A(n_710), .Y(n_787) );
INVxp67_ASAP7_75t_SL g852 ( .A(n_710), .Y(n_852) );
OR2x6_ASAP7_75t_L g888 ( .A(n_710), .B(n_889), .Y(n_888) );
OAI31xp33_ASAP7_75t_L g803 ( .A1(n_711), .A2(n_723), .A3(n_804), .B(n_805), .Y(n_803) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx2_ASAP7_75t_L g798 ( .A(n_712), .Y(n_798) );
INVx2_ASAP7_75t_L g881 ( .A(n_712), .Y(n_881) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_722), .B(n_728), .Y(n_714) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_717), .Y(n_891) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_718), .Y(n_753) );
INVx2_ASAP7_75t_L g776 ( .A(n_718), .Y(n_776) );
AOI33xp33_ASAP7_75t_L g771 ( .A1(n_719), .A2(n_772), .A3(n_773), .B1(n_774), .B2(n_775), .B3(n_777), .Y(n_771) );
AND2x2_ASAP7_75t_L g838 ( .A(n_719), .B(n_776), .Y(n_838) );
AND2x2_ASAP7_75t_L g840 ( .A(n_719), .B(n_841), .Y(n_840) );
AND2x4_ASAP7_75t_SL g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
NOR2x1p5_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g758 ( .A(n_725), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x4_ASAP7_75t_L g752 ( .A(n_727), .B(n_753), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g815 ( .A(n_727), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g876 ( .A(n_727), .B(n_770), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_735), .B1(n_738), .B2(n_740), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g796 ( .A(n_731), .B(n_770), .Y(n_796) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_733), .B(n_754), .Y(n_828) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g835 ( .A(n_734), .B(n_807), .Y(n_835) );
AND2x2_ASAP7_75t_L g869 ( .A(n_734), .B(n_807), .Y(n_869) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR2xp67_ASAP7_75t_SL g805 ( .A(n_739), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVxp67_ASAP7_75t_L g829 ( .A(n_742), .Y(n_829) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_764), .C(n_779), .Y(n_743) );
OAI21xp5_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_754), .B(n_755), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_749), .B1(n_750), .B2(n_752), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g896 ( .A(n_748), .Y(n_896) );
INVx2_ASAP7_75t_L g847 ( .A(n_750), .Y(n_847) );
INVx1_ASAP7_75t_L g880 ( .A(n_753), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_758), .B1(n_760), .B2(n_763), .Y(n_755) );
AND2x2_ASAP7_75t_L g769 ( .A(n_759), .B(n_770), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g874 ( .A1(n_760), .A2(n_875), .B(n_876), .Y(n_874) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_771), .Y(n_764) );
OAI21xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B(n_769), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g790 ( .A(n_770), .Y(n_790) );
AND2x2_ASAP7_75t_L g844 ( .A(n_770), .B(n_845), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g788 ( .A(n_772), .B(n_789), .C(n_790), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_772), .A2(n_833), .B1(n_836), .B2(n_837), .C(n_839), .Y(n_832) );
INVx2_ASAP7_75t_L g794 ( .A(n_774), .Y(n_794) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g841 ( .A(n_776), .Y(n_841) );
BUFx3_ASAP7_75t_L g866 ( .A(n_776), .Y(n_866) );
AND2x2_ASAP7_75t_L g875 ( .A(n_778), .B(n_826), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_785), .B(n_788), .Y(n_781) );
AND2x4_ASAP7_75t_SL g842 ( .A(n_783), .B(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g849 ( .A(n_789), .Y(n_849) );
NAND4xp25_ASAP7_75t_L g791 ( .A(n_792), .B(n_831), .C(n_859), .D(n_877), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_808), .Y(n_792) );
OAI221xp5_ASAP7_75t_SL g793 ( .A1(n_794), .A2(n_795), .B1(n_797), .B2(n_800), .C(n_803), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g823 ( .A(n_799), .Y(n_823) );
INVx1_ASAP7_75t_L g854 ( .A(n_799), .Y(n_854) );
INVxp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g825 ( .A(n_802), .Y(n_825) );
INVx1_ASAP7_75t_SL g836 ( .A(n_804), .Y(n_836) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g816 ( .A(n_807), .Y(n_816) );
OAI221xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_812), .B1(n_813), .B2(n_815), .C(n_817), .Y(n_808) );
AND2x2_ASAP7_75t_L g868 ( .A(n_811), .B(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g858 ( .A(n_815), .Y(n_858) );
O2A1O1Ixp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_822), .B(n_824), .C(n_827), .Y(n_817) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AND2x4_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B(n_830), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_846), .Y(n_831) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
OAI21xp33_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B(n_853), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
AND2x4_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_857), .B2(n_858), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_863), .B1(n_865), .B2(n_868), .C(n_870), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
AND2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_873), .B(n_874), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_884), .B1(n_890), .B2(n_892), .Y(n_877) );
OR2x2_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
AND2x4_ASAP7_75t_L g884 ( .A(n_885), .B(n_887), .Y(n_884) );
INVxp67_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVxp67_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
OAI21xp33_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .B(n_895), .Y(n_892) );
BUFx3_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
BUFx12f_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
CKINVDCx11_ASAP7_75t_R g899 ( .A(n_900), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OR2x6_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_903), .B(n_924), .Y(n_923) );
AOI21xp33_ASAP7_75t_L g911 ( .A1(n_904), .A2(n_912), .B(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
BUFx3_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
BUFx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
BUFx3_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
OR2x2_ASAP7_75t_L g920 ( .A(n_921), .B(n_925), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_922), .Y(n_921) );
BUFx12f_ASAP7_75t_L g950 ( .A(n_922), .Y(n_950) );
BUFx8_ASAP7_75t_L g953 ( .A(n_922), .Y(n_953) );
BUFx6f_ASAP7_75t_L g968 ( .A(n_922), .Y(n_968) );
BUFx6f_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_929), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_928), .Y(n_927) );
CKINVDCx6p67_ASAP7_75t_R g958 ( .A(n_928), .Y(n_958) );
OR2x2_ASAP7_75t_SL g956 ( .A(n_929), .B(n_957), .Y(n_956) );
CKINVDCx16_ASAP7_75t_R g929 ( .A(n_930), .Y(n_929) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_930), .A2(n_964), .B(n_966), .Y(n_963) );
NAND2xp5_ASAP7_75t_SL g932 ( .A(n_933), .B(n_951), .Y(n_932) );
INVxp67_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
AOI221x1_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_937), .B1(n_946), .B2(n_947), .C(n_948), .Y(n_934) );
INVx1_ASAP7_75t_L g947 ( .A(n_935), .Y(n_947) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g946 ( .A(n_937), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_941), .B1(n_942), .B2(n_945), .Y(n_937) );
INVx1_ASAP7_75t_L g945 ( .A(n_938), .Y(n_945) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_942), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_944), .B(n_960), .Y(n_959) );
BUFx3_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx3_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_SL g954 ( .A(n_955), .Y(n_954) );
BUFx3_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_961), .Y(n_960) );
BUFx6f_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
CKINVDCx8_ASAP7_75t_R g962 ( .A(n_963), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx5_ASAP7_75t_SL g967 ( .A(n_968), .Y(n_967) );
endmodule