module fake_jpeg_16740_n_361 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_361);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_361;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVxp33_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_19),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_56),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_0),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_48),
.A2(n_33),
.B(n_8),
.C(n_9),
.Y(n_111)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_53),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_1),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_14),
.B(n_1),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_62),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_58),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_64),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_1),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_22),
.B(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_2),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_68),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_70),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_27),
.B1(n_36),
.B2(n_32),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_73),
.A2(n_76),
.B1(n_81),
.B2(n_86),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_25),
.B1(n_36),
.B2(n_18),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_62),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_85),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_36),
.B1(n_32),
.B2(n_25),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_78),
.A2(n_73),
.B1(n_71),
.B2(n_86),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_83),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_29),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_60),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_84),
.A2(n_99),
.B1(n_103),
.B2(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_44),
.B(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_115),
.B1(n_12),
.B2(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_89),
.B(n_94),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_90),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_33),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_33),
.C(n_24),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_95),
.B(n_94),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_46),
.A2(n_30),
.B1(n_28),
.B2(n_23),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_28),
.B1(n_23),
.B2(n_4),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_33),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_113),
.B(n_75),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_118),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_70),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_111),
.A2(n_75),
.B(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_7),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_44),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_40),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_52),
.A2(n_11),
.B1(n_12),
.B2(n_63),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_121),
.A2(n_77),
.B1(n_115),
.B2(n_126),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_12),
.B1(n_58),
.B2(n_76),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_122),
.A2(n_137),
.B1(n_147),
.B2(n_163),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_123),
.Y(n_186)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_126),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_127),
.Y(n_188)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_130),
.Y(n_185)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_132),
.B(n_135),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_77),
.A2(n_88),
.B1(n_115),
.B2(n_79),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_140),
.B(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_158),
.Y(n_171)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_100),
.B1(n_111),
.B2(n_113),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_82),
.B(n_72),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_150),
.B(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_87),
.B(n_101),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_153),
.B1(n_161),
.B2(n_143),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_80),
.A2(n_116),
.B1(n_106),
.B2(n_100),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_93),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_156),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_128),
.C(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_87),
.B(n_101),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_85),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_160),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_71),
.B(n_96),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_126),
.B1(n_139),
.B2(n_141),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_73),
.A2(n_89),
.B1(n_107),
.B2(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_96),
.B(n_104),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_167),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_75),
.B(n_95),
.Y(n_169)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_169),
.A2(n_171),
.B(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_97),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_172),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_97),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_102),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_173),
.B(n_175),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_176),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_102),
.Y(n_175)
);

OAI22x1_ASAP7_75t_SL g180 ( 
.A1(n_148),
.A2(n_80),
.B1(n_157),
.B2(n_163),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_189),
.B1(n_171),
.B2(n_191),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_182),
.A2(n_189),
.B1(n_194),
.B2(n_196),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_147),
.B(n_121),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_136),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_191),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_136),
.B(n_131),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_133),
.A2(n_166),
.B1(n_137),
.B2(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_144),
.B(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_197),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_132),
.A2(n_167),
.B1(n_125),
.B2(n_129),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_123),
.B(n_134),
.C(n_161),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_152),
.B1(n_130),
.B2(n_140),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_168),
.B1(n_208),
.B2(n_198),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_127),
.A2(n_155),
.B(n_149),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_124),
.B(n_120),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_209),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_124),
.B(n_120),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_192),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_210),
.A2(n_211),
.B(n_238),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_215),
.Y(n_249)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_199),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_216),
.A2(n_227),
.B1(n_240),
.B2(n_200),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_237),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_180),
.B1(n_171),
.B2(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_230),
.A2(n_218),
.B1(n_213),
.B2(n_239),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_232),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_174),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_235),
.Y(n_273)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_169),
.A2(n_189),
.B(n_179),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_241),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_189),
.A2(n_180),
.B1(n_194),
.B2(n_177),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_202),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_181),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_245),
.B(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_170),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_202),
.B(n_179),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_181),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_188),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_175),
.B1(n_183),
.B2(n_172),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_247),
.A2(n_253),
.B1(n_267),
.B2(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_197),
.C(n_183),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_260),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_210),
.A2(n_174),
.B1(n_208),
.B2(n_203),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_271),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_238),
.B(n_216),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_256),
.A2(n_262),
.B(n_264),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_188),
.B(n_207),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_190),
.Y(n_263)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_178),
.B(n_190),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_230),
.B1(n_212),
.B2(n_217),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_200),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_231),
.A2(n_237),
.B(n_220),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_272),
.B(n_274),
.Y(n_283)
);

AOI221xp5_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_240),
.B1(n_229),
.B2(n_222),
.C(n_242),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_228),
.A2(n_234),
.B(n_226),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_229),
.A2(n_234),
.B1(n_235),
.B2(n_224),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_222),
.A3(n_221),
.B1(n_236),
.B2(n_211),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_296),
.Y(n_303)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_257),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_285),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_213),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_214),
.B1(n_219),
.B2(n_215),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_292),
.B1(n_297),
.B2(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_249),
.B(n_241),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_211),
.B1(n_250),
.B2(n_256),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_265),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_265),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

OAI322xp33_ASAP7_75t_L g300 ( 
.A1(n_249),
.A2(n_258),
.A3(n_260),
.B1(n_276),
.B2(n_274),
.C1(n_252),
.C2(n_254),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_255),
.C(n_272),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_252),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_251),
.B(n_247),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_302),
.A2(n_297),
.B(n_291),
.C(n_289),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_248),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_251),
.A3(n_250),
.B1(n_254),
.B2(n_253),
.C1(n_270),
.C2(n_255),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_283),
.Y(n_327)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_284),
.A2(n_266),
.B1(n_248),
.B2(n_262),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_312),
.B1(n_284),
.B2(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_281),
.A2(n_259),
.B1(n_261),
.B2(n_269),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_321),
.A2(n_306),
.B1(n_278),
.B2(n_296),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_303),
.A2(n_319),
.B1(n_314),
.B2(n_316),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_322),
.A2(n_324),
.B1(n_329),
.B2(n_308),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_288),
.B1(n_281),
.B2(n_279),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_287),
.C(n_283),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_331),
.C(n_332),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_312),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_316),
.B1(n_319),
.B2(n_308),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_279),
.B1(n_287),
.B2(n_282),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_311),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_301),
.C(n_282),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_261),
.C(n_294),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_324),
.B(n_318),
.Y(n_333)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_333),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_320),
.A2(n_302),
.B(n_309),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_340),
.B(n_341),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_342),
.B1(n_321),
.B2(n_322),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_317),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_339),
.A2(n_315),
.B(n_307),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_326),
.B(n_318),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_325),
.B(n_277),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_332),
.B1(n_331),
.B2(n_321),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_347),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_346),
.B(n_336),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_336),
.A2(n_323),
.B1(n_321),
.B2(n_307),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_349),
.B(n_342),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_354),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_333),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_341),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_352),
.C(n_346),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_350),
.B(n_345),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_359),
.A2(n_350),
.B(n_357),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_347),
.Y(n_361)
);


endmodule