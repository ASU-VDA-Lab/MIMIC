module fake_jpeg_3842_n_310 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_45),
.B(n_51),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_60),
.Y(n_73)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_56),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_25),
.B(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_19),
.B1(n_40),
.B2(n_35),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_64),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_67),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_30),
.B(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_30),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_74),
.Y(n_115)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_19),
.B1(n_41),
.B2(n_43),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_79),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_96),
.B1(n_101),
.B2(n_103),
.Y(n_117)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_19),
.B1(n_34),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_84),
.A2(n_95),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_35),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_5),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_37),
.B1(n_33),
.B2(n_42),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_91),
.B1(n_23),
.B2(n_31),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_40),
.B1(n_42),
.B2(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_33),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_94),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_25),
.B1(n_32),
.B2(n_28),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_32),
.B1(n_27),
.B2(n_26),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_38),
.B1(n_27),
.B2(n_26),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_10),
.B1(n_15),
.B2(n_2),
.Y(n_116)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_104),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_24),
.B1(n_22),
.B2(n_31),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_4),
.Y(n_124)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_38),
.B1(n_24),
.B2(n_22),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_114),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_116),
.A2(n_118),
.B1(n_134),
.B2(n_146),
.Y(n_176)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_120),
.Y(n_165)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_75),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_139),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_5),
.Y(n_129)
);

OR2x4_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_5),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_86),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_16),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_141),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_90),
.B(n_11),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_12),
.Y(n_141)
);

BUFx4f_ASAP7_75t_SL g143 ( 
.A(n_69),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_73),
.B(n_15),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_70),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_108),
.A2(n_13),
.B1(n_14),
.B2(n_104),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_81),
.A2(n_13),
.B1(n_76),
.B2(n_107),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_83),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2x1_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_91),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_168),
.B(n_132),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_81),
.B1(n_90),
.B2(n_105),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_159),
.B1(n_161),
.B2(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_158),
.B(n_138),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_89),
.B1(n_73),
.B2(n_77),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_160),
.B(n_135),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_92),
.B1(n_71),
.B2(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_92),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_102),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_129),
.B(n_80),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_178),
.Y(n_205)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_134),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_131),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_71),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_117),
.A2(n_125),
.B1(n_148),
.B2(n_135),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_119),
.B(n_124),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_196),
.B(n_208),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_131),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_149),
.C(n_151),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_191),
.Y(n_228)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_193),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_122),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_198),
.B(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_150),
.B(n_97),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_158),
.B1(n_155),
.B2(n_152),
.Y(n_214)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_85),
.B(n_125),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_210),
.B(n_212),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_155),
.A2(n_127),
.B(n_142),
.C(n_133),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_112),
.B(n_147),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_214),
.B(n_206),
.Y(n_242)
);

NOR4xp25_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_154),
.C(n_167),
.D(n_171),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_224),
.B(n_204),
.C(n_210),
.D(n_192),
.Y(n_239)
);

AO22x2_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_182),
.B1(n_149),
.B2(n_176),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_218),
.A2(n_186),
.B1(n_211),
.B2(n_183),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_221),
.C(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_199),
.C(n_202),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_154),
.B(n_181),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_225),
.B(n_184),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_154),
.B(n_182),
.C(n_177),
.D(n_171),
.Y(n_224)
);

AOI21x1_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_69),
.B(n_114),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_175),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_229),
.C(n_234),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_175),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_178),
.C(n_166),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_190),
.A2(n_120),
.B1(n_142),
.B2(n_172),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_210),
.B1(n_188),
.B2(n_211),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_195),
.B(n_82),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_195),
.C(n_198),
.Y(n_244)
);

OA21x2_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_223),
.B(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_242),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_190),
.B1(n_200),
.B2(n_187),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_248),
.B1(n_236),
.B2(n_219),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_254),
.C(n_221),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_253),
.B1(n_256),
.B2(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_186),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_207),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_183),
.C(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_205),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_237),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_264),
.C(n_267),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_244),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_232),
.B1(n_256),
.B2(n_255),
.Y(n_281)
);

NAND4xp25_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_239),
.C(n_224),
.D(n_246),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_252),
.B(n_230),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_226),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_230),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_220),
.C(n_234),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_278),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_274),
.Y(n_284)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_218),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_280),
.B(n_281),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_256),
.B1(n_245),
.B2(n_218),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_281),
.B1(n_275),
.B2(n_278),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_248),
.Y(n_278)
);

NAND4xp25_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_251),
.C(n_258),
.D(n_254),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_233),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_280),
.B(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_235),
.B1(n_231),
.B2(n_203),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_273),
.A2(n_240),
.B1(n_258),
.B2(n_247),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_197),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_289),
.B(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_197),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_257),
.C(n_264),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_269),
.C(n_267),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_276),
.A3(n_271),
.B1(n_279),
.B2(n_268),
.C1(n_282),
.C2(n_235),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_297),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_284),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_SL g302 ( 
.A1(n_295),
.A2(n_298),
.B(n_283),
.C(n_285),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_213),
.A3(n_191),
.B1(n_207),
.B2(n_82),
.C1(n_114),
.C2(n_100),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_191),
.C(n_79),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_300),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_288),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_302),
.A2(n_296),
.B(n_289),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_298),
.B1(n_288),
.B2(n_284),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_305),
.A3(n_301),
.B1(n_303),
.B2(n_291),
.C1(n_213),
.C2(n_114),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_308),
.CI(n_284),
.CON(n_309),
.SN(n_309)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_213),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_296),
.Y(n_310)
);


endmodule