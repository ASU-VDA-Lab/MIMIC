module fake_jpeg_12565_n_297 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_155;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g145 ( 
.A(n_52),
.Y(n_145)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_60),
.Y(n_134)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_22),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g99 ( 
.A(n_62),
.Y(n_99)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_72),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_82),
.Y(n_98)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_25),
.A2(n_2),
.B(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_30),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_29),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_32),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_80),
.Y(n_124)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_14),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g106 ( 
.A(n_83),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_6),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_24),
.B(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_26),
.B(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_90),
.Y(n_109)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_89),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_8),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_25),
.Y(n_116)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_94),
.B(n_95),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_40),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_46),
.B1(n_37),
.B2(n_38),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_112),
.B1(n_126),
.B2(n_51),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_46),
.B1(n_37),
.B2(n_38),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_118),
.B1(n_122),
.B2(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_49),
.A2(n_32),
.B1(n_39),
.B2(n_35),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_103),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_35),
.B1(n_39),
.B2(n_43),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_62),
.A2(n_87),
.B1(n_91),
.B2(n_90),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_50),
.A2(n_43),
.B1(n_41),
.B2(n_11),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_70),
.A2(n_41),
.B1(n_9),
.B2(n_8),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_140),
.B1(n_69),
.B2(n_54),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_55),
.A2(n_9),
.B1(n_16),
.B2(n_66),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_67),
.A2(n_92),
.B1(n_81),
.B2(n_75),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_95),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_57),
.B(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_59),
.B(n_76),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_134),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_148),
.A2(n_155),
.B1(n_157),
.B2(n_160),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_73),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_149),
.B(n_150),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_64),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_153),
.B(n_156),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_108),
.A2(n_52),
.B1(n_118),
.B2(n_126),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_121),
.B1(n_127),
.B2(n_146),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_99),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_165),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_127),
.B1(n_121),
.B2(n_146),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_110),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_104),
.B(n_109),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_110),
.B1(n_137),
.B2(n_102),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_106),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_167),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_100),
.A2(n_125),
.B1(n_119),
.B2(n_101),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_170),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_178),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_173),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_120),
.A2(n_139),
.B1(n_114),
.B2(n_123),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_182),
.B(n_167),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_182),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_119),
.A2(n_125),
.B1(n_114),
.B2(n_123),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_158),
.B1(n_172),
.B2(n_168),
.Y(n_203)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_111),
.B(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_179),
.B(n_181),
.Y(n_200)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_133),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_107),
.B1(n_126),
.B2(n_84),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_103),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_187),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_107),
.B(n_82),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_177),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_107),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_185),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_154),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_178),
.C(n_159),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_194),
.C(n_209),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_216),
.B(n_193),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_217),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_180),
.B(n_211),
.C(n_201),
.Y(n_221)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_161),
.A3(n_153),
.B1(n_151),
.B2(n_148),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_211),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_210),
.B(n_216),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_161),
.B(n_164),
.C(n_184),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_207),
.B(n_192),
.C(n_210),
.D(n_195),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_SL g209 ( 
.A(n_160),
.B(n_162),
.C(n_174),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_147),
.A2(n_152),
.B(n_171),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_172),
.A3(n_147),
.B1(n_176),
.B2(n_165),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_215),
.B(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_214),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_173),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_222),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_228),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_194),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_237),
.C(n_209),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_205),
.C(n_197),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_230),
.B(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_192),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_SL g235 ( 
.A(n_190),
.B(n_215),
.C(n_204),
.Y(n_235)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_200),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_216),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_200),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_220),
.C(n_237),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_245),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_201),
.C(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_228),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_203),
.B1(n_206),
.B2(n_198),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_253),
.B1(n_226),
.B2(n_231),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_222),
.A2(n_203),
.B1(n_206),
.B2(n_212),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_252),
.B1(n_247),
.B2(n_241),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_259),
.B1(n_262),
.B2(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_255),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_232),
.B(n_230),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_254),
.B(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_219),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_252),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_264),
.B(n_266),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_235),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_202),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_258),
.B(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_244),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_273),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_221),
.B1(n_248),
.B2(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_267),
.C(n_270),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_279),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_251),
.B1(n_253),
.B2(n_257),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_280),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_261),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_281),
.B(n_274),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_286),
.B(n_255),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_278),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_269),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_250),
.B(n_275),
.C(n_272),
.D(n_268),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_286),
.A2(n_277),
.B(n_284),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_290),
.B(n_285),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_248),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_279),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_246),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.C(n_289),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_293),
.B(n_224),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_294),
.Y(n_297)
);


endmodule