module fake_jpeg_12526_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_15),
.B1(n_34),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_38),
.B1(n_41),
.B2(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_55),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_41),
.C(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_44),
.Y(n_56)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_59),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_53),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_43),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_42),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_46),
.B1(n_37),
.B2(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_50),
.C(n_46),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_58),
.C(n_8),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_70),
.B1(n_76),
.B2(n_80),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_64),
.B1(n_60),
.B2(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_9),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_19),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_78),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_7),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_20),
.C(n_28),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_80),
.C(n_76),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_13),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_10),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_12),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_23),
.B1(n_26),
.B2(n_17),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_13),
.B1(n_14),
.B2(n_87),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_94),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_88),
.A3(n_84),
.B1(n_25),
.B2(n_30),
.C1(n_21),
.C2(n_14),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_98),
.C(n_96),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_106),
.A2(n_104),
.B(n_107),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

AOI221xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_95),
.B1(n_101),
.B2(n_97),
.C(n_88),
.Y(n_112)
);


endmodule