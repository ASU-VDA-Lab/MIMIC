module fake_netlist_5_1609_n_1168 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1168);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1168;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_316;
wire n_855;
wire n_389;
wire n_785;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_949;
wire n_854;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_1145;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_1163;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_1108;
wire n_908;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_1009;
wire n_1148;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_1149;
wire n_882;
wire n_243;
wire n_398;
wire n_1146;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_1020;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_1070;
wire n_777;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_990;
wire n_836;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_1093;
wire n_722;
wire n_907;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_1041;
wire n_989;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_846;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_1052;
wire n_963;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_607;
wire n_575;
wire n_354;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_647;
wire n_707;
wire n_710;
wire n_832;
wire n_695;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_1136;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1160;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1032;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_985;
wire n_904;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_104),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_74),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_91),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_217),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_130),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_164),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_126),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_162),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_155),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_89),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_31),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_37),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_117),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_61),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_38),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_31),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_29),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_57),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_24),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_131),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_84),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_122),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_13),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_151),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_11),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_27),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_133),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_146),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_36),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_115),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_169),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_77),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_54),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_109),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_113),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_190),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_127),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_88),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_189),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_163),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_213),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_144),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_85),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_129),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_14),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_166),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_119),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_110),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_5),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_68),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_192),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_64),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_81),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_181),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_23),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_142),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_52),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_179),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_145),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_46),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_34),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_254),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_235),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_230),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_227),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_242),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_251),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_279),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_243),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_252),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_285),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_243),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_223),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_222),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_225),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_232),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_262),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_224),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_271),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_252),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_252),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_252),
.Y(n_343)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_303),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_236),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_260),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_309),
.A2(n_228),
.B(n_226),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_307),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_303),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_317),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_317),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

OA21x2_ASAP7_75t_L g357 ( 
.A1(n_309),
.A2(n_231),
.B(n_229),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_325),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_234),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_295),
.A2(n_267),
.B1(n_249),
.B2(n_257),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_238),
.B(n_237),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_301),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

OAI22x1_ASAP7_75t_R g367 ( 
.A1(n_333),
.A2(n_273),
.B1(n_291),
.B2(n_289),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_318),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_298),
.B(n_239),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_333),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_295),
.A2(n_292),
.B1(n_287),
.B2(n_286),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_33),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_300),
.A2(n_282),
.B1(n_281),
.B2(n_280),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_294),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_343),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_320),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_296),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_302),
.B(n_240),
.Y(n_383)
);

CKINVDCx11_ASAP7_75t_R g384 ( 
.A(n_334),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_330),
.B(n_278),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_304),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_305),
.A2(n_246),
.B(n_241),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_314),
.A2(n_274),
.B1(n_270),
.B2(n_269),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_268),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_334),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_307),
.B(n_250),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_R g402 ( 
.A(n_396),
.B(n_338),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_324),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_384),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_374),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_397),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_397),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g409 ( 
.A(n_349),
.B(n_314),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_349),
.B(n_323),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_L g411 ( 
.A1(n_392),
.A2(n_331),
.B1(n_339),
.B2(n_340),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_397),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_361),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_398),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_R g416 ( 
.A(n_395),
.B(n_323),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_370),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_372),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_R g424 ( 
.A(n_359),
.B(n_324),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_345),
.B(n_346),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_398),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_387),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_387),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_367),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_387),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_377),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_375),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_385),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_392),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_362),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_382),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_362),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_367),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_345),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_352),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_398),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_394),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_394),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_352),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_365),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_365),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_394),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_383),
.B(n_312),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_386),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_394),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_365),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_383),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_383),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_383),
.B(n_315),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_393),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_393),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_393),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_388),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_388),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_L g467 ( 
.A1(n_381),
.A2(n_331),
.B1(n_306),
.B2(n_336),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_390),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_R g469 ( 
.A(n_391),
.B(n_335),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_347),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_371),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_391),
.B(n_336),
.Y(n_472)
);

AO21x2_ASAP7_75t_L g473 ( 
.A1(n_364),
.A2(n_312),
.B(n_256),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_417),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_425),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_420),
.B(n_380),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_419),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_422),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_406),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

CKINVDCx8_ASAP7_75t_R g483 ( 
.A(n_404),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_335),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_443),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_399),
.B(n_347),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_444),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_381),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_465),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_380),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_427),
.B(n_255),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_428),
.B(n_258),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_454),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_472),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_380),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_437),
.A2(n_347),
.B1(n_357),
.B2(n_391),
.Y(n_501)
);

NAND3x1_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_391),
.C(n_368),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_380),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_414),
.B(n_386),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_470),
.A2(n_435),
.B1(n_434),
.B2(n_411),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_432),
.B(n_264),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_460),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_463),
.B(n_347),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_461),
.B(n_357),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_467),
.B(n_357),
.Y(n_514)
);

AND2x6_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_386),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_455),
.B(n_380),
.Y(n_516)
);

AO22x2_ASAP7_75t_L g517 ( 
.A1(n_431),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_410),
.B(n_357),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_410),
.B(n_369),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_433),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_469),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_403),
.B(n_265),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_421),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_455),
.B(n_380),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_426),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_449),
.B(n_369),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_423),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_458),
.B(n_389),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_459),
.B(n_389),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_455),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_423),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_429),
.B(n_386),
.Y(n_533)
);

NOR3xp33_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_364),
.C(n_360),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_438),
.A2(n_360),
.B1(n_368),
.B2(n_356),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_457),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_429),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_447),
.B(n_390),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_407),
.B(n_356),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_448),
.B(n_390),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_413),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_456),
.B(n_390),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_408),
.B(n_412),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_442),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_452),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_452),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_416),
.B(n_363),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_426),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_473),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_473),
.B(n_386),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_431),
.B(n_390),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_416),
.B(n_373),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_469),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_424),
.Y(n_558)
);

INVxp33_ASAP7_75t_SL g559 ( 
.A(n_481),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_486),
.A2(n_440),
.B1(n_441),
.B2(n_418),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_505),
.B(n_424),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_478),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_L g566 ( 
.A(n_551),
.B(n_35),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_487),
.B(n_373),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_483),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_484),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_504),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_499),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_527),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_505),
.B(n_402),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_527),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_505),
.B(n_402),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_526),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_508),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_486),
.B(n_363),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_496),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_497),
.B(n_355),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_489),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_488),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_490),
.B(n_366),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_501),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_489),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_482),
.B(n_355),
.Y(n_588)
);

AOI211xp5_ASAP7_75t_L g589 ( 
.A1(n_535),
.A2(n_366),
.B(n_355),
.C(n_351),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_480),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_526),
.B(n_355),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_480),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_476),
.B(n_376),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_538),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_543),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_541),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_514),
.A2(n_376),
.B1(n_366),
.B2(n_358),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_513),
.A2(n_376),
.B1(n_351),
.B2(n_350),
.Y(n_598)
);

BUFx8_ASAP7_75t_L g599 ( 
.A(n_553),
.Y(n_599)
);

BUFx8_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_539),
.Y(n_601)
);

NAND2x1p5_ASAP7_75t_L g602 ( 
.A(n_526),
.B(n_348),
.Y(n_602)
);

AO22x2_ASAP7_75t_L g603 ( 
.A1(n_501),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_512),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_476),
.B(n_376),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_482),
.B(n_376),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_551),
.B(n_376),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_482),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_545),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_547),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_520),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_498),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_553),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_524),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_528),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_532),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_548),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_546),
.B(n_3),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_536),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_549),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_521),
.B(n_376),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_494),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_533),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_498),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_511),
.B(n_4),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_558),
.B(n_509),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_498),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_567),
.A2(n_500),
.B(n_554),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_613),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_567),
.A2(n_554),
.B(n_556),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_593),
.A2(n_556),
.B(n_503),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_619),
.B(n_509),
.C(n_627),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_562),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_578),
.A2(n_535),
.B(n_555),
.C(n_557),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_596),
.B(n_519),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_604),
.B(n_550),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_593),
.A2(n_531),
.B(n_479),
.Y(n_638)
);

BUFx12f_ASAP7_75t_L g639 ( 
.A(n_599),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_584),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_604),
.A2(n_518),
.B1(n_542),
.B2(n_552),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_606),
.A2(n_531),
.B(n_479),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_606),
.A2(n_525),
.B(n_516),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_623),
.B(n_563),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_607),
.A2(n_525),
.B(n_516),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_564),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_613),
.B(n_495),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_607),
.A2(n_544),
.B(n_540),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_620),
.B(n_537),
.C(n_522),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_570),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_559),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_572),
.B(n_495),
.Y(n_652)
);

O2A1O1Ixp5_ASAP7_75t_L g653 ( 
.A1(n_590),
.A2(n_530),
.B(n_529),
.C(n_552),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_565),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_599),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_580),
.B(n_575),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_597),
.A2(n_491),
.B(n_523),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_569),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_577),
.B(n_492),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_624),
.A2(n_510),
.B(n_493),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_582),
.A2(n_608),
.B(n_566),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_577),
.B(n_534),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_581),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_582),
.A2(n_507),
.B(n_354),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_592),
.A2(n_502),
.B1(n_517),
.B2(n_507),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_608),
.A2(n_507),
.B(n_354),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_626),
.B(n_517),
.C(n_358),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_568),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_566),
.A2(n_507),
.B(n_354),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_614),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_561),
.A2(n_348),
.B(n_350),
.C(n_8),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_585),
.B(n_515),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_595),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_583),
.B(n_515),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_588),
.A2(n_609),
.B(n_625),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_588),
.A2(n_354),
.B(n_344),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_598),
.A2(n_354),
.B(n_344),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_571),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_598),
.A2(n_354),
.B1(n_358),
.B2(n_515),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_587),
.B(n_515),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_622),
.A2(n_344),
.B(n_358),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_579),
.Y(n_683)
);

AO21x1_ASAP7_75t_L g684 ( 
.A1(n_589),
.A2(n_6),
.B(n_7),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_605),
.A2(n_40),
.B(n_39),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_589),
.B(n_358),
.C(n_6),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_573),
.A2(n_358),
.B1(n_8),
.B2(n_9),
.Y(n_687)
);

AOI21x1_ASAP7_75t_L g688 ( 
.A1(n_594),
.A2(n_344),
.B(n_43),
.Y(n_688)
);

OAI21xp33_ASAP7_75t_L g689 ( 
.A1(n_576),
.A2(n_7),
.B(n_9),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_613),
.A2(n_344),
.B1(n_114),
.B2(n_116),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_622),
.A2(n_344),
.B1(n_112),
.B2(n_118),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_601),
.A2(n_610),
.B(n_611),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_612),
.B(n_42),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_616),
.A2(n_45),
.B(n_44),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_600),
.Y(n_695)
);

OAI221xp5_ASAP7_75t_L g696 ( 
.A1(n_633),
.A2(n_617),
.B1(n_621),
.B2(n_618),
.C(n_615),
.Y(n_696)
);

AND2x2_ASAP7_75t_SL g697 ( 
.A(n_655),
.B(n_625),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_634),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_SL g699 ( 
.A(n_651),
.B(n_628),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_637),
.B(n_609),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_636),
.B(n_628),
.Y(n_701)
);

CKINVDCx14_ASAP7_75t_R g702 ( 
.A(n_640),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_635),
.A2(n_591),
.B(n_602),
.C(n_586),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_673),
.A2(n_628),
.B1(n_603),
.B2(n_586),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_631),
.A2(n_603),
.B(n_560),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_656),
.B(n_649),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_669),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_679),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_644),
.B(n_600),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_631),
.A2(n_560),
.B(n_48),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_683),
.B(n_47),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_652),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_687),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_660),
.B(n_10),
.C(n_12),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_629),
.A2(n_51),
.B(n_49),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_646),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_654),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_630),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_663),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_659),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_674),
.B(n_15),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_639),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_650),
.B(n_16),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_671),
.B(n_647),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_695),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_629),
.A2(n_55),
.B(n_53),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_662),
.A2(n_132),
.B(n_220),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_630),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_661),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_689),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_657),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_668),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_686),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_675),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_692),
.B(n_23),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_658),
.A2(n_138),
.B(n_219),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_632),
.B(n_24),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_681),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_684),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_672),
.B(n_25),
.C(n_26),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_666),
.B(n_25),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_632),
.B(n_26),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_685),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_653),
.Y(n_745)
);

NAND3xp33_ASAP7_75t_SL g746 ( 
.A(n_691),
.B(n_27),
.C(n_28),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_690),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_693),
.B(n_28),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_676),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_694),
.Y(n_750)
);

AO32x1_ASAP7_75t_L g751 ( 
.A1(n_641),
.A2(n_29),
.A3(n_30),
.B1(n_32),
.B2(n_56),
.Y(n_751)
);

AND2x6_ASAP7_75t_L g752 ( 
.A(n_648),
.B(n_58),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_645),
.B(n_30),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_694),
.B(n_32),
.Y(n_754)
);

OR2x6_ASAP7_75t_SL g755 ( 
.A(n_680),
.B(n_59),
.Y(n_755)
);

OAI21x1_ASAP7_75t_L g756 ( 
.A1(n_638),
.A2(n_60),
.B(n_62),
.Y(n_756)
);

BUFx8_ASAP7_75t_SL g757 ( 
.A(n_688),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_682),
.Y(n_758)
);

BUFx4_ASAP7_75t_SL g759 ( 
.A(n_707),
.Y(n_759)
);

INVx6_ASAP7_75t_L g760 ( 
.A(n_726),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_725),
.B(n_682),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_729),
.Y(n_762)
);

INVx5_ASAP7_75t_L g763 ( 
.A(n_729),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_725),
.B(n_667),
.Y(n_764)
);

CKINVDCx16_ASAP7_75t_R g765 ( 
.A(n_726),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_708),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_712),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_746),
.A2(n_643),
.B1(n_642),
.B2(n_665),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_732),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_698),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_740),
.B(n_678),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_729),
.B(n_670),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_697),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_705),
.B(n_678),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_702),
.Y(n_775)
);

INVx3_ASAP7_75t_SL g776 ( 
.A(n_722),
.Y(n_776)
);

BUFx8_ASAP7_75t_L g777 ( 
.A(n_723),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_739),
.B(n_677),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_753),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_745),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_716),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_747),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_717),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_720),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_722),
.Y(n_785)
);

INVx5_ASAP7_75t_L g786 ( 
.A(n_752),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_699),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_755),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_718),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_718),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_750),
.B(n_221),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_709),
.Y(n_792)
);

CKINVDCx8_ASAP7_75t_R g793 ( 
.A(n_749),
.Y(n_793)
);

BUFx6f_ASAP7_75t_SL g794 ( 
.A(n_711),
.Y(n_794)
);

NAND2x1p5_ASAP7_75t_L g795 ( 
.A(n_735),
.B(n_71),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_700),
.B(n_218),
.Y(n_796)
);

BUFx12f_ASAP7_75t_L g797 ( 
.A(n_711),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_724),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_701),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_742),
.B(n_72),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_706),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_752),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_752),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_738),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_743),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_752),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_704),
.B(n_215),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_696),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_754),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_758),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_721),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_744),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_736),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_719),
.B(n_748),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_758),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_756),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_710),
.B(n_73),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_714),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_757),
.Y(n_819)
);

BUFx12f_ASAP7_75t_L g820 ( 
.A(n_730),
.Y(n_820)
);

BUFx2_ASAP7_75t_SL g821 ( 
.A(n_728),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_703),
.B(n_733),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_734),
.Y(n_823)
);

CKINVDCx6p67_ASAP7_75t_R g824 ( 
.A(n_741),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_731),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_715),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_713),
.Y(n_827)
);

INVx5_ASAP7_75t_SL g828 ( 
.A(n_727),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_737),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_751),
.B(n_83),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_793),
.A2(n_751),
.B1(n_87),
.B2(n_90),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_804),
.A2(n_751),
.B(n_93),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_767),
.Y(n_833)
);

CKINVDCx16_ASAP7_75t_R g834 ( 
.A(n_765),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_784),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_816),
.A2(n_86),
.B(n_94),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_823),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_784),
.Y(n_838)
);

AOI221xp5_ASAP7_75t_L g839 ( 
.A1(n_827),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.C(n_101),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_780),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_783),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_827),
.B(n_102),
.C(n_103),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_774),
.A2(n_105),
.B(n_106),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_780),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_799),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_774),
.A2(n_107),
.B(n_108),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_770),
.Y(n_847)
);

AOI21xp33_ASAP7_75t_L g848 ( 
.A1(n_804),
.A2(n_827),
.B(n_822),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_805),
.B(n_111),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_769),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_815),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_809),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_824),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_813),
.B(n_124),
.Y(n_854)
);

AOI21xp33_ASAP7_75t_L g855 ( 
.A1(n_822),
.A2(n_125),
.B(n_128),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_781),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_798),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_771),
.A2(n_134),
.B(n_135),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_810),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_802),
.B(n_136),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_810),
.A2(n_139),
.B(n_140),
.Y(n_861)
);

AO31x2_ASAP7_75t_L g862 ( 
.A1(n_771),
.A2(n_141),
.A3(n_143),
.B(n_147),
.Y(n_862)
);

OA21x2_ASAP7_75t_L g863 ( 
.A1(n_768),
.A2(n_148),
.B(n_149),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_766),
.Y(n_864)
);

OAI21x1_ASAP7_75t_L g865 ( 
.A1(n_768),
.A2(n_150),
.B(n_152),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_812),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_809),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_812),
.Y(n_868)
);

AO21x2_ASAP7_75t_L g869 ( 
.A1(n_807),
.A2(n_153),
.B(n_154),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_809),
.B(n_214),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_801),
.B(n_156),
.Y(n_871)
);

BUFx10_ASAP7_75t_L g872 ( 
.A(n_760),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_761),
.Y(n_873)
);

AO21x2_ASAP7_75t_L g874 ( 
.A1(n_807),
.A2(n_157),
.B(n_158),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_818),
.A2(n_159),
.B(n_160),
.C(n_161),
.Y(n_875)
);

OAI221xp5_ASAP7_75t_L g876 ( 
.A1(n_782),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.C(n_170),
.Y(n_876)
);

OA21x2_ASAP7_75t_L g877 ( 
.A1(n_829),
.A2(n_830),
.B(n_778),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_786),
.A2(n_171),
.B(n_172),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_818),
.A2(n_173),
.B(n_174),
.C(n_176),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_817),
.A2(n_177),
.B(n_180),
.Y(n_880)
);

AO31x2_ASAP7_75t_L g881 ( 
.A1(n_808),
.A2(n_182),
.A3(n_183),
.B(n_185),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_820),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_786),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_817),
.A2(n_191),
.B(n_193),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_761),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_773),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_764),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_825),
.A2(n_197),
.B(n_198),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_773),
.Y(n_889)
);

INVx6_ASAP7_75t_L g890 ( 
.A(n_797),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_764),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_760),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_786),
.B(n_803),
.Y(n_893)
);

BUFx2_ASAP7_75t_R g894 ( 
.A(n_892),
.Y(n_894)
);

OAI22xp33_ASAP7_75t_L g895 ( 
.A1(n_876),
.A2(n_801),
.B1(n_788),
.B2(n_819),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_835),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_838),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_875),
.A2(n_788),
.B(n_782),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_841),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_833),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_840),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_840),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_848),
.B(n_779),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_844),
.Y(n_904)
);

AO21x1_ASAP7_75t_SL g905 ( 
.A1(n_832),
.A2(n_826),
.B(n_791),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_851),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_844),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_888),
.A2(n_791),
.B(n_796),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_889),
.Y(n_909)
);

AOI21xp33_ASAP7_75t_SL g910 ( 
.A1(n_834),
.A2(n_776),
.B(n_792),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_856),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_872),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_875),
.A2(n_801),
.B1(n_787),
.B2(n_794),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_845),
.Y(n_914)
);

CKINVDCx6p67_ASAP7_75t_R g915 ( 
.A(n_892),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_847),
.B(n_779),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_856),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_877),
.B(n_814),
.Y(n_918)
);

AO21x2_ASAP7_75t_L g919 ( 
.A1(n_865),
.A2(n_796),
.B(n_800),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_877),
.B(n_828),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_857),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_857),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_864),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_831),
.A2(n_800),
.B(n_795),
.Y(n_924)
);

AOI21x1_ASAP7_75t_L g925 ( 
.A1(n_863),
.A2(n_772),
.B(n_811),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_866),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_866),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_877),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_868),
.Y(n_929)
);

BUFx10_ASAP7_75t_L g930 ( 
.A(n_890),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_868),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_867),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_872),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_885),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_879),
.A2(n_826),
.B(n_795),
.Y(n_935)
);

INVx3_ASAP7_75t_SL g936 ( 
.A(n_872),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_885),
.Y(n_937)
);

BUFx12f_ASAP7_75t_L g938 ( 
.A(n_890),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_852),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_879),
.A2(n_794),
.B1(n_806),
.B2(n_775),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_873),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_923),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_898),
.A2(n_839),
.B(n_842),
.C(n_865),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_899),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_923),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_935),
.A2(n_905),
.B1(n_924),
.B2(n_895),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_911),
.Y(n_947)
);

NOR3xp33_ASAP7_75t_SL g948 ( 
.A(n_940),
.B(n_871),
.C(n_886),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_909),
.B(n_891),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_911),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_934),
.B(n_891),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_903),
.Y(n_952)
);

AOI211xp5_ASAP7_75t_L g953 ( 
.A1(n_913),
.A2(n_855),
.B(n_853),
.C(n_870),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_SL g954 ( 
.A(n_924),
.B(n_903),
.C(n_910),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_915),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_R g956 ( 
.A(n_915),
.B(n_883),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_902),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_905),
.A2(n_887),
.B1(n_873),
.B2(n_874),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_901),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_R g960 ( 
.A(n_916),
.B(n_852),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_900),
.B(n_850),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_R g962 ( 
.A(n_938),
.B(n_883),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_R g963 ( 
.A(n_918),
.B(n_863),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_914),
.B(n_887),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_921),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_938),
.B(n_883),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_932),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_937),
.B(n_859),
.Y(n_968)
);

NAND2xp33_ASAP7_75t_SL g969 ( 
.A(n_936),
.B(n_860),
.Y(n_969)
);

CKINVDCx16_ASAP7_75t_R g970 ( 
.A(n_912),
.Y(n_970)
);

CKINVDCx16_ASAP7_75t_R g971 ( 
.A(n_912),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_918),
.B(n_863),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_906),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_896),
.B(n_859),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_939),
.B(n_870),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_939),
.B(n_859),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_894),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_921),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_936),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_SL g980 ( 
.A(n_920),
.B(n_882),
.C(n_837),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_942),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_967),
.B(n_959),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_942),
.Y(n_983)
);

BUFx2_ASAP7_75t_SL g984 ( 
.A(n_973),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_979),
.B(n_933),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_972),
.B(n_928),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_957),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_955),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_945),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_952),
.B(n_920),
.Y(n_990)
);

OAI221xp5_ASAP7_75t_L g991 ( 
.A1(n_946),
.A2(n_890),
.B1(n_893),
.B2(n_933),
.C(n_931),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_L g992 ( 
.A1(n_954),
.A2(n_927),
.B1(n_929),
.B2(n_926),
.C(n_897),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_945),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_976),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_947),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_949),
.B(n_917),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_947),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_950),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_952),
.B(n_973),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_950),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_965),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_952),
.B(n_928),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_973),
.B(n_941),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_943),
.A2(n_878),
.B(n_919),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_987),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_988),
.B(n_961),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_995),
.Y(n_1007)
);

AOI221xp5_ASAP7_75t_L g1008 ( 
.A1(n_992),
.A2(n_943),
.B1(n_944),
.B2(n_974),
.C(n_964),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_1004),
.A2(n_925),
.B(n_958),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_998),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_983),
.Y(n_1011)
);

CKINVDCx14_ASAP7_75t_R g1012 ( 
.A(n_988),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_995),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_991),
.A2(n_953),
.B1(n_948),
.B2(n_970),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_988),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_983),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_985),
.A2(n_969),
.B(n_980),
.C(n_977),
.Y(n_1017)
);

OA21x2_ASAP7_75t_L g1018 ( 
.A1(n_1002),
.A2(n_1000),
.B(n_993),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_996),
.A2(n_969),
.B(n_874),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_997),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_993),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1001),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_990),
.B(n_956),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1006),
.B(n_999),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1005),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_1011),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1023),
.B(n_999),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1016),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_1015),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1018),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1021),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1023),
.B(n_990),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1008),
.B(n_982),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1007),
.B(n_1002),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1012),
.B(n_1010),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1022),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1012),
.B(n_994),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1035),
.B(n_971),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1035),
.B(n_1017),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1037),
.B(n_1017),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_1029),
.B(n_1032),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_1029),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1027),
.B(n_994),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1030),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1027),
.B(n_1014),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_1039),
.B(n_1040),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1041),
.B(n_1025),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1038),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_1041),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_1045),
.B(n_1033),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1042),
.B(n_1036),
.Y(n_1051)
);

AND3x2_ASAP7_75t_L g1052 ( 
.A(n_1044),
.B(n_1024),
.C(n_1043),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1049),
.B(n_1041),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_1046),
.B(n_1050),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_1048),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_1047),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1051),
.B(n_1024),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1052),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1050),
.B(n_1029),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1048),
.B(n_1029),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_1046),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1051),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1051),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1061),
.B(n_1034),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1056),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1056),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1055),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1061),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_1053),
.B(n_1044),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_1058),
.B(n_1028),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_1062),
.B(n_1063),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_1069),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1068),
.B(n_1054),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1065),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1066),
.A2(n_1054),
.B(n_1059),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1068),
.B(n_1057),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1070),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_1067),
.A2(n_1060),
.B(n_1019),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1073),
.B(n_1064),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_1072),
.B(n_1071),
.Y(n_1080)
);

NAND2xp33_ASAP7_75t_SL g1081 ( 
.A(n_1076),
.B(n_1077),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1074),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1075),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1083),
.B(n_1078),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1081),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_1079),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1080),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_SL g1088 ( 
.A(n_1082),
.B(n_785),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1079),
.Y(n_1089)
);

OAI21xp33_ASAP7_75t_SL g1090 ( 
.A1(n_1085),
.A2(n_1030),
.B(n_1026),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_SL g1091 ( 
.A1(n_1086),
.A2(n_1031),
.B1(n_984),
.B2(n_1007),
.C(n_1020),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1087),
.B(n_1026),
.Y(n_1092)
);

NAND4xp25_ASAP7_75t_L g1093 ( 
.A(n_1089),
.B(n_759),
.C(n_960),
.D(n_860),
.Y(n_1093)
);

HAxp5_ASAP7_75t_SL g1094 ( 
.A(n_1088),
.B(n_759),
.CON(n_1094),
.SN(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1084),
.B(n_1034),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1092),
.A2(n_1084),
.B1(n_1034),
.B2(n_890),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_1090),
.A2(n_777),
.B(n_849),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_R g1098 ( 
.A(n_1095),
.B(n_777),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1094),
.Y(n_1099)
);

NAND4xp25_ASAP7_75t_SL g1100 ( 
.A(n_1091),
.B(n_854),
.C(n_1020),
.D(n_1013),
.Y(n_1100)
);

OAI211xp5_ASAP7_75t_L g1101 ( 
.A1(n_1097),
.A2(n_1093),
.B(n_956),
.C(n_962),
.Y(n_1101)
);

AOI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1096),
.A2(n_860),
.B1(n_984),
.B2(n_854),
.C(n_874),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1099),
.Y(n_1103)
);

AOI222xp33_ASAP7_75t_L g1104 ( 
.A1(n_1100),
.A2(n_1009),
.B1(n_1013),
.B2(n_930),
.C1(n_828),
.C2(n_843),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1098),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1097),
.A2(n_869),
.B(n_1018),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1097),
.A2(n_880),
.B(n_884),
.C(n_843),
.Y(n_1107)
);

AOI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1097),
.A2(n_869),
.B1(n_762),
.B2(n_789),
.C(n_858),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1103),
.B(n_763),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_L g1110 ( 
.A(n_1105),
.B(n_763),
.C(n_762),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1101),
.Y(n_1111)
);

O2A1O1Ixp5_ASAP7_75t_L g1112 ( 
.A1(n_1106),
.A2(n_981),
.B(n_997),
.C(n_1000),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1107),
.A2(n_869),
.B(n_858),
.C(n_1018),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1108),
.A2(n_763),
.B1(n_963),
.B2(n_989),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_1104),
.A2(n_199),
.B(n_200),
.C(n_202),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1102),
.A2(n_762),
.B1(n_858),
.B2(n_989),
.C(n_981),
.Y(n_1116)
);

AOI321xp33_ASAP7_75t_L g1117 ( 
.A1(n_1103),
.A2(n_975),
.A3(n_968),
.B1(n_772),
.B2(n_951),
.C(n_1003),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_1103),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1118),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1111),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1110),
.Y(n_1121)
);

XNOR2xp5_ASAP7_75t_L g1122 ( 
.A(n_1109),
.B(n_203),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_L g1123 ( 
.A(n_1115),
.B(n_880),
.C(n_884),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_1112),
.B(n_861),
.C(n_846),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1116),
.B(n_881),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1114),
.Y(n_1126)
);

NAND4xp25_ASAP7_75t_SL g1127 ( 
.A(n_1113),
.B(n_986),
.C(n_1003),
.D(n_930),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_L g1128 ( 
.A(n_1117),
.B(n_861),
.C(n_846),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1109),
.A2(n_836),
.B(n_893),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1118),
.B(n_881),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_1118),
.B(n_986),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_1119),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_1120),
.Y(n_1133)
);

OAI21xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1127),
.A2(n_836),
.B(n_930),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1122),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1131),
.B(n_204),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1121),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1126),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_1130),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1132),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1138),
.A2(n_1123),
.B(n_1125),
.Y(n_1141)
);

AO22x2_ASAP7_75t_L g1142 ( 
.A1(n_1137),
.A2(n_1129),
.B1(n_1124),
.B2(n_1128),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1133),
.A2(n_968),
.B1(n_790),
.B2(n_919),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_1135),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_1139),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1136),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1145),
.B(n_1134),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1140),
.B(n_205),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1144),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1149),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1150),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1151),
.A2(n_1141),
.B(n_1147),
.Y(n_1152)
);

OA22x2_ASAP7_75t_L g1153 ( 
.A1(n_1152),
.A2(n_1146),
.B1(n_1142),
.B2(n_1143),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1152),
.A2(n_1148),
.B(n_1142),
.C(n_209),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1152),
.B(n_207),
.Y(n_1155)
);

AOI222xp33_ASAP7_75t_L g1156 ( 
.A1(n_1155),
.A2(n_790),
.B1(n_968),
.B2(n_211),
.C1(n_212),
.C2(n_208),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1153),
.A2(n_908),
.B1(n_790),
.B2(n_828),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1154),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1155),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_R g1160 ( 
.A1(n_1158),
.A2(n_1159),
.B1(n_1156),
.B2(n_1157),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_SL g1161 ( 
.A1(n_1158),
.A2(n_210),
.B1(n_962),
.B2(n_966),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1158),
.A2(n_966),
.B1(n_821),
.B2(n_919),
.Y(n_1162)
);

AOI222xp33_ASAP7_75t_L g1163 ( 
.A1(n_1158),
.A2(n_922),
.B1(n_965),
.B2(n_978),
.C1(n_904),
.C2(n_907),
.Y(n_1163)
);

OR2x6_ASAP7_75t_L g1164 ( 
.A(n_1160),
.B(n_908),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1161),
.A2(n_925),
.B(n_881),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1163),
.B(n_862),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1164),
.A2(n_1162),
.B(n_881),
.Y(n_1167)
);

AOI211xp5_ASAP7_75t_L g1168 ( 
.A1(n_1167),
.A2(n_1166),
.B(n_1165),
.C(n_881),
.Y(n_1168)
);


endmodule