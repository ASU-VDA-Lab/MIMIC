module fake_ariane_3173_n_1752 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1752);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1752;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_76),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_41),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_104),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_100),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_45),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_28),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_12),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_74),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_51),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_13),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_43),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_75),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_41),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_48),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_83),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_67),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_40),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_45),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_22),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_37),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_48),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_107),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_87),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_47),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_117),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_25),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_60),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_81),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_132),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_122),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_153),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_26),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_63),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_29),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_9),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_18),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_20),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_131),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_46),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_155),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_16),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_37),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_52),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_101),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_119),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_136),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_30),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_65),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_86),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_89),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_62),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_4),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_103),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_109),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_125),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_42),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_55),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_133),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_143),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_93),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_108),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_121),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_23),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_47),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_22),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_32),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_14),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_113),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_88),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_10),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_5),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_72),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_9),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_66),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_82),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_105),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_73),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_49),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_54),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_80),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_20),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_140),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_126),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_29),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_21),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_137),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_12),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_141),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_129),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_77),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_59),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_25),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_106),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_91),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_61),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_71),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_154),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_40),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_60),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_34),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_151),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_32),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_139),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_27),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_49),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_46),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_0),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_59),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_54),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_92),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_79),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_2),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_78),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_27),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_55),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_128),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_36),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_7),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_111),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_150),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_112),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_50),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_43),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_17),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_0),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_162),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_222),
.B(n_1),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_252),
.B(n_2),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_165),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_198),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_179),
.B(n_3),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_185),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_191),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_299),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_229),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_181),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_178),
.B(n_182),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_181),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_181),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_194),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_240),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_201),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_179),
.B(n_6),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_181),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_238),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_181),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_210),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_210),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_166),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_281),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_203),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_210),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_210),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_210),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_211),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_211),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_211),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_189),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_309),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_211),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_204),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_296),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_276),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_303),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_205),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_276),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_208),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_276),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_212),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_215),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_183),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_183),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_186),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_307),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_220),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_206),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_238),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_221),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_159),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_206),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_249),
.B(n_6),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

CKINVDCx6p67_ASAP7_75t_R g382 ( 
.A(n_378),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_314),
.B(n_224),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_166),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_316),
.B(n_227),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_249),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_260),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_325),
.B(n_228),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_260),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_326),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_327),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_234),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_340),
.B(n_163),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_235),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_340),
.B(n_163),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_331),
.A2(n_306),
.B(n_250),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_377),
.B(n_289),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_318),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_352),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_352),
.B(n_289),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_345),
.B(n_167),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_349),
.B(n_236),
.Y(n_439)
);

CKINVDCx6p67_ASAP7_75t_R g440 ( 
.A(n_311),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_349),
.B(n_265),
.Y(n_441)
);

NOR2x1_ASAP7_75t_L g442 ( 
.A(n_350),
.B(n_306),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_368),
.B(n_370),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_350),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_351),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_398),
.Y(n_446)
);

OR2x6_ASAP7_75t_L g447 ( 
.A(n_411),
.B(n_322),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_384),
.B(n_319),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_423),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_354),
.Y(n_450)
);

AND3x1_ASAP7_75t_L g451 ( 
.A(n_386),
.B(n_313),
.C(n_312),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_361),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_363),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_396),
.B(n_366),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_396),
.B(n_322),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_384),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_403),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_385),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_411),
.B(n_367),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_430),
.B(n_339),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_386),
.B(n_310),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_396),
.B(n_337),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_385),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_387),
.B(n_408),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_389),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_396),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_L g477 ( 
.A(n_387),
.B(n_156),
.Y(n_477)
);

NOR2x1p5_ASAP7_75t_L g478 ( 
.A(n_382),
.B(n_320),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_381),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_392),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_411),
.B(n_337),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_403),
.Y(n_484)
);

BUFx6f_ASAP7_75t_SL g485 ( 
.A(n_396),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_389),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_390),
.B(n_380),
.C(n_353),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_396),
.A2(n_380),
.B1(n_255),
.B2(n_300),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_390),
.B(n_376),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_408),
.B(n_295),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_397),
.A2(n_160),
.B1(n_291),
.B2(n_284),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_442),
.B(n_163),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_397),
.A2(n_184),
.B1(n_302),
.B2(n_271),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_399),
.B(n_351),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_430),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_403),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_SL g506 ( 
.A1(n_438),
.A2(n_344),
.B1(n_358),
.B2(n_329),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_438),
.B(n_305),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_399),
.B(n_406),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_438),
.B(n_156),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_436),
.B(n_157),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_384),
.B(n_171),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_399),
.B(n_353),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_395),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_395),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_406),
.B(n_355),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_403),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_406),
.B(n_202),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_436),
.B(n_157),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_401),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_407),
.B(n_355),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_389),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_442),
.B(n_401),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_401),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_397),
.A2(n_261),
.B1(n_188),
.B2(n_175),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_407),
.A2(n_359),
.B(n_357),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_389),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_440),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_393),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_393),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_440),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_404),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_404),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_393),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_409),
.B(n_232),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_393),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_393),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_409),
.B(n_359),
.C(n_357),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_393),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_412),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_383),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_393),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_409),
.B(n_368),
.Y(n_553)
);

AND3x4_ASAP7_75t_L g554 ( 
.A(n_442),
.B(n_254),
.C(n_168),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_397),
.A2(n_247),
.B1(n_195),
.B2(n_254),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_394),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_412),
.B(n_362),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_388),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_394),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_412),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_404),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_405),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_388),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_405),
.B(n_158),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_405),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_394),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_394),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_394),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_394),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_388),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_410),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_414),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_402),
.A2(n_254),
.B1(n_244),
.B2(n_159),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_388),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_394),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_412),
.B(n_370),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_402),
.B(n_371),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_405),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_383),
.B(n_364),
.C(n_362),
.Y(n_579)
);

NOR2x1p5_ASAP7_75t_L g580 ( 
.A(n_382),
.B(n_170),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_412),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_405),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_413),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_413),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_422),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_422),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_413),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_444),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_383),
.A2(n_172),
.B1(n_309),
.B2(n_308),
.Y(n_589)
);

INVx8_ASAP7_75t_L g590 ( 
.A(n_414),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_402),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_444),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_402),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_467),
.B(n_382),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_550),
.B(n_391),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_446),
.B(n_454),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_458),
.A2(n_526),
.B1(n_570),
.B2(n_558),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_527),
.B(n_391),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_520),
.B(n_391),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_551),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_450),
.B(n_382),
.Y(n_602)
);

NOR2xp67_ASAP7_75t_L g603 ( 
.A(n_449),
.B(n_410),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_561),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_453),
.B(n_335),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_471),
.B(n_360),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_541),
.B(n_400),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_561),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_456),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_507),
.A2(n_400),
.B1(n_410),
.B2(n_415),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_504),
.B(n_591),
.Y(n_612)
);

AND3x2_ASAP7_75t_L g613 ( 
.A(n_532),
.B(n_440),
.C(n_372),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_578),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_L g615 ( 
.A(n_449),
.B(n_415),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_504),
.B(n_400),
.Y(n_616)
);

AND2x6_ASAP7_75t_SL g617 ( 
.A(n_498),
.B(n_443),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_468),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_468),
.Y(n_619)
);

BUFx6f_ASAP7_75t_SL g620 ( 
.A(n_447),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_578),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_591),
.B(n_420),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_593),
.B(n_420),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_451),
.A2(n_415),
.B1(n_420),
.B2(n_214),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_527),
.B(n_419),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_487),
.Y(n_627)
);

NOR2x1_ASAP7_75t_L g628 ( 
.A(n_462),
.B(n_447),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_527),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_593),
.B(n_420),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_527),
.B(n_560),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_518),
.B(n_439),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_583),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_551),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_459),
.B(n_440),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_582),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_560),
.B(n_419),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_466),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_448),
.B(n_511),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_511),
.B(n_172),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_448),
.B(n_439),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_582),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_455),
.B(n_439),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_509),
.B(n_176),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_583),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_560),
.B(n_581),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_558),
.B(n_443),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_461),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_461),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_510),
.B(n_176),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_570),
.B(n_443),
.Y(n_651)
);

BUFx5_ASAP7_75t_L g652 ( 
.A(n_572),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_521),
.B(n_290),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_574),
.B(n_443),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_574),
.B(n_441),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_463),
.B(n_441),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_563),
.B(n_290),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_474),
.B(n_441),
.Y(n_658)
);

NOR2xp67_ASAP7_75t_L g659 ( 
.A(n_494),
.B(n_416),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_474),
.B(n_419),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_551),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_447),
.A2(n_292),
.B1(n_293),
.B2(n_297),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_551),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_458),
.B(n_576),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_458),
.B(n_419),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_584),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_451),
.A2(n_214),
.B1(n_161),
.B2(n_304),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_458),
.B(n_444),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_463),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_560),
.B(n_158),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_526),
.A2(n_159),
.B1(n_244),
.B2(n_445),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_SL g672 ( 
.A(n_485),
.B(n_292),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_553),
.A2(n_445),
.B(n_416),
.C(n_421),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_545),
.B(n_549),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_577),
.B(n_444),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_577),
.B(n_444),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_447),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_584),
.Y(n_678)
);

O2A1O1Ixp5_ASAP7_75t_L g679 ( 
.A1(n_479),
.A2(n_444),
.B(n_445),
.C(n_425),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_464),
.A2(n_425),
.B(n_421),
.C(n_435),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_464),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_497),
.B(n_444),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_581),
.B(n_161),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_469),
.B(n_416),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_447),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_495),
.B(n_421),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_466),
.B(n_425),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_581),
.B(n_164),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_465),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_587),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_466),
.B(n_426),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_587),
.Y(n_692)
);

BUFx5_ASAP7_75t_L g693 ( 
.A(n_572),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_457),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_483),
.B(n_293),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_493),
.B(n_548),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_493),
.B(n_426),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_526),
.A2(n_244),
.B1(n_435),
.B2(n_433),
.Y(n_698)
);

AND2x6_ASAP7_75t_SL g699 ( 
.A(n_554),
.B(n_371),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_465),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_493),
.B(n_548),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_548),
.B(n_426),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_470),
.B(n_472),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_470),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_457),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_519),
.A2(n_432),
.B(n_428),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_500),
.B(n_373),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_535),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_472),
.B(n_428),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_484),
.B(n_297),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_473),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_508),
.A2(n_432),
.B(n_428),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g713 ( 
.A(n_532),
.B(n_308),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_475),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_473),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_551),
.B(n_164),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_475),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_476),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_588),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_476),
.B(n_432),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_480),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_480),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_481),
.B(n_482),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_481),
.B(n_433),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_SL g725 ( 
.A(n_554),
.B(n_279),
.C(n_246),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_477),
.B(n_219),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_482),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_488),
.B(n_490),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_526),
.A2(n_554),
.B1(n_485),
.B2(n_555),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_489),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_590),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_489),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_499),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_488),
.B(n_433),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_589),
.B(n_225),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_571),
.B(n_485),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_484),
.B(n_486),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_484),
.B(n_169),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_564),
.B(n_277),
.C(n_230),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_499),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_526),
.A2(n_180),
.B1(n_177),
.B2(n_174),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_525),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_490),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_525),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_590),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_491),
.Y(n_746)
);

AOI221xp5_ASAP7_75t_L g747 ( 
.A1(n_502),
.A2(n_282),
.B1(n_263),
.B2(n_243),
.C(n_242),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_526),
.A2(n_180),
.B1(n_177),
.B2(n_174),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_491),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_492),
.B(n_514),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_529),
.B(n_373),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_573),
.B(n_239),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_492),
.B(n_435),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_531),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_514),
.B(n_169),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_506),
.B(n_375),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_515),
.B(n_173),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_515),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_517),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_505),
.B(n_546),
.Y(n_760)
);

O2A1O1Ixp5_ASAP7_75t_L g761 ( 
.A1(n_586),
.A2(n_437),
.B(n_434),
.C(n_431),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_517),
.B(n_173),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_522),
.B(n_294),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_522),
.B(n_294),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_523),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_596),
.B(n_523),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_528),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_594),
.A2(n_526),
.B1(n_580),
.B2(n_478),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_633),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_629),
.B(n_484),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_602),
.B(n_505),
.Y(n_771)
);

OAI21xp33_ASAP7_75t_L g772 ( 
.A1(n_735),
.A2(n_257),
.B(n_241),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_761),
.A2(n_536),
.B(n_528),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_607),
.B(n_656),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_611),
.A2(n_562),
.B(n_537),
.C(n_536),
.Y(n_775)
);

AO21x1_ASAP7_75t_L g776 ( 
.A1(n_625),
.A2(n_512),
.B(n_503),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_610),
.Y(n_777)
);

AO21x1_ASAP7_75t_L g778 ( 
.A1(n_625),
.A2(n_524),
.B(n_516),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_736),
.A2(n_539),
.B(n_562),
.C(n_565),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_645),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_598),
.A2(n_586),
.B(n_460),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_598),
.A2(n_586),
.B(n_460),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_666),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_629),
.B(n_484),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_656),
.B(n_537),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_641),
.B(n_539),
.Y(n_786)
);

CKINVDCx6p67_ASAP7_75t_R g787 ( 
.A(n_635),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_731),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_651),
.B(n_565),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_595),
.A2(n_460),
.B(n_452),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_678),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_669),
.B(n_478),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_651),
.B(n_531),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_669),
.B(n_580),
.Y(n_794)
);

AOI21x1_ASAP7_75t_L g795 ( 
.A1(n_637),
.A2(n_530),
.B(n_557),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_690),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_692),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_610),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_629),
.B(n_597),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_635),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_616),
.B(n_640),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_612),
.B(n_603),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_729),
.A2(n_579),
.B1(n_494),
.B2(n_501),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_615),
.B(n_533),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_694),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_622),
.B(n_533),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_614),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_696),
.A2(n_452),
.B(n_505),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_623),
.B(n_534),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_696),
.A2(n_452),
.B(n_505),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_701),
.A2(n_546),
.B(n_588),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_630),
.B(n_534),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_701),
.A2(n_546),
.B(n_592),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_632),
.B(n_540),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_627),
.B(n_486),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_637),
.A2(n_660),
.B(n_665),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_760),
.A2(n_646),
.B(n_638),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_639),
.B(n_540),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_679),
.A2(n_673),
.B(n_680),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_647),
.B(n_542),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_654),
.B(n_542),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_SL g822 ( 
.A1(n_673),
.A2(n_592),
.B(n_543),
.C(n_575),
.Y(n_822)
);

NAND2x1p5_ASAP7_75t_L g823 ( 
.A(n_731),
.B(n_543),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_731),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_614),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_646),
.A2(n_546),
.B(n_513),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_726),
.B(n_547),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_655),
.B(n_547),
.Y(n_828)
);

AND2x2_ASAP7_75t_SL g829 ( 
.A(n_671),
.B(n_163),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_605),
.A2(n_559),
.B1(n_556),
.B2(n_552),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_705),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_680),
.A2(n_668),
.B(n_643),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_631),
.A2(n_538),
.B(n_513),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_711),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_631),
.A2(n_538),
.B(n_513),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_628),
.B(n_552),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_703),
.A2(n_538),
.B(n_513),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_657),
.B(n_556),
.Y(n_839)
);

NOR2x1_ASAP7_75t_R g840 ( 
.A(n_713),
.B(n_267),
.Y(n_840)
);

AOI222xp33_ASAP7_75t_L g841 ( 
.A1(n_606),
.A2(n_268),
.B1(n_275),
.B2(n_280),
.C1(n_287),
.C2(n_288),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_731),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_723),
.A2(n_513),
.B(n_486),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_721),
.Y(n_844)
);

AO21x1_ASAP7_75t_L g845 ( 
.A1(n_716),
.A2(n_530),
.B(n_437),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_728),
.A2(n_538),
.B(n_486),
.Y(n_846)
);

AND2x2_ASAP7_75t_SL g847 ( 
.A(n_698),
.B(n_163),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_674),
.B(n_624),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_664),
.A2(n_566),
.B(n_559),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_627),
.A2(n_658),
.B1(n_601),
.B2(n_618),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_707),
.B(n_566),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_750),
.A2(n_496),
.B(n_538),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_674),
.B(n_375),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_621),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_722),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_707),
.B(n_567),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_709),
.A2(n_568),
.B(n_575),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_730),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_627),
.A2(n_567),
.B1(n_568),
.B2(n_569),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_604),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_751),
.B(n_675),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_725),
.A2(n_579),
.B1(n_501),
.B2(n_544),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_687),
.A2(n_496),
.B(n_486),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_676),
.A2(n_644),
.B(n_662),
.C(n_682),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_667),
.A2(n_569),
.B(n_544),
.C(n_437),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_708),
.B(n_379),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_691),
.A2(n_496),
.B(n_585),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_617),
.B(n_496),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_697),
.A2(n_496),
.B(n_585),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_636),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_706),
.A2(n_501),
.B(n_418),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_636),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_751),
.B(n_501),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_702),
.A2(n_585),
.B(n_590),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_731),
.Y(n_875)
);

AND2x6_ASAP7_75t_SL g876 ( 
.A(n_650),
.B(n_379),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_737),
.A2(n_670),
.B(n_684),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_737),
.A2(n_585),
.B(n_590),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_670),
.A2(n_585),
.B(n_590),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_613),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_677),
.B(n_298),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_609),
.B(n_501),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_685),
.B(n_501),
.Y(n_883)
);

BUFx8_ASAP7_75t_L g884 ( 
.A(n_620),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_732),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_619),
.B(n_626),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_642),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_642),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_733),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_600),
.B(n_572),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_756),
.B(n_418),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_648),
.A2(n_298),
.B(n_301),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_648),
.A2(n_301),
.B(n_304),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_649),
.B(n_501),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_649),
.B(n_681),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_740),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_681),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_689),
.B(n_418),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_689),
.A2(n_418),
.B(n_437),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_712),
.A2(n_427),
.B(n_437),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_600),
.B(n_572),
.Y(n_901)
);

AOI22x1_ASAP7_75t_L g902 ( 
.A1(n_700),
.A2(n_434),
.B1(n_431),
.B2(n_427),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_700),
.B(n_418),
.Y(n_903)
);

AOI21x1_ASAP7_75t_L g904 ( 
.A1(n_720),
.A2(n_434),
.B(n_431),
.Y(n_904)
);

OAI321xp33_ASAP7_75t_L g905 ( 
.A1(n_752),
.A2(n_365),
.A3(n_364),
.B1(n_427),
.B2(n_434),
.C(n_431),
.Y(n_905)
);

BUFx2_ASAP7_75t_SL g906 ( 
.A(n_620),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_704),
.A2(n_434),
.B(n_431),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_704),
.A2(n_427),
.B(n_248),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_714),
.B(n_427),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_714),
.A2(n_424),
.B1(n_422),
.B2(n_237),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_717),
.B(n_187),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_653),
.B(n_7),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_717),
.A2(n_251),
.B(n_192),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_718),
.B(n_190),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_718),
.B(n_193),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_756),
.B(n_8),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_727),
.B(n_196),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_727),
.A2(n_365),
.B(n_414),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_745),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_743),
.A2(n_256),
.B(n_199),
.Y(n_920)
);

OAI21xp33_ASAP7_75t_L g921 ( 
.A1(n_741),
.A2(n_253),
.B(n_200),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_743),
.B(n_197),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_699),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_745),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_746),
.A2(n_424),
.B(n_422),
.C(n_283),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_746),
.A2(n_262),
.B(n_209),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_695),
.B(n_11),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_749),
.A2(n_765),
.B(n_758),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_620),
.B(n_11),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_749),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_634),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_745),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_604),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_742),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_745),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_634),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_745),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_758),
.A2(n_264),
.B(n_213),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_759),
.B(n_207),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_672),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_759),
.B(n_765),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_744),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_754),
.Y(n_943)
);

OAI22xp33_ASAP7_75t_L g944 ( 
.A1(n_748),
.A2(n_259),
.B1(n_217),
.B2(n_226),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_683),
.A2(n_270),
.B(n_231),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_608),
.B(n_719),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_672),
.A2(n_272),
.B1(n_233),
.B2(n_245),
.Y(n_947)
);

INVxp67_ASAP7_75t_R g948 ( 
.A(n_608),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_600),
.B(n_424),
.Y(n_949)
);

O2A1O1Ixp5_ASAP7_75t_L g950 ( 
.A1(n_738),
.A2(n_424),
.B(n_422),
.C(n_15),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_683),
.A2(n_216),
.B(n_258),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_719),
.B(n_266),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_724),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_912),
.A2(n_719),
.B(n_661),
.C(n_663),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_912),
.A2(n_688),
.B(n_763),
.C(n_762),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_771),
.A2(n_688),
.B(n_716),
.Y(n_956)
);

BUFx8_ASAP7_75t_L g957 ( 
.A(n_800),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_769),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_801),
.B(n_739),
.Y(n_959)
);

OAI22x1_ASAP7_75t_L g960 ( 
.A1(n_916),
.A2(n_927),
.B1(n_768),
.B2(n_848),
.Y(n_960)
);

AO32x1_ASAP7_75t_L g961 ( 
.A1(n_850),
.A2(n_710),
.A3(n_738),
.B1(n_659),
.B2(n_764),
.Y(n_961)
);

BUFx12f_ASAP7_75t_L g962 ( 
.A(n_884),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_771),
.A2(n_753),
.B(n_734),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_906),
.B(n_634),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_897),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_L g966 ( 
.A(n_927),
.B(n_747),
.C(n_710),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_766),
.A2(n_600),
.B(n_661),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_884),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_780),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_798),
.Y(n_970)
);

BUFx12f_ASAP7_75t_L g971 ( 
.A(n_880),
.Y(n_971)
);

INVxp33_ASAP7_75t_L g972 ( 
.A(n_798),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_767),
.A2(n_774),
.B(n_877),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_916),
.B(n_686),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_777),
.B(n_600),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_827),
.A2(n_663),
.B(n_661),
.Y(n_976)
);

AOI22x1_ASAP7_75t_L g977 ( 
.A1(n_817),
.A2(n_663),
.B1(n_634),
.B2(n_755),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_876),
.B(n_757),
.Y(n_978)
);

BUFx10_ASAP7_75t_L g979 ( 
.A(n_881),
.Y(n_979)
);

BUFx6f_ASAP7_75t_SL g980 ( 
.A(n_792),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_848),
.B(n_787),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_931),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_861),
.B(n_652),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_940),
.A2(n_652),
.B1(n_693),
.B2(n_269),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_924),
.B(n_693),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_822),
.A2(n_693),
.B(n_652),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_883),
.B(n_422),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_883),
.B(n_693),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_923),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_853),
.Y(n_990)
);

INVx3_ASAP7_75t_SL g991 ( 
.A(n_792),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_924),
.B(n_693),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_794),
.B(n_693),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_931),
.B(n_424),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_864),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_995)
);

INVx3_ASAP7_75t_SL g996 ( 
.A(n_794),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_904),
.A2(n_424),
.B(n_422),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_953),
.B(n_652),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_891),
.B(n_652),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_841),
.B(n_422),
.C(n_424),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_785),
.A2(n_693),
.B1(n_652),
.B2(n_274),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_802),
.B(n_652),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_866),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_881),
.B(n_17),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_822),
.A2(n_424),
.B(n_422),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_832),
.A2(n_422),
.B(n_424),
.C(n_283),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_829),
.A2(n_424),
.B1(n_417),
.B2(n_414),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_897),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_775),
.A2(n_18),
.B(n_19),
.C(n_21),
.Y(n_1009)
);

AO32x1_ASAP7_75t_L g1010 ( 
.A1(n_942),
.A2(n_943),
.A3(n_859),
.B1(n_910),
.B2(n_930),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_936),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_838),
.A2(n_223),
.B(n_273),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_930),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_783),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_868),
.B(n_223),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_816),
.A2(n_417),
.B(n_414),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_843),
.A2(n_223),
.B(n_273),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_772),
.B(n_19),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_936),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_791),
.B(n_23),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_868),
.A2(n_417),
.B1(n_414),
.B2(n_283),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_921),
.A2(n_223),
.B(n_273),
.Y(n_1022)
);

OAI22x1_ASAP7_75t_L g1023 ( 
.A1(n_929),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_840),
.B(n_24),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_948),
.B(n_30),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_836),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_796),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_797),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_944),
.B(n_31),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_944),
.B(n_223),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_875),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_788),
.B(n_842),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_805),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_825),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_846),
.A2(n_273),
.B(n_283),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_SL g1036 ( 
.A1(n_829),
.A2(n_273),
.B1(n_283),
.B2(n_38),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_860),
.B(n_31),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_831),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_933),
.B(n_33),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_875),
.B(n_33),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_847),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_775),
.A2(n_39),
.B(n_44),
.C(n_50),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_852),
.A2(n_44),
.B(n_51),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_836),
.B(n_52),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_847),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_933),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_SL g1047 ( 
.A1(n_862),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_834),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_776),
.A2(n_58),
.B(n_64),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_875),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_778),
.A2(n_928),
.B(n_867),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_851),
.B(n_417),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_873),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_779),
.A2(n_417),
.B(n_414),
.C(n_85),
.Y(n_1054)
);

XOR2x2_ASAP7_75t_L g1055 ( 
.A(n_947),
.B(n_70),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_837),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_789),
.A2(n_417),
.B1(n_414),
.B2(n_97),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_844),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_855),
.B(n_417),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_942),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_875),
.B(n_417),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_854),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_858),
.B(n_417),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_885),
.B(n_417),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_863),
.A2(n_84),
.B(n_90),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_856),
.B(n_417),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_889),
.B(n_896),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_869),
.A2(n_98),
.B(n_102),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_932),
.B(n_417),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_SL g1070 ( 
.A(n_892),
.B(n_417),
.C(n_414),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_934),
.B(n_417),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_793),
.B(n_414),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_886),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_943),
.A2(n_414),
.B1(n_115),
.B2(n_127),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_818),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_824),
.B(n_114),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_804),
.B(n_130),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_857),
.A2(n_414),
.B(n_138),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_786),
.A2(n_414),
.B1(n_145),
.B2(n_147),
.Y(n_1079)
);

NAND2x1_ASAP7_75t_L g1080 ( 
.A(n_824),
.B(n_414),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_830),
.B(n_134),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_807),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_870),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_870),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_790),
.A2(n_148),
.B(n_874),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_779),
.A2(n_799),
.B(n_839),
.C(n_905),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_828),
.A2(n_941),
.B1(n_895),
.B2(n_820),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_865),
.A2(n_799),
.B(n_819),
.C(n_821),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_814),
.B(n_911),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_932),
.B(n_788),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_865),
.A2(n_950),
.B(n_871),
.C(n_862),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_932),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_872),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_795),
.A2(n_770),
.B(n_784),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_990),
.B(n_888),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_1046),
.Y(n_1096)
);

AO31x2_ASAP7_75t_L g1097 ( 
.A1(n_1051),
.A2(n_845),
.A3(n_925),
.B(n_908),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_963),
.A2(n_973),
.B(n_986),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_966),
.B(n_945),
.C(n_951),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_963),
.A2(n_781),
.B(n_782),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_997),
.A2(n_900),
.B(n_835),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_966),
.A2(n_915),
.B(n_939),
.C(n_922),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_988),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_970),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_1051),
.A2(n_925),
.A3(n_872),
.B(n_888),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_959),
.A2(n_803),
.B(n_893),
.C(n_917),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_973),
.A2(n_770),
.B(n_784),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1085),
.A2(n_833),
.B(n_773),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1003),
.B(n_981),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1085),
.A2(n_902),
.B(n_879),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_962),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_960),
.A2(n_803),
.B1(n_914),
.B2(n_812),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_956),
.A2(n_813),
.B(n_811),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_989),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_958),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_1091),
.A2(n_1006),
.A3(n_1087),
.B(n_1012),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_968),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1029),
.A2(n_952),
.B(n_815),
.C(n_809),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1086),
.A2(n_1088),
.B(n_956),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1005),
.A2(n_899),
.B(n_907),
.Y(n_1120)
);

BUFx4_ASAP7_75t_SL g1121 ( 
.A(n_964),
.Y(n_1121)
);

OAI22x1_ASAP7_75t_L g1122 ( 
.A1(n_1018),
.A2(n_887),
.B1(n_815),
.B2(n_949),
.Y(n_1122)
);

OAI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_1004),
.A2(n_806),
.B(n_849),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_955),
.A2(n_920),
.B(n_913),
.C(n_926),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_L g1125 ( 
.A1(n_1030),
.A2(n_949),
.B(n_901),
.C(n_890),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_SL g1126 ( 
.A(n_1031),
.B(n_932),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1073),
.B(n_887),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1088),
.A2(n_808),
.B(n_810),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_986),
.A2(n_878),
.B(n_826),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_988),
.B(n_890),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_955),
.A2(n_909),
.B(n_903),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_974),
.A2(n_882),
.B(n_894),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_1012),
.A2(n_946),
.A3(n_898),
.B(n_938),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1073),
.B(n_842),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_967),
.A2(n_901),
.B(n_823),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_965),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_969),
.Y(n_1137)
);

AO21x1_ASAP7_75t_L g1138 ( 
.A1(n_1041),
.A2(n_823),
.B(n_918),
.Y(n_1138)
);

AO21x1_ASAP7_75t_L g1139 ( 
.A1(n_1045),
.A2(n_919),
.B(n_935),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1014),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1005),
.A2(n_919),
.B(n_935),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1001),
.A2(n_937),
.B(n_998),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1027),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_978),
.A2(n_937),
.B(n_1089),
.C(n_995),
.Y(n_1144)
);

OA21x2_ASAP7_75t_L g1145 ( 
.A1(n_1049),
.A2(n_1035),
.B(n_1017),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_964),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1049),
.A2(n_1035),
.B(n_1017),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_957),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_995),
.A2(n_1042),
.B(n_1009),
.C(n_1024),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_SL g1150 ( 
.A1(n_954),
.A2(n_985),
.B(n_1040),
.C(n_975),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_983),
.A2(n_967),
.B(n_976),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_977),
.A2(n_976),
.B(n_1094),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_982),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1043),
.A2(n_999),
.B(n_1072),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1078),
.A2(n_1016),
.B(n_1065),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1008),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_961),
.A2(n_1002),
.B(n_1077),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1083),
.A2(n_1084),
.A3(n_1093),
.B(n_1034),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1013),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_957),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1028),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1009),
.A2(n_1042),
.B(n_1020),
.C(n_1039),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1036),
.A2(n_1047),
.B1(n_1055),
.B2(n_1075),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1000),
.A2(n_1037),
.B(n_984),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1075),
.B(n_1067),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1026),
.B(n_964),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1060),
.B(n_979),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_979),
.B(n_1048),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1033),
.B(n_1058),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1081),
.A2(n_996),
.B1(n_991),
.B2(n_1007),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1038),
.B(n_1056),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1062),
.A2(n_1010),
.A3(n_1068),
.B(n_1065),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1068),
.A2(n_1043),
.B(n_1090),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_1044),
.B(n_980),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_982),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_982),
.B(n_1019),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_994),
.A2(n_1052),
.B(n_1066),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1053),
.B(n_1025),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_961),
.A2(n_1022),
.B(n_988),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_994),
.A2(n_1054),
.B(n_1080),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1054),
.A2(n_993),
.B(n_1076),
.C(n_1015),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1070),
.A2(n_1069),
.B(n_1061),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_980),
.B(n_1019),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_961),
.A2(n_1010),
.B(n_1076),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1082),
.B(n_987),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1079),
.A2(n_1059),
.B(n_1063),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1010),
.A2(n_1031),
.B(n_1050),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1023),
.A2(n_1057),
.A3(n_1050),
.B(n_992),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1031),
.A2(n_987),
.B(n_1092),
.Y(n_1189)
);

O2A1O1Ixp5_ASAP7_75t_L g1190 ( 
.A1(n_1064),
.A2(n_1071),
.B(n_1032),
.C(n_1019),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1074),
.A2(n_1011),
.B(n_1021),
.Y(n_1191)
);

NOR4xp25_ASAP7_75t_L g1192 ( 
.A(n_1011),
.B(n_995),
.C(n_1042),
.D(n_1009),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1011),
.A2(n_912),
.B(n_927),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_971),
.A2(n_997),
.B(n_1051),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_990),
.B(n_594),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_990),
.B(n_594),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_959),
.A2(n_927),
.B(n_912),
.C(n_966),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_963),
.A2(n_771),
.B(n_737),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_963),
.A2(n_771),
.B(n_737),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_L g1200 ( 
.A1(n_997),
.A2(n_1051),
.B(n_1017),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_972),
.B(n_606),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_SL g1202 ( 
.A(n_1036),
.B(n_829),
.Y(n_1202)
);

AO21x1_ASAP7_75t_L g1203 ( 
.A1(n_1041),
.A2(n_1045),
.B(n_912),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_959),
.A2(n_927),
.B(n_912),
.C(n_966),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_997),
.A2(n_1051),
.B(n_1085),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1051),
.A2(n_778),
.A3(n_776),
.B(n_1091),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1051),
.A2(n_778),
.A3(n_776),
.B(n_1091),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_959),
.A2(n_927),
.B(n_912),
.C(n_966),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1051),
.A2(n_778),
.A3(n_776),
.B(n_1091),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_963),
.A2(n_771),
.B(n_737),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1051),
.A2(n_778),
.A3(n_776),
.B(n_1091),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_990),
.B(n_594),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_965),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_959),
.A2(n_594),
.B1(n_912),
.B2(n_801),
.Y(n_1214)
);

NAND2x1_ASAP7_75t_L g1215 ( 
.A(n_1050),
.B(n_988),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_962),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1003),
.B(n_798),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1086),
.A2(n_1091),
.B(n_1088),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_965),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1026),
.B(n_964),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_958),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_990),
.B(n_594),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_962),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_990),
.B(n_594),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_990),
.B(n_594),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_982),
.B(n_708),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_990),
.B(n_639),
.Y(n_1227)
);

AOI221xp5_ASAP7_75t_SL g1228 ( 
.A1(n_995),
.A2(n_1042),
.B1(n_1009),
.B2(n_1029),
.C(n_912),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_958),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_990),
.B(n_594),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_958),
.Y(n_1231)
);

AO32x2_ASAP7_75t_L g1232 ( 
.A1(n_1047),
.A2(n_1036),
.A3(n_1041),
.B1(n_1045),
.B2(n_1087),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_972),
.B(n_606),
.Y(n_1233)
);

OR2x2_ASAP7_75t_L g1234 ( 
.A(n_1003),
.B(n_798),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_966),
.A2(n_912),
.B(n_927),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_SL g1236 ( 
.A(n_966),
.B(n_449),
.C(n_423),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1146),
.B(n_1215),
.Y(n_1237)
);

BUFx10_ASAP7_75t_L g1238 ( 
.A(n_1114),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1217),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1202),
.A2(n_1163),
.B1(n_1214),
.B2(n_1235),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1169),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1227),
.B(n_1201),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1202),
.A2(n_1203),
.B1(n_1218),
.B2(n_1233),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1195),
.B(n_1196),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1218),
.A2(n_1164),
.B1(n_1236),
.B2(n_1119),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1146),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1115),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1119),
.A2(n_1193),
.B1(n_1212),
.B2(n_1222),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1224),
.A2(n_1230),
.B1(n_1225),
.B2(n_1112),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1137),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1117),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1165),
.B(n_1096),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1140),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1112),
.A2(n_1109),
.B1(n_1234),
.B2(n_1232),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1098),
.Y(n_1255)
);

INVx6_ASAP7_75t_L g1256 ( 
.A(n_1146),
.Y(n_1256)
);

OAI22x1_ASAP7_75t_SL g1257 ( 
.A1(n_1148),
.A2(n_1223),
.B1(n_1216),
.B2(n_1111),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1123),
.A2(n_1178),
.B1(n_1170),
.B2(n_1174),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1228),
.A2(n_1208),
.B1(n_1204),
.B2(n_1197),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1153),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1153),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_1104),
.Y(n_1262)
);

CKINVDCx14_ASAP7_75t_R g1263 ( 
.A(n_1160),
.Y(n_1263)
);

INVx8_ASAP7_75t_L g1264 ( 
.A(n_1130),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1232),
.A2(n_1095),
.B1(n_1168),
.B2(n_1167),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1123),
.A2(n_1127),
.B1(n_1232),
.B2(n_1143),
.Y(n_1266)
);

INVx6_ASAP7_75t_L g1267 ( 
.A(n_1153),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1192),
.A2(n_1104),
.B1(n_1183),
.B2(n_1226),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1161),
.A2(n_1231),
.B1(n_1229),
.B2(n_1221),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1144),
.A2(n_1149),
.B1(n_1106),
.B2(n_1162),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_R g1271 ( 
.A1(n_1228),
.A2(n_1192),
.B1(n_1099),
.B2(n_1121),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1175),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_1102),
.A2(n_1124),
.B(n_1134),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1136),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1166),
.A2(n_1220),
.B1(n_1130),
.B2(n_1103),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1198),
.A2(n_1199),
.B1(n_1210),
.B2(n_1181),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1185),
.A2(n_1138),
.B1(n_1219),
.B2(n_1213),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1175),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1118),
.A2(n_1130),
.B1(n_1186),
.B2(n_1157),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1156),
.A2(n_1159),
.B1(n_1179),
.B2(n_1139),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1175),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1176),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1194),
.Y(n_1283)
);

INVx8_ASAP7_75t_L g1284 ( 
.A(n_1220),
.Y(n_1284)
);

BUFx2_ASAP7_75t_SL g1285 ( 
.A(n_1103),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1122),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1189),
.B(n_1190),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1180),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_1187),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1126),
.B(n_1188),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1182),
.Y(n_1291)
);

INVx6_ASAP7_75t_L g1292 ( 
.A(n_1182),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1186),
.A2(n_1154),
.B1(n_1131),
.B2(n_1142),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1184),
.A2(n_1131),
.B1(n_1154),
.B2(n_1191),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1107),
.A2(n_1128),
.B1(n_1135),
.B2(n_1145),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1135),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1188),
.B(n_1211),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1188),
.B(n_1211),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1105),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1132),
.A2(n_1145),
.B1(n_1147),
.B2(n_1177),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1105),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1206),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1147),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1128),
.A2(n_1151),
.B1(n_1113),
.B2(n_1100),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1206),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1150),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1129),
.A2(n_1152),
.B1(n_1200),
.B2(n_1116),
.Y(n_1307)
);

CKINVDCx11_ASAP7_75t_R g1308 ( 
.A(n_1125),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1152),
.A2(n_1116),
.B1(n_1209),
.B2(n_1211),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1141),
.Y(n_1310)
);

AOI22x1_ASAP7_75t_L g1311 ( 
.A1(n_1206),
.A2(n_1209),
.B1(n_1207),
.B2(n_1173),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1207),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1108),
.A2(n_1116),
.B1(n_1110),
.B2(n_1155),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1205),
.A2(n_1207),
.B1(n_1209),
.B2(n_1101),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1133),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1133),
.Y(n_1316)
);

INVx4_ASAP7_75t_SL g1317 ( 
.A(n_1133),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1097),
.B(n_1172),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1097),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1097),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1172),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1120),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1172),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1202),
.A2(n_916),
.B1(n_1163),
.B2(n_1036),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1117),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1146),
.B(n_1215),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1202),
.A2(n_1214),
.B1(n_1235),
.B2(n_1045),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1202),
.A2(n_594),
.B1(n_606),
.B2(n_1214),
.Y(n_1328)
);

CKINVDCx6p67_ASAP7_75t_R g1329 ( 
.A(n_1148),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1171),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1158),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1146),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1202),
.A2(n_1214),
.B1(n_1235),
.B2(n_1045),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1214),
.A2(n_1204),
.B1(n_1208),
.B2(n_1197),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1171),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1217),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1146),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1202),
.A2(n_1036),
.B1(n_916),
.B2(n_1214),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1148),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1214),
.B(n_990),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1153),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1226),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1171),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1153),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1202),
.A2(n_594),
.B1(n_606),
.B2(n_1214),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1117),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1153),
.Y(n_1347)
);

INVx6_ASAP7_75t_L g1348 ( 
.A(n_1146),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1202),
.A2(n_594),
.B1(n_606),
.B2(n_1214),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1202),
.A2(n_916),
.B1(n_1163),
.B2(n_1036),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1202),
.A2(n_1036),
.B1(n_916),
.B2(n_1214),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1148),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1171),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1226),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1202),
.A2(n_1036),
.B1(n_916),
.B2(n_1214),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1214),
.A2(n_1204),
.B(n_1197),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1171),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1244),
.B(n_1252),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1302),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1305),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1288),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1288),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1288),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1239),
.B(n_1336),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1267),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1264),
.B(n_1289),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1318),
.B(n_1296),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1247),
.B(n_1250),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1253),
.B(n_1242),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1328),
.A2(n_1349),
.B(n_1345),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1240),
.A2(n_1324),
.B1(n_1350),
.B2(n_1338),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1288),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1331),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1356),
.B(n_1243),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1243),
.B(n_1304),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1269),
.B(n_1320),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1262),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1276),
.A2(n_1334),
.B(n_1327),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1267),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1266),
.B(n_1321),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1249),
.B(n_1241),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1278),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1283),
.B(n_1317),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1249),
.B(n_1248),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1290),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1307),
.A2(n_1311),
.B(n_1300),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1297),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1323),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1298),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1312),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1312),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1301),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1265),
.A2(n_1309),
.B(n_1254),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1300),
.A2(n_1295),
.B(n_1322),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1259),
.A2(n_1333),
.B1(n_1327),
.B2(n_1254),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1293),
.A2(n_1270),
.A3(n_1279),
.B(n_1323),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1264),
.B(n_1287),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1264),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1265),
.A2(n_1294),
.B(n_1321),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1280),
.A2(n_1255),
.B(n_1273),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1316),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1292),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1340),
.B(n_1330),
.Y(n_1403)
);

AO21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1240),
.A2(n_1280),
.B(n_1245),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1324),
.A2(n_1350),
.B(n_1355),
.C(n_1351),
.Y(n_1405)
);

BUFx4f_ASAP7_75t_SL g1406 ( 
.A(n_1325),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1248),
.B(n_1357),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1299),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1316),
.Y(n_1409)
);

AOI21xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1294),
.A2(n_1257),
.B(n_1268),
.Y(n_1410)
);

OAI222xp33_ASAP7_75t_L g1411 ( 
.A1(n_1258),
.A2(n_1266),
.B1(n_1291),
.B2(n_1275),
.C1(n_1343),
.C2(n_1335),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_SL g1412 ( 
.A1(n_1346),
.A2(n_1271),
.B(n_1282),
.C(n_1306),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1319),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1284),
.B(n_1319),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1255),
.A2(n_1310),
.B(n_1353),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1315),
.A2(n_1261),
.B(n_1260),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1319),
.B(n_1314),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1277),
.A2(n_1237),
.B(n_1326),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1317),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1267),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1272),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1303),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1274),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1286),
.B(n_1285),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1313),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1292),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1272),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1308),
.A2(n_1332),
.B(n_1348),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1341),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1341),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1344),
.B(n_1347),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1256),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1246),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1344),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1347),
.B(n_1354),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1369),
.B(n_1263),
.Y(n_1436)
);

AOI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1371),
.A2(n_1342),
.B1(n_1263),
.B2(n_1284),
.C(n_1246),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1369),
.B(n_1238),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1364),
.B(n_1329),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1373),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1405),
.A2(n_1281),
.B1(n_1251),
.B2(n_1256),
.Y(n_1441)
);

A2O1A1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1378),
.A2(n_1370),
.B(n_1374),
.C(n_1410),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1366),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1367),
.B(n_1238),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1374),
.B(n_1339),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1367),
.B(n_1352),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1410),
.A2(n_1337),
.B(n_1348),
.C(n_1375),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1395),
.A2(n_1375),
.B1(n_1384),
.B2(n_1381),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1397),
.B(n_1417),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1400),
.A2(n_1425),
.B(n_1426),
.Y(n_1450)
);

OAI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1425),
.A2(n_1412),
.B(n_1407),
.C(n_1400),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1393),
.A2(n_1399),
.B(n_1386),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1402),
.B(n_1424),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1415),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1406),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_SL g1456 ( 
.A(n_1366),
.B(n_1397),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1368),
.B(n_1403),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1358),
.B(n_1377),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1402),
.B(n_1424),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1397),
.B(n_1417),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1368),
.B(n_1403),
.Y(n_1461)
);

OAI211xp5_ASAP7_75t_L g1462 ( 
.A1(n_1400),
.A2(n_1429),
.B(n_1434),
.C(n_1430),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1400),
.A2(n_1415),
.B(n_1399),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1386),
.A2(n_1366),
.B(n_1393),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1394),
.A2(n_1411),
.B(n_1418),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1422),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1380),
.A2(n_1376),
.B1(n_1387),
.B2(n_1389),
.C(n_1385),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1382),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1383),
.B(n_1401),
.Y(n_1469)
);

AO32x2_ASAP7_75t_L g1470 ( 
.A1(n_1421),
.A2(n_1427),
.A3(n_1379),
.B1(n_1420),
.B2(n_1365),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1396),
.B(n_1431),
.Y(n_1471)
);

AO32x2_ASAP7_75t_L g1472 ( 
.A1(n_1380),
.A2(n_1385),
.A3(n_1396),
.B1(n_1389),
.B2(n_1387),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1431),
.B(n_1396),
.Y(n_1473)
);

CKINVDCx14_ASAP7_75t_R g1474 ( 
.A(n_1435),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1404),
.A2(n_1418),
.B(n_1396),
.C(n_1394),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1422),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1392),
.B(n_1359),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1423),
.Y(n_1478)
);

CKINVDCx16_ASAP7_75t_R g1479 ( 
.A(n_1398),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1404),
.A2(n_1435),
.B(n_1416),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1428),
.A2(n_1398),
.B(n_1414),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1383),
.B(n_1401),
.Y(n_1482)
);

OAI211xp5_ASAP7_75t_L g1483 ( 
.A1(n_1388),
.A2(n_1372),
.B(n_1361),
.C(n_1363),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1423),
.Y(n_1484)
);

AOI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1360),
.A2(n_1383),
.B1(n_1390),
.B2(n_1391),
.C(n_1408),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1448),
.A2(n_1428),
.B1(n_1398),
.B2(n_1383),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1440),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1471),
.B(n_1388),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1473),
.B(n_1388),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1457),
.B(n_1461),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1445),
.A2(n_1428),
.B1(n_1413),
.B2(n_1414),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1477),
.Y(n_1492)
);

OR2x6_ASAP7_75t_SL g1493 ( 
.A(n_1458),
.B(n_1413),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1478),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1484),
.Y(n_1495)
);

NOR2x1_ASAP7_75t_L g1496 ( 
.A(n_1483),
.B(n_1361),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1466),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1445),
.A2(n_1414),
.B1(n_1419),
.B2(n_1432),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1466),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1476),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1476),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1469),
.Y(n_1502)
);

NOR2xp67_ASAP7_75t_L g1503 ( 
.A(n_1462),
.B(n_1409),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1482),
.B(n_1456),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1470),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1470),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1470),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1472),
.B(n_1362),
.Y(n_1508)
);

NOR2xp67_ASAP7_75t_L g1509 ( 
.A(n_1463),
.B(n_1409),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1467),
.B(n_1362),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1470),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1472),
.B(n_1409),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1454),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1493),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1487),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1509),
.A2(n_1452),
.B(n_1475),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1496),
.B(n_1479),
.Y(n_1517)
);

OAI31xp33_ASAP7_75t_L g1518 ( 
.A1(n_1510),
.A2(n_1442),
.A3(n_1451),
.B(n_1475),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1454),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1505),
.B(n_1452),
.Y(n_1520)
);

OAI322xp33_ASAP7_75t_L g1521 ( 
.A1(n_1505),
.A2(n_1441),
.A3(n_1464),
.B1(n_1474),
.B2(n_1442),
.C1(n_1439),
.C2(n_1459),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1508),
.B(n_1472),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1499),
.B(n_1474),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1494),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1508),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1504),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1508),
.B(n_1488),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1504),
.B(n_1449),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1512),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1486),
.A2(n_1450),
.B1(n_1465),
.B2(n_1437),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1506),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1488),
.B(n_1472),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1494),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1495),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1488),
.B(n_1449),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1512),
.B(n_1460),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1506),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1495),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1507),
.B(n_1511),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1497),
.B(n_1485),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1513),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1513),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1493),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1500),
.B(n_1480),
.Y(n_1545)
);

AND4x1_ASAP7_75t_L g1546 ( 
.A(n_1496),
.B(n_1447),
.C(n_1446),
.D(n_1459),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1500),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1541),
.Y(n_1548)
);

AND2x4_ASAP7_75t_SL g1549 ( 
.A(n_1528),
.B(n_1504),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1514),
.B(n_1502),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1514),
.B(n_1502),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1525),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1524),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1514),
.B(n_1502),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1514),
.B(n_1504),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1526),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1536),
.B(n_1537),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1532),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1524),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1525),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1531),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1546),
.B(n_1465),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1526),
.B(n_1507),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1540),
.B(n_1541),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1531),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1540),
.B(n_1490),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1525),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1547),
.B(n_1511),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1547),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1528),
.B(n_1503),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1481),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1540),
.B(n_1490),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1545),
.B(n_1492),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1542),
.B(n_1501),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1534),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1543),
.B(n_1492),
.Y(n_1577)
);

NAND2x1p5_ASAP7_75t_L g1578 ( 
.A(n_1546),
.B(n_1443),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1535),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_1537),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_1545),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1564),
.B(n_1455),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1581),
.B(n_1533),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1581),
.B(n_1533),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1548),
.B(n_1564),
.Y(n_1585)
);

NAND2x1p5_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1517),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1549),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1557),
.B(n_1544),
.Y(n_1589)
);

NOR2x1_ASAP7_75t_L g1590 ( 
.A(n_1555),
.B(n_1517),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1553),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1566),
.B(n_1538),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1528),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1562),
.B(n_1518),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1566),
.B(n_1538),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1548),
.B(n_1533),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1559),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1549),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1574),
.B(n_1522),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1559),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1573),
.B(n_1538),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1555),
.B(n_1528),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1574),
.B(n_1522),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1552),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1561),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1557),
.B(n_1580),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1561),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1573),
.B(n_1532),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1562),
.B(n_1522),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1552),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1569),
.B(n_1518),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1560),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1555),
.Y(n_1614)
);

NAND2xp33_ASAP7_75t_SL g1615 ( 
.A(n_1563),
.B(n_1526),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1569),
.B(n_1539),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1565),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1569),
.B(n_1539),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1560),
.Y(n_1619)
);

OAI21xp33_ASAP7_75t_L g1620 ( 
.A1(n_1550),
.A2(n_1525),
.B(n_1523),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1565),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1527),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1576),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1586),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1614),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1582),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1596),
.B(n_1577),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1585),
.B(n_1577),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1590),
.B(n_1578),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1588),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1586),
.B(n_1555),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1594),
.B(n_1558),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1597),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1586),
.B(n_1550),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1612),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1597),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1583),
.B(n_1558),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_SL g1638 ( 
.A(n_1614),
.B(n_1521),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1589),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1607),
.B(n_1551),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1598),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1587),
.Y(n_1642)
);

INVxp33_ASAP7_75t_L g1643 ( 
.A(n_1589),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1587),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1610),
.B(n_1571),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1598),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1593),
.B(n_1578),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1608),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1607),
.B(n_1551),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1584),
.A2(n_1530),
.B1(n_1516),
.B2(n_1521),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1608),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1591),
.B(n_1576),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1593),
.B(n_1554),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1621),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1621),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1600),
.A2(n_1530),
.B1(n_1516),
.B2(n_1604),
.Y(n_1656)
);

OAI21xp33_ASAP7_75t_L g1657 ( 
.A1(n_1616),
.A2(n_1568),
.B(n_1554),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1593),
.B(n_1570),
.Y(n_1658)
);

NAND2x1p5_ASAP7_75t_L g1659 ( 
.A(n_1624),
.B(n_1570),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1639),
.B(n_1592),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1633),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1632),
.B(n_1622),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1656),
.A2(n_1613),
.B1(n_1588),
.B2(n_1619),
.C(n_1611),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1626),
.B(n_1599),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1640),
.B(n_1603),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1650),
.A2(n_1578),
.B1(n_1595),
.B2(n_1602),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1632),
.B(n_1592),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1642),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1643),
.A2(n_1578),
.B1(n_1602),
.B2(n_1595),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1635),
.A2(n_1493),
.B1(n_1609),
.B2(n_1599),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1642),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1672)
);

AND2x4_ASAP7_75t_SL g1673 ( 
.A(n_1658),
.B(n_1436),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1625),
.B(n_1622),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1633),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1625),
.B(n_1618),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1640),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1644),
.B(n_1603),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1644),
.Y(n_1679)
);

XNOR2xp5_ASAP7_75t_L g1680 ( 
.A(n_1658),
.B(n_1486),
.Y(n_1680)
);

OAI322xp33_ASAP7_75t_L g1681 ( 
.A1(n_1638),
.A2(n_1520),
.A3(n_1623),
.B1(n_1601),
.B2(n_1617),
.C1(n_1606),
.C2(n_1563),
.Y(n_1681)
);

BUFx2_ASAP7_75t_SL g1682 ( 
.A(n_1624),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1636),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1668),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1665),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1666),
.A2(n_1638),
.B1(n_1634),
.B2(n_1624),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1666),
.A2(n_1657),
.B1(n_1624),
.B2(n_1637),
.C(n_1654),
.Y(n_1687)
);

AOI21xp33_ASAP7_75t_L g1688 ( 
.A1(n_1667),
.A2(n_1630),
.B(n_1636),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1663),
.A2(n_1634),
.B1(n_1631),
.B2(n_1630),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1681),
.A2(n_1657),
.B1(n_1637),
.B2(n_1655),
.C(n_1654),
.Y(n_1690)
);

AOI21xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1670),
.A2(n_1629),
.B(n_1647),
.Y(n_1691)
);

INVxp33_ASAP7_75t_L g1692 ( 
.A(n_1678),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1682),
.B(n_1630),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1661),
.Y(n_1694)
);

O2A1O1Ixp5_ASAP7_75t_L g1695 ( 
.A1(n_1670),
.A2(n_1631),
.B(n_1655),
.C(n_1646),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1660),
.B(n_1628),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1675),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1671),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1683),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1672),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1659),
.A2(n_1572),
.B1(n_1627),
.B2(n_1658),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1679),
.B(n_1658),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1698),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1684),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1700),
.B(n_1677),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1696),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1685),
.B(n_1662),
.Y(n_1707)
);

OA22x2_ASAP7_75t_L g1708 ( 
.A1(n_1686),
.A2(n_1680),
.B1(n_1674),
.B2(n_1669),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1695),
.A2(n_1669),
.B(n_1676),
.C(n_1664),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1691),
.A2(n_1659),
.B1(n_1570),
.B2(n_1645),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1694),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1697),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1689),
.A2(n_1627),
.B1(n_1673),
.B2(n_1646),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1699),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1706),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1703),
.Y(n_1716)
);

OAI21xp33_ASAP7_75t_L g1717 ( 
.A1(n_1710),
.A2(n_1692),
.B(n_1702),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_L g1718 ( 
.A(n_1709),
.B(n_1688),
.C(n_1701),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1704),
.B(n_1687),
.C(n_1690),
.Y(n_1719)
);

NAND4xp25_ASAP7_75t_SL g1720 ( 
.A(n_1705),
.B(n_1653),
.C(n_1649),
.D(n_1651),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1707),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1713),
.B(n_1653),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_L g1723 ( 
.A(n_1713),
.B(n_1648),
.C(n_1641),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_R g1724 ( 
.A(n_1715),
.B(n_1711),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1718),
.A2(n_1714),
.B1(n_1712),
.B2(n_1708),
.C(n_1641),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1719),
.A2(n_1693),
.B1(n_1651),
.B2(n_1648),
.Y(n_1726)
);

AOI21xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1721),
.A2(n_1693),
.B(n_1649),
.Y(n_1727)
);

A2O1A1Ixp33_ASAP7_75t_SL g1728 ( 
.A1(n_1716),
.A2(n_1693),
.B(n_1652),
.C(n_1623),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1726),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1725),
.A2(n_1722),
.B1(n_1717),
.B2(n_1723),
.Y(n_1730)
);

AOI222xp33_ASAP7_75t_L g1731 ( 
.A1(n_1728),
.A2(n_1613),
.B1(n_1605),
.B2(n_1611),
.C1(n_1619),
.C2(n_1720),
.Y(n_1731)
);

AND4x2_ASAP7_75t_L g1732 ( 
.A(n_1727),
.B(n_1615),
.C(n_1652),
.D(n_1556),
.Y(n_1732)
);

AOI322xp5_ASAP7_75t_L g1733 ( 
.A1(n_1724),
.A2(n_1605),
.A3(n_1620),
.B1(n_1529),
.B2(n_1615),
.C1(n_1560),
.C2(n_1567),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1725),
.A2(n_1568),
.B1(n_1520),
.B2(n_1567),
.C(n_1529),
.Y(n_1734)
);

NAND4xp75_ASAP7_75t_L g1735 ( 
.A(n_1729),
.B(n_1503),
.C(n_1444),
.D(n_1438),
.Y(n_1735)
);

NAND4xp75_ASAP7_75t_L g1736 ( 
.A(n_1734),
.B(n_1527),
.C(n_1567),
.D(n_1537),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1730),
.B(n_1603),
.Y(n_1737)
);

XNOR2xp5_ASAP7_75t_L g1738 ( 
.A(n_1732),
.B(n_1468),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1731),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1739),
.B(n_1733),
.C(n_1572),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1738),
.A2(n_1572),
.B1(n_1529),
.B2(n_1520),
.C(n_1556),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1737),
.B(n_1572),
.C(n_1570),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1740),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1742),
.B1(n_1741),
.B2(n_1736),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1744),
.A2(n_1735),
.B1(n_1556),
.B2(n_1579),
.Y(n_1745)
);

XOR2x2_ASAP7_75t_L g1746 ( 
.A(n_1745),
.B(n_1491),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1746),
.Y(n_1747)
);

OAI21xp33_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1556),
.B(n_1572),
.Y(n_1748)
);

AOI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1516),
.B(n_1515),
.Y(n_1749)
);

NOR2xp67_ASAP7_75t_SL g1750 ( 
.A(n_1749),
.B(n_1433),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_R g1751 ( 
.A1(n_1750),
.A2(n_1498),
.B1(n_1579),
.B2(n_1491),
.C(n_1575),
.Y(n_1751)
);

AOI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1453),
.B(n_1519),
.C(n_1523),
.Y(n_1752)
);


endmodule