module fake_jpeg_4227_n_189 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_31),
.B(n_2),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_50),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_46),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_22),
.B1(n_14),
.B2(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_64),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_22),
.B1(n_14),
.B2(n_20),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_59),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_14),
.B1(n_25),
.B2(n_20),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_18),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_69),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_29),
.C(n_18),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_68),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_29),
.C(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_23),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_70),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_76),
.B(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_84),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_65),
.B1(n_67),
.B2(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_10),
.C(n_13),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_58),
.B1(n_11),
.B2(n_12),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_21),
.B1(n_24),
.B2(n_6),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_120)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_48),
.B(n_45),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_83),
.B(n_78),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_49),
.C(n_59),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_91),
.B(n_93),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_51),
.C(n_66),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.C(n_78),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_82),
.C(n_90),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2x1_ASAP7_75t_R g119 ( 
.A(n_83),
.B(n_72),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_76),
.B(n_87),
.C(n_97),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_87),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_72),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_11),
.B1(n_9),
.B2(n_8),
.Y(n_122)
);

BUFx12f_ASAP7_75t_SL g123 ( 
.A(n_119),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_139),
.B(n_111),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_134),
.C(n_111),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_131),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_83),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_102),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_46),
.B(n_100),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_101),
.B(n_79),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_106),
.B1(n_105),
.B2(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_125),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_146),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_113),
.B(n_116),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_147),
.B(n_150),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_151),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_86),
.B(n_114),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_96),
.B1(n_107),
.B2(n_103),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_146),
.Y(n_168)
);

OAI31xp33_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_130),
.A3(n_132),
.B(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_162),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_132),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_163),
.C(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_127),
.B1(n_144),
.B2(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_167),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_161),
.C(n_155),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_144),
.B1(n_145),
.B2(n_129),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_171),
.B(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_142),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_175),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_178),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_168),
.C(n_172),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_133),
.B(n_81),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_180),
.B(n_182),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_165),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_186),
.B(n_183),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_86),
.A3(n_174),
.B1(n_112),
.B2(n_107),
.C(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_117),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);


endmodule