module fake_jpeg_22566_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_0),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_19),
.B1(n_15),
.B2(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_19),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_13),
.B1(n_14),
.B2(n_24),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_18),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_48),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_52),
.B(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_60),
.B1(n_63),
.B2(n_36),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_28),
.B(n_15),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_57),
.B(n_58),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_28),
.B(n_16),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_30),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_64),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_28),
.B1(n_27),
.B2(n_16),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_14),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_69),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_39),
.B(n_47),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_71),
.B(n_60),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_34),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_74),
.B(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_36),
.B1(n_50),
.B2(n_49),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_79),
.B1(n_61),
.B2(n_55),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_49),
.C(n_51),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_73),
.B1(n_68),
.B2(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_87),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_83),
.A2(n_73),
.B1(n_56),
.B2(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_85),
.B1(n_21),
.B2(n_10),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_85),
.B(n_86),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_R g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_91),
.B1(n_7),
.B2(n_11),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_93),
.B(n_5),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_5),
.C(n_7),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_99),
.Y(n_101)
);


endmodule