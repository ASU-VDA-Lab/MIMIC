module real_jpeg_29444_n_17 (n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_323;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_0),
.A2(n_35),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_0),
.A2(n_46),
.B1(n_101),
.B2(n_102),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_0),
.A2(n_46),
.B1(n_159),
.B2(n_160),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

A2O1A1O1Ixp25_ASAP7_75t_L g39 ( 
.A1(n_1),
.A2(n_36),
.B(n_37),
.C(n_40),
.D(n_44),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_1),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_62),
.B(n_66),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_101),
.B(n_103),
.C(n_104),
.D(n_106),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_1),
.B(n_101),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_1),
.B(n_132),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_134),
.B(n_158),
.C(n_159),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_1),
.A2(n_83),
.B1(n_159),
.B2(n_160),
.Y(n_167)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_3),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_156),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_3),
.A2(n_101),
.B1(n_102),
.B2(n_156),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_3),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_301)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_5),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_5),
.A2(n_35),
.B1(n_37),
.B2(n_219),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_5),
.A2(n_101),
.B1(n_102),
.B2(n_219),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_5),
.A2(n_159),
.B1(n_160),
.B2(n_219),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_35),
.B1(n_37),
.B2(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_58),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_7),
.A2(n_58),
.B1(n_101),
.B2(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_7),
.A2(n_58),
.B1(n_159),
.B2(n_160),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_8),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_8),
.A2(n_35),
.B1(n_37),
.B2(n_116),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_8),
.A2(n_101),
.B1(n_102),
.B2(n_116),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_8),
.A2(n_116),
.B1(n_159),
.B2(n_160),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_35),
.B1(n_37),
.B2(n_65),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_65),
.B1(n_101),
.B2(n_102),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_10),
.A2(n_65),
.B1(n_159),
.B2(n_160),
.Y(n_212)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_11),
.B(n_37),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_12),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_12),
.A2(n_35),
.B1(n_37),
.B2(n_201),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_12),
.A2(n_101),
.B1(n_102),
.B2(n_201),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_12),
.A2(n_159),
.B1(n_160),
.B2(n_201),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_13),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_138),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_13),
.A2(n_101),
.B1(n_102),
.B2(n_138),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_13),
.A2(n_138),
.B1(n_159),
.B2(n_160),
.Y(n_291)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_15),
.A2(n_53),
.B1(n_101),
.B2(n_102),
.Y(n_105)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_333),
.B(n_336),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_328),
.B(n_332),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_315),
.B(n_327),
.Y(n_19)
);

OAI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_279),
.A3(n_308),
.B1(n_313),
.B2(n_314),
.C(n_340),
.Y(n_20)
);

AOI321xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_229),
.A3(n_268),
.B1(n_273),
.B2(n_278),
.C(n_341),
.Y(n_21)
);

NOR3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_180),
.C(n_225),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_147),
.B(n_179),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_121),
.B(n_146),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_96),
.B(n_120),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_70),
.B(n_95),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_48),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_28),
.B(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_39),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_39),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.A3(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_30),
.B(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_31),
.B(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_35),
.B(n_54),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_37),
.A2(n_102),
.A3(n_103),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_40),
.A2(n_43),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_40),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_40),
.A2(n_43),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_40),
.A2(n_43),
.B1(n_245),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_44),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_57),
.B(n_59),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_47),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_47),
.A2(n_59),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_47),
.A2(n_143),
.B1(n_178),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_47),
.A2(n_143),
.B1(n_203),
.B2(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_47),
.A2(n_143),
.B(n_254),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_61),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_56),
.C(n_61),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_52),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_52),
.A2(n_104),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_52),
.A2(n_104),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_52),
.A2(n_104),
.B1(n_257),
.B2(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_52),
.A2(n_104),
.B(n_320),
.Y(n_319)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B(n_66),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_62),
.A2(n_115),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_62),
.A2(n_78),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_62),
.A2(n_78),
.B1(n_200),
.B2(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_62),
.A2(n_78),
.B(n_218),
.Y(n_247)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_74),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_86),
.B(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_SL g139 ( 
.A(n_69),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_69),
.A2(n_75),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_80),
.B(n_94),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_79),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_93),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_83),
.A2(n_101),
.B(n_133),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_98),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_109),
.C(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_102),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_108),
.A2(n_127),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_108),
.A2(n_188),
.B1(n_215),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_108),
.A2(n_188),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_123),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_140),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_141),
.C(n_142),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_130),
.C(n_136),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_126),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_132),
.A2(n_165),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_132),
.A2(n_165),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_132),
.A2(n_165),
.B1(n_323),
.B2(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_132),
.A2(n_165),
.B(n_330),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_134),
.B1(n_159),
.B2(n_160),
.Y(n_166)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_149),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_163),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_151),
.B(n_152),
.C(n_163),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_161),
.Y(n_184)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_173),
.C(n_176),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B(n_168),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_165),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_169),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_181),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_205),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_182),
.B(n_205),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_197),
.C(n_204),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_186),
.C(n_196),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_196),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B(n_190),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_191),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_194),
.B(n_195),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_194),
.A2(n_195),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_194),
.A2(n_236),
.B1(n_264),
.B2(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_194),
.A2(n_236),
.B1(n_291),
.B2(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_204),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_202),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_216),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_207),
.B(n_216),
.C(n_224),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_220),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_226),
.B(n_227),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_249),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_241),
.C(n_248),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_241),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_240),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_232),
.Y(n_240)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_238),
.C(n_240),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_247),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_247),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_247),
.A2(n_262),
.B(n_265),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_267),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_259),
.B1(n_260),
.B2(n_266),
.Y(n_250)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_255),
.B(n_258),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_255),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_258),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_281),
.B1(n_282),
.B2(n_293),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_259),
.B(n_266),
.C(n_267),
.Y(n_309)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_274),
.B(n_277),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_270),
.B(n_271),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_296),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_296),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_293),
.C(n_294),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_290),
.B2(n_292),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_285),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_289),
.C(n_290),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_286),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_287),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_289),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_300),
.C(n_304),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_290),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_292),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_299),
.C(n_307),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_294),
.A2(n_295),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_307),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_301),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_317),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_326),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_319),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_321),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_325),
.C(n_326),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_329),
.B(n_331),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_329),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);


endmodule