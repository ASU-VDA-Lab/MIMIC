module fake_jpeg_1367_n_152 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx6p67_ASAP7_75t_R g74 ( 
.A(n_33),
.Y(n_74)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_28),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_8),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_43),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_11),
.B(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_47),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_9),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_10),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_55),
.B(n_80),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_80),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_75),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_23),
.B1(n_14),
.B2(n_4),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_45),
.C(n_48),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_74),
.Y(n_98)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_38),
.A2(n_23),
.B1(n_39),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_59),
.B1(n_74),
.B2(n_67),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_47),
.B(n_41),
.C(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_92),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_42),
.B1(n_49),
.B2(n_81),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_86),
.B1(n_96),
.B2(n_87),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_76),
.B1(n_61),
.B2(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_69),
.B1(n_67),
.B2(n_60),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_96),
.B(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_64),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_78),
.B1(n_68),
.B2(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_58),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_72),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_83),
.B(n_97),
.Y(n_102)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_113),
.B1(n_102),
.B2(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_91),
.B1(n_84),
.B2(n_82),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_110),
.B1(n_113),
.B2(n_112),
.Y(n_124)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_104),
.Y(n_118)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_123),
.C(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_127),
.B1(n_115),
.B2(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_126),
.B(n_121),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_103),
.B1(n_115),
.B2(n_110),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_109),
.B(n_106),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_117),
.B(n_120),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_107),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_133),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_127),
.C(n_122),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_131),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_117),
.CI(n_120),
.CON(n_137),
.SN(n_137)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_137),
.B(n_135),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_139),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_142),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_129),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_134),
.Y(n_143)
);

AOI21x1_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_136),
.B(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_144),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_146),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_132),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_149),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_148),
.Y(n_152)
);


endmodule