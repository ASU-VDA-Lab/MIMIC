module fake_jpeg_11452_n_529 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_529);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_529;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_51),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_52),
.B(n_68),
.Y(n_144)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_61),
.B(n_64),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_18),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_65),
.Y(n_140)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_0),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_70),
.B(n_75),
.Y(n_150)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_85),
.B(n_87),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_89),
.Y(n_154)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_26),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_0),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_34),
.B(n_0),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_26),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_36),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_96),
.B(n_97),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_27),
.Y(n_97)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

AND2x4_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_27),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_23),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_65),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_73),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_36),
.B1(n_49),
.B2(n_47),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_112),
.A2(n_155),
.B1(n_54),
.B2(n_74),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_62),
.B1(n_92),
.B2(n_84),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_113),
.A2(n_115),
.B1(n_116),
.B2(n_123),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_60),
.A2(n_37),
.B1(n_40),
.B2(n_29),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_114),
.A2(n_121),
.B1(n_122),
.B2(n_151),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_27),
.B1(n_29),
.B2(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_68),
.A2(n_50),
.B1(n_38),
.B2(n_37),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_50),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_126),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_29),
.B1(n_45),
.B2(n_30),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_63),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_46),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_146),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_77),
.A2(n_29),
.B1(n_41),
.B2(n_43),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_135),
.A2(n_8),
.B(n_9),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_30),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_100),
.A2(n_45),
.B1(n_30),
.B2(n_23),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_94),
.A2(n_30),
.B1(n_23),
.B2(n_45),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_72),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_95),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_67),
.A2(n_30),
.B1(n_23),
.B2(n_43),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_162),
.B1(n_54),
.B2(n_5),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_67),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_164),
.B(n_166),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_165),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_75),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_129),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_175),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_108),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_173),
.A2(n_131),
.B1(n_135),
.B2(n_116),
.Y(n_222)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_176),
.B(n_191),
.Y(n_254)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_93),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_129),
.Y(n_180)
);

NAND2xp33_ASAP7_75t_SL g259 ( 
.A(n_180),
.B(n_186),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_78),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_181),
.B(n_188),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_73),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_76),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_129),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_127),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_2),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_3),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_126),
.B(n_98),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_58),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_194),
.A2(n_160),
.B(n_124),
.Y(n_257)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_198),
.A2(n_203),
.B1(n_219),
.B2(n_221),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_124),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_202),
.Y(n_246)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_200),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_124),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_109),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_7),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_216),
.Y(n_230)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_105),
.B(n_7),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_208),
.B(n_213),
.Y(n_264)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_209),
.Y(n_262)
);

INVx11_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

BUFx24_ASAP7_75t_L g255 ( 
.A(n_210),
.Y(n_255)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_212),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_140),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_111),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_214),
.Y(n_253)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_111),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_146),
.B(n_7),
.C(n_8),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_109),
.C(n_124),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_117),
.B1(n_145),
.B2(n_118),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_8),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_220),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_222),
.A2(n_233),
.B1(n_239),
.B2(n_263),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_226),
.B(n_266),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_107),
.B1(n_134),
.B2(n_110),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_228),
.A2(n_176),
.B1(n_184),
.B2(n_182),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_171),
.B1(n_178),
.B2(n_169),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_134),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_238),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_107),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_191),
.A2(n_120),
.B1(n_153),
.B2(n_110),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_131),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_SL g245 ( 
.A(n_194),
.B(n_117),
.C(n_145),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_176),
.C(n_257),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_257),
.B(n_125),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_191),
.A2(n_102),
.B1(n_120),
.B2(n_142),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_153),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_186),
.B1(n_180),
.B2(n_200),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_273),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_254),
.B(n_244),
.C(n_270),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_291),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_185),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_275),
.B(n_276),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_230),
.B(n_182),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_225),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_283),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_279),
.A2(n_301),
.B(n_309),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_280),
.A2(n_286),
.B1(n_290),
.B2(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_179),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_232),
.B(n_194),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_285),
.B(n_296),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_228),
.A2(n_218),
.B1(n_184),
.B2(n_142),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_179),
.B1(n_216),
.B2(n_209),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_288),
.A2(n_295),
.B1(n_308),
.B2(n_311),
.Y(n_361)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_243),
.A2(n_136),
.B1(n_147),
.B2(n_196),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_230),
.B(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_229),
.Y(n_292)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_246),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_294),
.B(n_299),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_254),
.B1(n_235),
.B2(n_239),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_258),
.B(n_174),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_214),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_297),
.B(n_259),
.Y(n_324)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_298),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_167),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_163),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_313),
.C(n_249),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_302),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_219),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_303),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_211),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_269),
.Y(n_332)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_305),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_226),
.B(n_204),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_306),
.A2(n_307),
.B(n_317),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_247),
.B(n_205),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_263),
.A2(n_136),
.B1(n_147),
.B2(n_195),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_231),
.B(n_172),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

NOR2x1_ASAP7_75t_R g352 ( 
.A(n_310),
.B(n_314),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_261),
.A2(n_189),
.B1(n_103),
.B2(n_193),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_255),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_312),
.A2(n_315),
.B(n_316),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_165),
.C(n_212),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_255),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_237),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_240),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_245),
.B(n_125),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_318),
.A2(n_255),
.B(n_210),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_240),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_320),
.B(n_12),
.C(n_13),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_281),
.A2(n_265),
.B1(n_251),
.B2(n_267),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_322),
.A2(n_330),
.B1(n_339),
.B2(n_315),
.Y(n_381)
);

XNOR2x1_ASAP7_75t_L g392 ( 
.A(n_324),
.B(n_331),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_281),
.A2(n_251),
.B1(n_183),
.B2(n_170),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_287),
.B(n_247),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_354),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_334),
.B(n_298),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_286),
.A2(n_271),
.B1(n_256),
.B2(n_250),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_340),
.B1(n_345),
.B2(n_348),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_278),
.B(n_269),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_350),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_295),
.A2(n_187),
.B1(n_256),
.B2(n_250),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_280),
.A2(n_224),
.B1(n_227),
.B2(n_252),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_342),
.B(n_354),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_306),
.A2(n_224),
.B1(n_252),
.B2(n_253),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_318),
.A2(n_249),
.B(n_241),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_346),
.A2(n_301),
.B(n_285),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_260),
.C(n_236),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_349),
.C(n_351),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_284),
.A2(n_234),
.B1(n_241),
.B2(n_236),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_149),
.C(n_234),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_278),
.B(n_125),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_284),
.B(n_207),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_299),
.A2(n_149),
.B(n_177),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_274),
.B(n_9),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_301),
.C(n_276),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_279),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_359),
.A2(n_312),
.B1(n_292),
.B2(n_282),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_360),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_368),
.Y(n_402)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_304),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_366),
.B(n_369),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_297),
.Y(n_368)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_351),
.B(n_288),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_329),
.A2(n_291),
.B1(n_308),
.B2(n_296),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_371),
.A2(n_381),
.B1(n_386),
.B2(n_387),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_333),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_374),
.Y(n_409)
);

BUFx12_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_377),
.Y(n_400)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_328),
.B(n_307),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_378),
.A2(n_383),
.B1(n_357),
.B2(n_339),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_289),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_385),
.C(n_350),
.Y(n_397)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_384),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_329),
.A2(n_317),
.B1(n_316),
.B2(n_314),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_336),
.A2(n_310),
.B(n_305),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_322),
.A2(n_290),
.B1(n_293),
.B2(n_309),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_361),
.A2(n_309),
.B1(n_302),
.B2(n_12),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_328),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_388),
.A2(n_390),
.B1(n_393),
.B2(n_394),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_357),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_389),
.B(n_391),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_10),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_11),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_17),
.B1(n_13),
.B2(n_14),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_335),
.B1(n_343),
.B2(n_323),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_359),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_398),
.C(n_406),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_347),
.C(n_326),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_403),
.A2(n_367),
.B1(n_380),
.B2(n_376),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_405),
.B(n_396),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_325),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_326),
.C(n_320),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_408),
.C(n_412),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_331),
.C(n_338),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_325),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_410),
.B(n_330),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_349),
.C(n_355),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_332),
.C(n_324),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_418),
.C(n_419),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_381),
.A2(n_337),
.B1(n_348),
.B2(n_327),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_371),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_346),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_342),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_344),
.C(n_340),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_423),
.C(n_424),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_327),
.C(n_353),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_353),
.C(n_354),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_363),
.B(n_345),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_383),
.C(n_384),
.Y(n_442)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_426),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_442),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_436),
.Y(n_455)
);

AO22x1_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_378),
.B1(n_363),
.B2(n_389),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_432),
.A2(n_448),
.B(n_423),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_402),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_433),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_372),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_434),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_362),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_435),
.B(n_446),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_403),
.A2(n_394),
.B1(n_387),
.B2(n_422),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_368),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_443),
.A2(n_447),
.B(n_416),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_400),
.A2(n_386),
.B1(n_391),
.B2(n_395),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_445),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_SL g448 ( 
.A(n_407),
.B(n_382),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_398),
.B(n_408),
.C(n_397),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_452),
.C(n_412),
.Y(n_453)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

INVx11_ASAP7_75t_L g471 ( 
.A(n_450),
.Y(n_471)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

NOR3xp33_ASAP7_75t_SL g468 ( 
.A(n_451),
.B(n_375),
.C(n_393),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_459),
.C(n_437),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_450),
.A2(n_401),
.B(n_420),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_456),
.A2(n_460),
.B(n_438),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_442),
.A2(n_425),
.B(n_419),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_461),
.A2(n_463),
.B(n_443),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_406),
.C(n_418),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_469),
.C(n_470),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_443),
.A2(n_375),
.B(n_410),
.Y(n_463)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_445),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_472),
.Y(n_487)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_468),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_413),
.C(n_405),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_364),
.C(n_323),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_343),
.C(n_335),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_477),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_459),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_478),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_438),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_461),
.A2(n_451),
.B1(n_429),
.B2(n_428),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_479),
.A2(n_457),
.B1(n_443),
.B2(n_455),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_456),
.A2(n_449),
.B(n_437),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_480),
.A2(n_455),
.B(n_471),
.Y(n_501)
);

XNOR2x1_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_452),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_482),
.C(n_453),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_462),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_486),
.Y(n_492)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_465),
.Y(n_495)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_463),
.B(n_432),
.CI(n_433),
.CON(n_485),
.SN(n_485)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_486),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_447),
.Y(n_486)
);

OAI221xp5_ASAP7_75t_L g488 ( 
.A1(n_473),
.A2(n_430),
.B1(n_432),
.B2(n_439),
.C(n_440),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_488),
.A2(n_465),
.B1(n_458),
.B2(n_471),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_499),
.B(n_501),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_489),
.B(n_472),
.C(n_470),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_494),
.B(n_497),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_474),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_496),
.A2(n_478),
.B(n_483),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_464),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_464),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_498),
.B(n_494),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_469),
.C(n_457),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_500),
.A2(n_503),
.B1(n_477),
.B2(n_485),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_475),
.A2(n_471),
.B(n_468),
.Y(n_503)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_479),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_509),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g510 ( 
.A1(n_492),
.A2(n_482),
.B(n_485),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_510),
.B(n_511),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_493),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_481),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_502),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_502),
.C(n_492),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_518),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_516),
.A2(n_490),
.B(n_509),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_520),
.Y(n_524)
);

AOI321xp33_ASAP7_75t_L g525 ( 
.A1(n_521),
.A2(n_523),
.A3(n_519),
.B1(n_515),
.B2(n_500),
.C(n_375),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_517),
.A2(n_512),
.B(n_505),
.Y(n_523)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_525),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_522),
.B(n_524),
.Y(n_527)
);

AOI221xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_12),
.B1(n_16),
.B2(n_17),
.C(n_515),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_12),
.Y(n_529)
);


endmodule