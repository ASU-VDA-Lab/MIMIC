module fake_jpeg_3433_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_47),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_53),
.Y(n_59)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_62),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_56),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_42),
.B1(n_41),
.B2(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_43),
.B1(n_45),
.B2(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_41),
.B1(n_46),
.B2(n_44),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_43),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_52),
.B(n_49),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_87),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_63),
.B1(n_61),
.B2(n_44),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_84),
.B1(n_88),
.B2(n_4),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_66),
.B(n_68),
.C(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_55),
.B1(n_52),
.B2(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_21),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_1),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_74),
.B(n_2),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_103),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_73),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_104),
.B(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_101),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_45),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_2),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_45),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_107),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_96),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_23),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_86),
.B(n_81),
.C(n_24),
.D(n_26),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_14),
.C(n_15),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_20),
.B1(n_38),
.B2(n_37),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_8),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_19),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_29),
.B1(n_36),
.B2(n_35),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_9),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_100),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_107),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_138),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_14),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_109),
.B1(n_129),
.B2(n_128),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_110),
.B1(n_123),
.B2(n_108),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_138),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_148),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_130),
.C(n_136),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_139),
.B(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_147),
.B1(n_139),
.B2(n_130),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_120),
.B(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_149),
.B1(n_137),
.B2(n_135),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_30),
.B(n_31),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_32),
.C(n_34),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_39),
.Y(n_158)
);


endmodule