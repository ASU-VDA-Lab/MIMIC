module real_jpeg_29668_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_288;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_299;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_0),
.B(n_52),
.Y(n_84)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_0),
.B(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_0),
.B(n_230),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_30),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_46),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_57),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_21),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_2),
.A2(n_10),
.B(n_46),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_2),
.A2(n_51),
.B(n_53),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_63),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_32),
.B1(n_46),
.B2(n_49),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_4),
.A2(n_32),
.B1(n_51),
.B2(n_52),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_6),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_135),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_6),
.A2(n_46),
.B1(n_49),
.B2(n_135),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_135),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_7),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_46),
.B1(n_49),
.B2(n_67),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_67),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_51),
.B1(n_52),
.B2(n_67),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_11),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_110),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_109),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_16),
.B(n_92),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_71),
.C(n_79),
.Y(n_16)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_17),
.B(n_71),
.CI(n_79),
.CON(n_141),
.SN(n_141)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_18),
.A2(n_19),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_19),
.B(n_41),
.C(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_20),
.B(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_21),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_23),
.B(n_30),
.C(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_22),
.A2(n_35),
.B(n_37),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_22),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_24),
.B(n_27),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_25),
.B(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_25),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_25),
.A2(n_57),
.B(n_195),
.C(n_196),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_29),
.B(n_35),
.Y(n_99)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_34),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_35),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_36),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_37),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_38),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_58),
.B2(n_59),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_41),
.B(n_155),
.C(n_157),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_41),
.A2(n_42),
.B1(n_157),
.B2(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_54),
.B(n_55),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_44),
.B(n_56),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_44),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_49),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_46),
.A2(n_48),
.B(n_57),
.C(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_50),
.B(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_50),
.B(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_52),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_54),
.A2(n_77),
.B(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_54),
.B(n_57),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_57),
.B(n_86),
.Y(n_245)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B(n_68),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_60),
.B(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_60),
.B(n_160),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_60),
.Y(n_276)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_63),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_69),
.B(n_168),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_73),
.A2(n_104),
.B(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_76),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_77),
.B(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_91),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_81),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_82),
.A2(n_83),
.B1(n_91),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_82),
.A2(n_83),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_83),
.B(n_194),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_87),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_84),
.B(n_87),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_84),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_87),
.Y(n_117)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_85),
.Y(n_175)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_88),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_90),
.B(n_212),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_91),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_108),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_107),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_99),
.B(n_156),
.Y(n_273)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_103),
.B(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_142),
.B(n_299),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_141),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_112),
.B(n_141),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_136),
.C(n_137),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_113),
.A2(n_114),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.C(n_127),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_115),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_116),
.B(n_123),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_117),
.B(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_118),
.A2(n_150),
.B(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_119),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_124),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_126),
.B(n_159),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_136),
.B(n_137),
.Y(n_297)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_141),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_293),
.B(n_298),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_280),
.B(n_292),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_188),
.B(n_263),
.C(n_279),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_176),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_146),
.B(n_176),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_161),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_148),
.B(n_154),
.C(n_161),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_149),
.B(n_152),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_151),
.B(n_229),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_153),
.B(n_202),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_169),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_163),
.B(n_166),
.C(n_169),
.Y(n_277)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.C(n_182),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_177),
.A2(n_178),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_262),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_255),
.B(n_261),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_214),
.B(n_254),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_204),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_192),
.B(n_204),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.C(n_200),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_193),
.B(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_194),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_252)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_211),
.C(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_249),
.B(n_253),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_231),
.B(n_248),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_238),
.B(n_247),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_236),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_242),
.B(n_246),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_251),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_256),
.B(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_277),
.B2(n_278),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_269),
.C(n_278),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_273),
.C(n_274),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_291),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_288),
.B2(n_289),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_289),
.C(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);


endmodule