module fake_jpeg_24669_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_25),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_57),
.Y(n_107)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_67),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_34),
.B1(n_30),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_66),
.B1(n_83),
.B2(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_70),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_32),
.B1(n_23),
.B2(n_28),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

CKINVDCx6p67_ASAP7_75t_R g81 ( 
.A(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_81),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_24),
.B(n_36),
.C(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_35),
.B1(n_28),
.B2(n_36),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_59),
.Y(n_118)
);

OR2x6_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_24),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_103),
.B(n_81),
.Y(n_122)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_3),
.Y(n_148)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_61),
.B(n_24),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_24),
.C(n_27),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_115),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_25),
.B1(n_21),
.B2(n_19),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_67),
.B1(n_76),
.B2(n_51),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_118),
.B(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_120),
.B(n_121),
.Y(n_173)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_105),
.B(n_116),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_95),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_85),
.B(n_19),
.C(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_73),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_132),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_136),
.B1(n_137),
.B2(n_99),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_139),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_84),
.B1(n_51),
.B2(n_68),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_68),
.B1(n_53),
.B2(n_65),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_2),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_16),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_2),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_65),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_161),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_106),
.C(n_90),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_158),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_103),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_138),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_99),
.B1(n_90),
.B2(n_116),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_112),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_127),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_176),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_144),
.B(n_140),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_89),
.B1(n_98),
.B2(n_93),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_182),
.B(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_119),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_187),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_137),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_196),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_133),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_156),
.B(n_157),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_191),
.B(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_152),
.A2(n_120),
.B(n_121),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_98),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_154),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_199),
.C(n_205),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_175),
.C(n_153),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_131),
.B1(n_150),
.B2(n_169),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_179),
.B1(n_213),
.B2(n_186),
.Y(n_223)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_191),
.B1(n_184),
.B2(n_178),
.C(n_196),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_161),
.C(n_163),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_171),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_186),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_151),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_190),
.B(n_183),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_212),
.B(n_213),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_196),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_199),
.B1(n_203),
.B2(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_207),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_201),
.B1(n_204),
.B2(n_211),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_179),
.B1(n_177),
.B2(n_151),
.Y(n_224)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

BUFx12f_ASAP7_75t_SL g225 ( 
.A(n_201),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

OA21x2_ASAP7_75t_SL g226 ( 
.A1(n_214),
.A2(n_172),
.B(n_159),
.Y(n_226)
);

OAI322xp33_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_166),
.A3(n_93),
.B1(n_149),
.B2(n_128),
.C1(n_16),
.C2(n_15),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_177),
.B1(n_193),
.B2(n_173),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_162),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_236),
.Y(n_245)
);

AOI31xp67_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_201),
.A3(n_202),
.B(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_235),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_215),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_228),
.B1(n_221),
.B2(n_224),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_238),
.A2(n_14),
.B(n_165),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_244),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_216),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_247),
.B(n_237),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_166),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_149),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_248),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_254),
.C(n_155),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_232),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_240),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_233),
.A3(n_236),
.B1(n_232),
.B2(n_230),
.C1(n_215),
.C2(n_222),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_218),
.Y(n_255)
);

OAI211xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_256),
.B(n_5),
.C(n_6),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_162),
.B1(n_89),
.B2(n_155),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_258),
.C(n_4),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_155),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_4),
.C(n_5),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_4),
.C(n_6),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_262),
.Y(n_265)
);


endmodule