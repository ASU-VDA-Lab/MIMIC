module fake_jpeg_4789_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_240;
wire n_131;
wire n_56;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_19),
.B1(n_25),
.B2(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_47),
.B1(n_58),
.B2(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_19),
.B1(n_25),
.B2(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_55),
.Y(n_73)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_22),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_17),
.B1(n_18),
.B2(n_24),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_32),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_63),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_29),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_14),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_10),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_39),
.B(n_38),
.C(n_43),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_69),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_71),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_38),
.B1(n_39),
.B2(n_32),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_85),
.B1(n_60),
.B2(n_51),
.Y(n_107)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_29),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_45),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_29),
.C(n_27),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_88),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_29),
.C(n_26),
.Y(n_88)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_14),
.B(n_13),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_50),
.CI(n_59),
.CON(n_101),
.SN(n_101)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_101),
.B(n_116),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_105),
.Y(n_142)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_108),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_60),
.B1(n_51),
.B2(n_47),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_56),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_45),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_54),
.Y(n_130)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_72),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_70),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_58),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_123),
.A2(n_149),
.B(n_13),
.Y(n_179)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_129),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_81),
.B(n_46),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_127),
.A2(n_148),
.B(n_53),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_98),
.Y(n_156)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_133),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_75),
.B1(n_91),
.B2(n_78),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_136),
.B1(n_143),
.B2(n_102),
.Y(n_164)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_140),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_83),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_147),
.C(n_141),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_88),
.B1(n_87),
.B2(n_77),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_69),
.B(n_67),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_112),
.B(n_99),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_65),
.C(n_63),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_145),
.C(n_101),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_66),
.B1(n_77),
.B2(n_70),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_49),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_102),
.B1(n_120),
.B2(n_97),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_49),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_119),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_44),
.B(n_54),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_101),
.A2(n_98),
.B1(n_104),
.B2(n_99),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_158),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_98),
.C(n_112),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_156),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_168),
.B(n_180),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_100),
.C(n_118),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_166),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_165),
.B1(n_143),
.B2(n_137),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_125),
.A2(n_102),
.B1(n_108),
.B2(n_100),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_136),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_173),
.Y(n_203)
);

OAI22x1_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_94),
.B1(n_53),
.B2(n_54),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_171),
.A2(n_131),
.B1(n_148),
.B2(n_129),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_61),
.C(n_53),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_174),
.Y(n_206)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_44),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_89),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_124),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_0),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_105),
.B1(n_9),
.B2(n_10),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_140),
.B(n_134),
.Y(n_191)
);

XOR2x1_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_126),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_149),
.B1(n_125),
.B2(n_127),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_189),
.B1(n_191),
.B2(n_200),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_128),
.B(n_123),
.C(n_124),
.D(n_144),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_174),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_171),
.B1(n_176),
.B2(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_193),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_187),
.A2(n_199),
.B1(n_0),
.B2(n_1),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_144),
.B(n_138),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_198),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_170),
.B(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_128),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_153),
.A2(n_89),
.B1(n_137),
.B2(n_96),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_199),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_158),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_213),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_180),
.C(n_152),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_210),
.C(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_172),
.C(n_177),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_159),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_161),
.C(n_162),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_161),
.C(n_157),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_222),
.C(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_164),
.B1(n_193),
.B2(n_165),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_203),
.B1(n_186),
.B2(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_166),
.C(n_173),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_183),
.B(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_224),
.B(n_187),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_137),
.C(n_89),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_191),
.B(n_203),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_205),
.C(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_228),
.C(n_185),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_0),
.C(n_1),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_184),
.B(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_237),
.Y(n_254)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_235),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_241),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_244),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_182),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_243),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_210),
.C(n_208),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_220),
.B1(n_201),
.B2(n_12),
.Y(n_255)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_243),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_256),
.B(n_258),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_212),
.B1(n_213),
.B2(n_209),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_245),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_236),
.B1(n_12),
.B2(n_11),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_1),
.C(n_2),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_1),
.C(n_2),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_12),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_238),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_230),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_257),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_268),
.C(n_270),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_239),
.B1(n_231),
.B2(n_247),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_272),
.B1(n_262),
.B2(n_258),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_248),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_269),
.B(n_271),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_261),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_267),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_237),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_252),
.A2(n_233),
.B1(n_245),
.B2(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_255),
.B(n_11),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_284),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_2),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_254),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_280),
.A2(n_278),
.B(n_277),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_256),
.B(n_252),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_3),
.C(n_4),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_259),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_286),
.B(n_287),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_11),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_288),
.A2(n_6),
.B1(n_7),
.B2(n_290),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_3),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_5),
.Y(n_294)
);

AOI31xp67_ASAP7_75t_SL g292 ( 
.A1(n_291),
.A2(n_283),
.A3(n_4),
.B(n_5),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_282),
.C2(n_266),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_296),
.C(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_298),
.Y(n_301)
);


endmodule