module real_jpeg_26868_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_0),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_0),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_0),
.A2(n_54),
.B1(n_56),
.B2(n_75),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_75),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_75),
.Y(n_212)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_1),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_37),
.B1(n_70),
.B2(n_71),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_37),
.B1(n_54),
.B2(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_2),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_3),
.A2(n_34),
.B1(n_54),
.B2(n_56),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_70),
.B1(n_71),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_7),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_7),
.A2(n_54),
.B1(n_56),
.B2(n_132),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_132),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_225)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_9),
.B(n_73),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_56),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_9),
.A2(n_56),
.B(n_176),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_121),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_9),
.A2(n_28),
.B(n_43),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_9),
.B(n_57),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_9),
.A2(n_31),
.B1(n_82),
.B2(n_225),
.Y(n_228)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_70),
.B1(n_71),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_12),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_12),
.A2(n_54),
.B1(n_56),
.B2(n_107),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_107),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_107),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_13),
.A2(n_47),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_14),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_63)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_14),
.Y(n_175)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_19),
.B(n_109),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_90),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_78),
.B2(n_79),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_38),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_25),
.A2(n_83),
.B(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_26),
.A2(n_36),
.B(n_95),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_26),
.A2(n_30),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_27),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_30),
.Y(n_226)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_31),
.A2(n_82),
.B1(n_93),
.B2(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_33),
.B(n_83),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_35),
.A2(n_82),
.B(n_212),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_39),
.A2(n_48),
.B(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_39),
.A2(n_86),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_39),
.A2(n_45),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_39),
.A2(n_184),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_39),
.A2(n_45),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_39),
.A2(n_45),
.B1(n_183),
.B2(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_41),
.A2(n_54),
.A3(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_42),
.B(n_174),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_42),
.A2(n_44),
.B(n_121),
.C(n_204),
.Y(n_203)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_46),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_45),
.B(n_121),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_64),
.B2(n_65),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B(n_60),
.Y(n_52)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_56),
.B1(n_68),
.B2(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_54),
.A2(n_72),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_68),
.Y(n_119)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_58),
.A2(n_62),
.B1(n_126),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_58),
.A2(n_62),
.B1(n_147),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_58),
.A2(n_62),
.B1(n_160),
.B2(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B(n_76),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_74),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_66),
.A2(n_106),
.B1(n_108),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_67),
.A2(n_73),
.B1(n_120),
.B2(n_131),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B(n_72),
.C(n_73),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_70),
.Y(n_72)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g120 ( 
.A(n_70),
.B(n_121),
.CON(n_120),
.SN(n_120)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_82),
.A2(n_217),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_88),
.B(n_144),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.C(n_104),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_96),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_99),
.A2(n_104),
.B1(n_105),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_103),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_115),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_110),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_115),
.A2(n_116),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_124),
.C(n_128),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_121),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_128),
.B1(n_129),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_164),
.B(n_251),
.C(n_257),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_152),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_137),
.B(n_152),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_149),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_139),
.B(n_140),
.C(n_149),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.C(n_148),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_153),
.A2(n_154),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_158),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_250),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_243),
.B(n_249),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_195),
.B(n_242),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_185),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_168),
.B(n_185),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_178),
.C(n_181),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_169),
.A2(n_170),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_172),
.Y(n_192)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_186),
.B(n_192),
.C(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_236),
.B(n_241),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_213),
.B(n_235),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_205),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_198),
.B(n_205),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_221),
.B(n_234),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_219),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_233),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);


endmodule