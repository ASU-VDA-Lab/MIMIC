module fake_jpeg_9539_n_78 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_20),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_17),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_10),
.C(n_13),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_20),
.B(n_21),
.C(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_27),
.B1(n_19),
.B2(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_20),
.B(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_37),
.B1(n_32),
.B2(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_15),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_8),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_8),
.C(n_11),
.Y(n_55)
);

XNOR2x1_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_18),
.Y(n_42)
);

XNOR2x1_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_34),
.B1(n_30),
.B2(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_55),
.B(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_40),
.B1(n_46),
.B2(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_42),
.C(n_41),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_43),
.B(n_45),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_54),
.B(n_9),
.Y(n_67)
);

OAI321xp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_50),
.A3(n_21),
.B1(n_18),
.B2(n_19),
.C(n_40),
.Y(n_66)
);

NAND4xp25_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_25),
.C(n_18),
.D(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_53),
.Y(n_65)
);

FAx1_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.CI(n_67),
.CON(n_69),
.SN(n_69)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_58),
.B1(n_9),
.B2(n_55),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_62),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_1),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_0),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_73),
.B(n_2),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.A3(n_71),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_2),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_6),
.Y(n_78)
);


endmodule