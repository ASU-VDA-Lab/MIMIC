module real_jpeg_32657_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

OAI22x1_ASAP7_75t_SL g23 ( 
.A1(n_0),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_0),
.B(n_68),
.Y(n_67)
);

OAI22x1_ASAP7_75t_SL g95 ( 
.A1(n_0),
.A2(n_27),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

AOI22x1_ASAP7_75t_L g178 ( 
.A1(n_0),
.A2(n_27),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_0),
.A2(n_205),
.A3(n_211),
.B1(n_215),
.B2(n_223),
.Y(n_204)
);

NAND2xp67_ASAP7_75t_SL g278 ( 
.A(n_0),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_0),
.B(n_242),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_1),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_2),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_4),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_5),
.A2(n_327),
.B1(n_328),
.B2(n_331),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_5),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_6),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_6),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_6),
.A2(n_318),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_9),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22x1_ASAP7_75t_L g81 ( 
.A1(n_9),
.A2(n_62),
.B1(n_82),
.B2(n_86),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_62),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_62),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_10),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_358),
.Y(n_12)
);

INVxp67_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_299),
.B(n_351),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_233),
.B(n_296),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_188),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_17),
.B(n_188),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_101),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_19),
.B(n_134),
.C(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_66),
.C(n_73),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_20),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_20),
.B(n_307),
.Y(n_343)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_21),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_32),
.B1(n_46),
.B2(n_57),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g338 ( 
.A1(n_22),
.A2(n_46),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22x1_ASAP7_75t_L g185 ( 
.A1(n_23),
.A2(n_33),
.B1(n_47),
.B2(n_58),
.Y(n_185)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_27),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_27),
.A2(n_123),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_27),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_27),
.B(n_34),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_27),
.B(n_264),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g269 ( 
.A1(n_27),
.A2(n_169),
.B(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_48),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_34),
.Y(n_339)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_35),
.B(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_35),
.Y(n_266)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_37),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_37),
.Y(n_201)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_40),
.Y(n_219)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_51),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_65),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_66),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_192)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_68),
.B(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_L g259 ( 
.A(n_73),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_73),
.B(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_74),
.B(n_277),
.Y(n_276)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_80),
.B(n_90),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_79),
.Y(n_279)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_91),
.B1(n_95),
.B2(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_85),
.Y(n_274)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_89),
.Y(n_321)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_89),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_89),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_90),
.A2(n_315),
.B(n_322),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_91),
.Y(n_231)
);

NOR2x1_ASAP7_75t_R g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g232 ( 
.A(n_92),
.Y(n_232)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_95),
.B(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_97),
.Y(n_317)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_101),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_128),
.B1(n_129),
.B2(n_133),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_103),
.B(n_128),
.Y(n_305)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.A3(n_111),
.B1(n_116),
.B2(n_123),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_108),
.A3(n_111),
.B1(n_116),
.B2(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_128),
.B(n_194),
.C(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_128),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_R g282 ( 
.A(n_129),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_129),
.B(n_283),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_158),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_135),
.B(n_385),
.C(n_386),
.Y(n_384)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_137),
.B(n_159),
.C(n_187),
.Y(n_345)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_138),
.B(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_146),
.B(n_147),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_139),
.A2(n_146),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_139),
.A2(n_146),
.B1(n_309),
.B2(n_310),
.Y(n_370)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_148),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_151),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_177),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_169),
.B(n_172),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_168),
.B1(n_178),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_161),
.Y(n_382)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_162),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_163),
.Y(n_281)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_R g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_176),
.Y(n_381)
);

AOI22x1_ASAP7_75t_L g240 ( 
.A1(n_177),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_240)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_178),
.A2(n_376),
.B1(n_382),
.B2(n_383),
.Y(n_375)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_183),
.Y(n_378)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_184),
.A2(n_187),
.B1(n_239),
.B2(n_253),
.Y(n_252)
);

AO22x1_ASAP7_75t_L g368 ( 
.A1(n_184),
.A2(n_185),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.C(n_202),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_193),
.B(n_305),
.C(n_306),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_194),
.A2(n_202),
.B1(n_203),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_194),
.A2(n_195),
.B1(n_255),
.B2(n_290),
.Y(n_289)
);

AO22x1_ASAP7_75t_L g312 ( 
.A1(n_194),
.A2(n_247),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_194),
.B(n_314),
.Y(n_371)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_229),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_229),
.Y(n_244)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_230),
.B(n_326),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_231),
.A2(n_315),
.B1(n_322),
.B2(n_325),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_248),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_236),
.B(n_245),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.C(n_244),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_239),
.A2(n_253),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_239),
.B(n_262),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_239),
.B(n_336),
.Y(n_335)
);

XOR2x2_ASAP7_75t_L g344 ( 
.A(n_239),
.B(n_336),
.Y(n_344)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_243),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_294),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_256),
.B(n_292),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_286),
.B(n_291),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_275),
.B(n_285),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_267),
.B(n_269),
.Y(n_262)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_282),
.B(n_284),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_346),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_301),
.B(n_354),
.Y(n_353)
);

NAND2x1_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_340),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_311),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_311),
.Y(n_356)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_304),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_343),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_334),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_361),
.C(n_363),
.Y(n_360)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx4f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_334),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.C(n_345),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_345),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_349),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_R g358 ( 
.A(n_359),
.B(n_387),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_364),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_360),
.B(n_364),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_384),
.Y(n_364)
);

OAI22x1_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_372),
.B2(n_373),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XOR2x2_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);


endmodule