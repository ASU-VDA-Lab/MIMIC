module fake_jpeg_30283_n_78 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_2),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_45),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_43),
.B1(n_16),
.B2(n_23),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_15),
.B1(n_25),
.B2(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_3),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_55),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_54),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_13),
.B(n_22),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_11),
.C(n_19),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_61),
.C(n_63),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_9),
.C(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_55),
.B1(n_49),
.B2(n_5),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_64),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_7),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.C(n_62),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_26),
.C(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_67),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_72),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_66),
.C(n_60),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_60),
.C(n_71),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_71),
.Y(n_78)
);


endmodule