module fake_netlist_6_359_n_1904 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1904);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1904;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_174),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_21),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_57),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_46),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_93),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_87),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_49),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_11),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_134),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_48),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_38),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_36),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_6),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_50),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_66),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_28),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_136),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_71),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_47),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_83),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_76),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_55),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_63),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_112),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_47),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_104),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_75),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_43),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_42),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_68),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_169),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_148),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_44),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_48),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_143),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_40),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_124),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_113),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_54),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_18),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_0),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_27),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_125),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_173),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_100),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_157),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_65),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_12),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_21),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_1),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_56),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_103),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_16),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_42),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_131),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_118),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_121),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_19),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_144),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_9),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_68),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_161),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_145),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_84),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_90),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_25),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_18),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_82),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_51),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_102),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_5),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_139),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_38),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_132),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_111),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_10),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_162),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_65),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_171),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_80),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_110),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_117),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_176),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_6),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_41),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_109),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_44),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_101),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_57),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_55),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_5),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_52),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_106),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_114),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_98),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_13),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_152),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_14),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_53),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_16),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_66),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_67),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_72),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_15),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_116),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_138),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_33),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_8),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_77),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_107),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_154),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_137),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_140),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_95),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_60),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_24),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_40),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_0),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_91),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_155),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_26),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_168),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_61),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_175),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_35),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_164),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_73),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_158),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_58),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_7),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_96),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_70),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_59),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_22),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_23),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_46),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_156),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_45),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_25),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_167),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_10),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_54),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_51),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_2),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_126),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_32),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_30),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_32),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_26),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_23),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_208),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_254),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_204),
.B(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_208),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_181),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_182),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_208),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_208),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_248),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_184),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_187),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_190),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_204),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_249),
.B(n_1),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_209),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_208),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_300),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_208),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_208),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_208),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_332),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_333),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_193),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_249),
.B(n_2),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_340),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_203),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_205),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_275),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_185),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_209),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_206),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_249),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_270),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_270),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_298),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_215),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_298),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_217),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_218),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_328),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_321),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_192),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_224),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_227),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_228),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_192),
.Y(n_411)
);

INVxp33_ASAP7_75t_SL g412 ( 
.A(n_186),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_189),
.B(n_3),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_235),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_336),
.B(n_3),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_207),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_237),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_232),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_238),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_244),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_245),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_260),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_265),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_269),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_207),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_229),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_229),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_277),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_279),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_280),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_273),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_230),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_230),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_273),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_282),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_328),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_251),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_251),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_284),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_338),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_287),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_338),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_288),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_291),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_252),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_189),
.B(n_4),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_303),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_380),
.B(n_234),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_179),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_257),
.Y(n_454)
);

CKINVDCx8_ASAP7_75t_R g455 ( 
.A(n_361),
.Y(n_455)
);

INVxp33_ASAP7_75t_SL g456 ( 
.A(n_362),
.Y(n_456)
);

NAND2x1_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_328),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_309),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_396),
.B(n_257),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_311),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

AOI22x1_ASAP7_75t_L g463 ( 
.A1(n_371),
.A2(n_307),
.B1(n_355),
.B2(n_354),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_396),
.B(n_179),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_407),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_312),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_387),
.A2(n_198),
.B(n_183),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_359),
.B(n_183),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_416),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_436),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_416),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_357),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_357),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_360),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_427),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_413),
.B(n_315),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_360),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_363),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_363),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_364),
.B(n_198),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_364),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_372),
.B(n_316),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_372),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_437),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_438),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_438),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_374),
.B(n_317),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_L g504 ( 
.A(n_370),
.B(n_328),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_374),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_376),
.B(n_319),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_369),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_376),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_381),
.B(n_320),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_359),
.B(n_274),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_381),
.B(n_326),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_382),
.Y(n_513)
);

INVxp33_ASAP7_75t_SL g514 ( 
.A(n_366),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_393),
.A2(n_324),
.B1(n_226),
.B2(n_256),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_382),
.B(n_330),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_383),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_370),
.B(n_328),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_445),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_383),
.B(n_386),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_388),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_388),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_391),
.B(n_201),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_447),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_494),
.B(n_201),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_447),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_367),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_448),
.B(n_412),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_448),
.B(n_368),
.Y(n_531)
);

OAI21xp33_ASAP7_75t_SL g532 ( 
.A1(n_472),
.A2(n_365),
.B(n_253),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_447),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_481),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_511),
.B(n_379),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_494),
.B(n_210),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_481),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_488),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_451),
.A2(n_252),
.B1(n_255),
.B2(n_253),
.Y(n_540)
);

INVx4_ASAP7_75t_SL g541 ( 
.A(n_520),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_447),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_488),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_518),
.C(n_463),
.Y(n_544)
);

CKINVDCx11_ASAP7_75t_R g545 ( 
.A(n_455),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_451),
.A2(n_255),
.B1(n_276),
.B2(n_261),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_497),
.B(n_385),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_389),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_447),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_494),
.B(n_210),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_520),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_447),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_452),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_495),
.Y(n_555)
);

AOI21x1_ASAP7_75t_L g556 ( 
.A1(n_457),
.A2(n_394),
.B(n_392),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_495),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_L g560 ( 
.A(n_468),
.B(n_400),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_469),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_452),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_488),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_469),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_451),
.B(n_397),
.Y(n_565)
);

BUFx8_ASAP7_75t_SL g566 ( 
.A(n_472),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_521),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_458),
.B(n_403),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_449),
.B(n_390),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_520),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_521),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_452),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_452),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_453),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_511),
.B(n_404),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_515),
.B(n_358),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_478),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_453),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_478),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_L g582 ( 
.A(n_468),
.B(n_408),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_494),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_461),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_461),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_504),
.B(n_394),
.C(n_392),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_461),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_461),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_455),
.B(n_410),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_478),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_482),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_458),
.B(n_414),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_515),
.A2(n_225),
.B1(n_415),
.B2(n_246),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_461),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_494),
.B(n_211),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_454),
.B(n_211),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_464),
.B(n_397),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_482),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_L g600 ( 
.A1(n_449),
.A2(n_415),
.B1(n_296),
.B2(n_295),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_524),
.A2(n_278),
.B1(n_188),
.B2(n_267),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_454),
.A2(n_283),
.B1(n_276),
.B2(n_355),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_503),
.B(n_420),
.Y(n_603)
);

NOR2x1p5_ASAP7_75t_L g604 ( 
.A(n_487),
.B(n_261),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_461),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_461),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_471),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_454),
.B(n_212),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_491),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_467),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_491),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_460),
.B(n_421),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_460),
.B(n_422),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_491),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_471),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_454),
.A2(n_289),
.B1(n_306),
.B2(n_307),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_464),
.B(n_398),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_455),
.B(n_423),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_471),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_488),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_456),
.B(n_424),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_471),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_456),
.B(n_430),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_454),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_520),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_492),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_471),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_492),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_507),
.B(n_435),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_520),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_492),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_477),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_499),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_477),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_472),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_499),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_507),
.B(n_439),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_477),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_517),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_477),
.Y(n_644)
);

AND2x6_ASAP7_75t_L g645 ( 
.A(n_464),
.B(n_212),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_488),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_467),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_510),
.B(n_512),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_450),
.B(n_465),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_510),
.B(n_443),
.Y(n_650)
);

XOR2xp5_ASAP7_75t_L g651 ( 
.A(n_514),
.B(n_373),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_517),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_477),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_508),
.Y(n_655)
);

BUFx4f_ASAP7_75t_L g656 ( 
.A(n_520),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_512),
.B(n_262),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_517),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_516),
.B(n_411),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_463),
.A2(n_294),
.B1(n_258),
.B2(n_318),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_516),
.Y(n_661)
);

BUFx6f_ASAP7_75t_SL g662 ( 
.A(n_459),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_518),
.A2(n_314),
.B1(n_289),
.B2(n_306),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_514),
.B(n_395),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_522),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_520),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_522),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_477),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_477),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_487),
.B(n_334),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_522),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_524),
.B(n_337),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_488),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_523),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_SL g676 ( 
.A(n_459),
.B(n_444),
.Y(n_676)
);

AND3x4_ASAP7_75t_L g677 ( 
.A(n_459),
.B(n_418),
.C(n_378),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_570),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_661),
.B(n_520),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_661),
.B(n_520),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_648),
.B(n_505),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_530),
.A2(n_428),
.B1(n_409),
.B2(n_417),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_627),
.A2(n_656),
.B(n_551),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_531),
.B(n_505),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_568),
.B(n_505),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_567),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_592),
.B(n_505),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_613),
.B(n_505),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_614),
.B(n_627),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_529),
.B(n_513),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_659),
.B(n_429),
.C(n_419),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_611),
.B(n_411),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_547),
.B(n_513),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_537),
.B(n_450),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_649),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_672),
.B(n_441),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_621),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_611),
.B(n_377),
.Y(n_698)
);

AO21x1_ASAP7_75t_L g699 ( 
.A1(n_660),
.A2(n_222),
.B(n_219),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_551),
.B(n_488),
.Y(n_700)
);

BUFx6f_ASAP7_75t_SL g701 ( 
.A(n_657),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_657),
.A2(n_346),
.B1(n_262),
.B2(n_268),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_548),
.B(n_513),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_571),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_609),
.B(n_526),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_593),
.B(n_342),
.C(n_194),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_551),
.B(n_509),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_656),
.B(n_509),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_603),
.B(n_632),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_640),
.B(n_513),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_649),
.Y(n_711)
);

NOR2x1p5_ASAP7_75t_L g712 ( 
.A(n_659),
.B(n_191),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_528),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_650),
.B(n_513),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_571),
.Y(n_715)
);

BUFx8_ASAP7_75t_L g716 ( 
.A(n_574),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_545),
.B(n_195),
.Y(n_717)
);

OAI221xp5_ASAP7_75t_L g718 ( 
.A1(n_532),
.A2(n_180),
.B1(n_264),
.B2(n_348),
.C(n_354),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_583),
.Y(n_719)
);

INVxp33_ASAP7_75t_L g720 ( 
.A(n_654),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_656),
.B(n_509),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_537),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_638),
.B(n_670),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_574),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_638),
.B(n_465),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_528),
.B(n_509),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_534),
.B(n_509),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_534),
.B(n_509),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_570),
.B(n_509),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_552),
.B(n_523),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_552),
.B(n_459),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_570),
.B(n_459),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_555),
.B(n_219),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_579),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_645),
.A2(n_222),
.B1(n_223),
.B2(n_243),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_655),
.B(n_565),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_566),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_621),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_671),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_555),
.B(n_223),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_SL g741 ( 
.A(n_604),
.B(n_243),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_597),
.B(n_473),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_558),
.B(n_247),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_570),
.B(n_266),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_653),
.A2(n_558),
.B(n_570),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_570),
.B(n_247),
.Y(n_746)
);

AOI221xp5_ASAP7_75t_L g747 ( 
.A1(n_601),
.A2(n_283),
.B1(n_310),
.B2(n_314),
.C(n_323),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_565),
.B(n_604),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_595),
.B(n_258),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_624),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_595),
.B(n_285),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_595),
.B(n_285),
.Y(n_752)
);

NAND2x1p5_ASAP7_75t_L g753 ( 
.A(n_628),
.B(n_633),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_597),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_628),
.B(n_633),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_595),
.B(n_286),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_626),
.B(n_196),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_596),
.B(n_286),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_671),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_666),
.B(n_294),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_673),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_596),
.B(n_299),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_673),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_619),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_544),
.A2(n_299),
.B1(n_351),
.B2(n_318),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_666),
.B(n_325),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_601),
.B(n_199),
.C(n_197),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_541),
.B(n_325),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_645),
.A2(n_343),
.B1(n_351),
.B2(n_310),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_596),
.B(n_343),
.Y(n_770)
);

NAND2x1_ASAP7_75t_L g771 ( 
.A(n_583),
.B(n_462),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_541),
.B(n_301),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_596),
.B(n_473),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_619),
.B(n_476),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_645),
.B(n_476),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_541),
.B(n_301),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_583),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_589),
.B(n_479),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_662),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_535),
.B(n_200),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_675),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_620),
.B(n_540),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_583),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_645),
.B(n_479),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_657),
.A2(n_519),
.B1(n_506),
.B2(n_502),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_645),
.B(n_480),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_645),
.B(n_480),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_675),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_645),
.B(n_483),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_578),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_657),
.B(n_483),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_657),
.B(n_484),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_541),
.B(n_301),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_560),
.B(n_484),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_526),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_651),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_578),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_559),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_582),
.B(n_485),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_L g800 ( 
.A(n_609),
.B(n_485),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_544),
.B(n_486),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_600),
.B(n_532),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_576),
.B(n_202),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_525),
.B(n_533),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_559),
.A2(n_457),
.B(n_474),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_561),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_SL g807 ( 
.A(n_546),
.B(n_323),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_561),
.B(n_486),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_569),
.B(n_220),
.C(n_353),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_525),
.B(n_489),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_SL g811 ( 
.A(n_676),
.B(n_216),
.C(n_213),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_609),
.A2(n_348),
.B1(n_506),
.B2(n_502),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_533),
.B(n_489),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_584),
.Y(n_814)
);

NAND2x1p5_ASAP7_75t_L g815 ( 
.A(n_564),
.B(n_457),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_539),
.B(n_490),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_564),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_664),
.B(n_490),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_662),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_539),
.B(n_493),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_549),
.B(n_493),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_581),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_581),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_549),
.B(n_496),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_647),
.B(n_214),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_553),
.B(n_496),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_553),
.B(n_498),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_554),
.B(n_557),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_590),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_609),
.B(n_498),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_591),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_602),
.A2(n_519),
.B(n_501),
.C(n_500),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_591),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_618),
.B(n_500),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_554),
.B(n_501),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_557),
.B(n_462),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_562),
.B(n_466),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_598),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_562),
.B(n_466),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_584),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_572),
.B(n_466),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_598),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_662),
.B(n_527),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_572),
.B(n_470),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_573),
.B(n_470),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_573),
.B(n_470),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_686),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_729),
.A2(n_556),
.B(n_575),
.Y(n_848)
);

AO21x1_ASAP7_75t_L g849 ( 
.A1(n_802),
.A2(n_660),
.B(n_610),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_691),
.B(n_586),
.C(n_231),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_729),
.A2(n_808),
.B(n_680),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_683),
.A2(n_543),
.B(n_538),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_709),
.B(n_609),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_681),
.A2(n_586),
.B(n_580),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_689),
.A2(n_543),
.B(n_538),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_686),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_723),
.A2(n_609),
.B1(n_677),
.B2(n_536),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_757),
.A2(n_663),
.B(n_580),
.C(n_669),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_755),
.A2(n_543),
.B(n_538),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_679),
.A2(n_585),
.B(n_575),
.Y(n_860)
);

INVx6_ASAP7_75t_L g861 ( 
.A(n_716),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_725),
.B(n_609),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_697),
.B(n_585),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_753),
.A2(n_677),
.B1(n_587),
.B2(n_669),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_774),
.B(n_526),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_755),
.A2(n_543),
.B(n_538),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_692),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_737),
.B(n_577),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_697),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_742),
.B(n_526),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_801),
.A2(n_594),
.B(n_587),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_696),
.B(n_677),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_697),
.B(n_738),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_734),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_736),
.B(n_577),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_704),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_697),
.B(n_594),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_738),
.B(n_801),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_738),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_742),
.B(n_526),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_722),
.B(n_526),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_704),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_748),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_715),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_715),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_802),
.A2(n_803),
.B(n_780),
.C(n_782),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_778),
.A2(n_550),
.B1(n_536),
.B2(n_526),
.Y(n_887)
);

INVx11_ASAP7_75t_L g888 ( 
.A(n_716),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_742),
.B(n_536),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_738),
.B(n_795),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_684),
.B(n_536),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_700),
.A2(n_646),
.B(n_563),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_722),
.B(n_695),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_724),
.B(n_651),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_700),
.A2(n_646),
.B(n_563),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_801),
.A2(n_630),
.B(n_605),
.C(n_606),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_747),
.A2(n_599),
.B(n_610),
.C(n_667),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_720),
.B(n_674),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_713),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_685),
.B(n_536),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_687),
.B(n_536),
.Y(n_901)
);

AO21x1_ASAP7_75t_L g902 ( 
.A1(n_741),
.A2(n_612),
.B(n_599),
.Y(n_902)
);

BUFx4f_ASAP7_75t_L g903 ( 
.A(n_779),
.Y(n_903)
);

NOR2xp67_ASAP7_75t_L g904 ( 
.A(n_682),
.B(n_556),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_790),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_745),
.A2(n_805),
.B(n_804),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_818),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_690),
.B(n_605),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_808),
.A2(n_617),
.B(n_608),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_711),
.B(n_232),
.Y(n_910)
);

OAI21xp33_ASAP7_75t_SL g911 ( 
.A1(n_798),
.A2(n_615),
.B(n_612),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_791),
.A2(n_550),
.B1(n_536),
.B2(n_527),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_688),
.B(n_550),
.Y(n_913)
);

INVx11_ASAP7_75t_L g914 ( 
.A(n_716),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_718),
.A2(n_615),
.B(n_629),
.C(n_667),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_693),
.B(n_550),
.Y(n_916)
);

NOR2x1_ASAP7_75t_R g917 ( 
.A(n_794),
.B(n_221),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_767),
.B(n_617),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_797),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_703),
.B(n_622),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_710),
.B(n_622),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_714),
.B(n_550),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_707),
.A2(n_646),
.B(n_563),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_754),
.B(n_764),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_694),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_694),
.B(n_550),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_707),
.A2(n_646),
.B(n_563),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_792),
.A2(n_550),
.B1(n_668),
.B2(n_527),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_708),
.A2(n_584),
.B(n_588),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_L g930 ( 
.A(n_779),
.B(n_584),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_708),
.A2(n_584),
.B(n_588),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_741),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_721),
.A2(n_588),
.B(n_637),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_775),
.A2(n_637),
.B(n_625),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_721),
.A2(n_588),
.B(n_644),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_717),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_784),
.A2(n_787),
.B(n_786),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_779),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_712),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_797),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_789),
.A2(n_773),
.B(n_806),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_678),
.A2(n_588),
.B(n_644),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_779),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_678),
.A2(n_625),
.B(n_668),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_SL g945 ( 
.A1(n_796),
.A2(n_233),
.B1(n_236),
.B2(n_239),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_807),
.A2(n_629),
.B(n_631),
.C(n_665),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_694),
.B(n_631),
.Y(n_947)
);

AO22x1_ASAP7_75t_L g948 ( 
.A1(n_706),
.A2(n_341),
.B1(n_240),
.B2(n_241),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_819),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_678),
.A2(n_668),
.B(n_542),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_834),
.B(n_634),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_814),
.A2(n_542),
.B(n_607),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_719),
.B(n_542),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_814),
.A2(n_607),
.B(n_616),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_719),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_799),
.B(n_634),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_817),
.A2(n_607),
.B1(n_616),
.B2(n_635),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_720),
.B(n_674),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_814),
.A2(n_635),
.B(n_616),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_840),
.A2(n_635),
.B(n_642),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_807),
.A2(n_636),
.B(n_665),
.C(n_658),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_822),
.B(n_636),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_840),
.A2(n_642),
.B(n_674),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_832),
.A2(n_658),
.B(n_652),
.C(n_643),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_783),
.A2(n_642),
.B1(n_623),
.B2(n_643),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_750),
.B(n_639),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_840),
.A2(n_652),
.B(n_641),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_731),
.A2(n_641),
.B(n_639),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_823),
.B(n_623),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_828),
.A2(n_475),
.B(n_474),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_750),
.B(n_623),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_831),
.B(n_475),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_842),
.B(n_475),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_829),
.B(n_474),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_829),
.B(n_242),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_819),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_705),
.A2(n_406),
.B(n_402),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_719),
.B(n_250),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_702),
.A2(n_322),
.B(n_259),
.C(n_263),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_777),
.B(n_272),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_833),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_726),
.A2(n_406),
.B(n_402),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_749),
.A2(n_401),
.B(n_399),
.C(n_398),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_833),
.B(n_838),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_727),
.A2(n_401),
.B(n_399),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_832),
.A2(n_313),
.B(n_352),
.C(n_350),
.Y(n_986)
);

NOR2x1_ASAP7_75t_L g987 ( 
.A(n_777),
.B(n_232),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_728),
.A2(n_281),
.B(n_349),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_730),
.A2(n_290),
.B(n_347),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_800),
.A2(n_292),
.B(n_345),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_777),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_760),
.A2(n_766),
.B(n_785),
.C(n_752),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_810),
.B(n_293),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_813),
.B(n_297),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_819),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_750),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_765),
.A2(n_356),
.B1(n_339),
.B2(n_271),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_771),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_821),
.A2(n_86),
.B(n_172),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_821),
.A2(n_85),
.B(n_170),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_830),
.A2(n_302),
.B(n_335),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_816),
.B(n_304),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_751),
.A2(n_305),
.B(n_331),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_820),
.B(n_308),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_732),
.A2(n_327),
.B(n_329),
.Y(n_1005)
);

AO21x1_ASAP7_75t_L g1006 ( 
.A1(n_756),
.A2(n_758),
.B(n_770),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_760),
.A2(n_356),
.B(n_339),
.C(n_271),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_762),
.A2(n_356),
.B(n_339),
.C(n_271),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_701),
.A2(n_766),
.B1(n_843),
.B2(n_809),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_826),
.B(n_7),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_739),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_819),
.B(n_9),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_824),
.A2(n_165),
.B(n_160),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_835),
.B(n_11),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_732),
.A2(n_153),
.B(n_147),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_739),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_759),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_759),
.B(n_12),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_815),
.A2(n_146),
.B(n_141),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_815),
.A2(n_135),
.B(n_133),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_825),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_698),
.B(n_13),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_836),
.A2(n_130),
.B(n_128),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_841),
.A2(n_127),
.B(n_120),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_761),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_761),
.B(n_14),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_701),
.B(n_119),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_763),
.B(n_19),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_765),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_844),
.A2(n_115),
.B(n_105),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_763),
.Y(n_1031)
);

CKINVDCx10_ASAP7_75t_R g1032 ( 
.A(n_811),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_781),
.B(n_20),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_869),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_867),
.B(n_733),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_874),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_853),
.A2(n_846),
.B(n_776),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_856),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_886),
.A2(n_740),
.B(n_743),
.C(n_827),
.Y(n_1039)
);

INVxp67_ASAP7_75t_SL g1040 ( 
.A(n_878),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_861),
.B(n_795),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_872),
.B(n_772),
.C(n_776),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_907),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1011),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_867),
.B(n_793),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_SL g1046 ( 
.A(n_1022),
.B(n_699),
.C(n_735),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_986),
.A2(n_827),
.B(n_824),
.C(n_772),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_883),
.B(n_765),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_925),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_893),
.B(n_768),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_875),
.B(n_793),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_937),
.A2(n_812),
.B(n_839),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_891),
.A2(n_845),
.B(n_839),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_900),
.A2(n_845),
.B(n_837),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_901),
.A2(n_837),
.B(n_768),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_913),
.A2(n_788),
.B(n_781),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1011),
.Y(n_1057)
);

BUFx12f_ASAP7_75t_L g1058 ( 
.A(n_861),
.Y(n_1058)
);

INVx6_ASAP7_75t_L g1059 ( 
.A(n_943),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_916),
.A2(n_769),
.B(n_746),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_883),
.B(n_746),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_861),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_986),
.A2(n_744),
.B(n_22),
.C(n_24),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1016),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_876),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_943),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1016),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1021),
.B(n_744),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_893),
.Y(n_1069)
);

INVx6_ASAP7_75t_L g1070 ( 
.A(n_943),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1021),
.B(n_20),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_922),
.A2(n_99),
.B(n_97),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_858),
.A2(n_896),
.B(n_871),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_894),
.B(n_27),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_878),
.A2(n_890),
.B1(n_865),
.B2(n_862),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_925),
.B(n_94),
.Y(n_1076)
);

AND3x1_ASAP7_75t_SL g1077 ( 
.A(n_899),
.B(n_28),
.C(n_29),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_890),
.A2(n_89),
.B1(n_88),
.B2(n_81),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_872),
.A2(n_78),
.B1(n_74),
.B2(n_69),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_924),
.B(n_966),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_941),
.A2(n_29),
.B(n_30),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_936),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_919),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_966),
.B(n_31),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_932),
.B(n_31),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_992),
.A2(n_34),
.B(n_35),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_904),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_939),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_855),
.A2(n_37),
.B(n_39),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_943),
.B(n_45),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_951),
.B(n_898),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_956),
.A2(n_50),
.B(n_52),
.Y(n_1092)
);

INVx3_ASAP7_75t_SL g1093 ( 
.A(n_996),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_898),
.B(n_53),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_857),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_946),
.A2(n_62),
.B(n_64),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_869),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_910),
.B(n_62),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_940),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1029),
.A2(n_64),
.B1(n_67),
.B2(n_850),
.Y(n_1100)
);

CKINVDCx11_ASAP7_75t_R g1101 ( 
.A(n_1012),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_884),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_958),
.B(n_917),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_949),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_946),
.A2(n_961),
.B(n_854),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_958),
.B(n_945),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_949),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_888),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_991),
.A2(n_887),
.B1(n_889),
.B2(n_880),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_885),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_991),
.A2(n_870),
.B1(n_926),
.B2(n_947),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_981),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_847),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_SL g1114 ( 
.A1(n_1022),
.A2(n_997),
.B1(n_1012),
.B2(n_1009),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_948),
.B(n_850),
.C(n_1007),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_993),
.B(n_994),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_882),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_852),
.A2(n_921),
.B(n_908),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1025),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_873),
.A2(n_879),
.B1(n_984),
.B2(n_905),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_933),
.A2(n_935),
.B(n_851),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_987),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1002),
.B(n_1004),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1031),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_975),
.B(n_978),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_920),
.A2(n_921),
.B(n_860),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1017),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_SL g1128 ( 
.A(n_1008),
.B(n_979),
.C(n_864),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_1012),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_978),
.B(n_980),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_903),
.B(n_949),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_SL g1132 ( 
.A(n_903),
.B(n_938),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_997),
.B(n_989),
.C(n_1003),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_949),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_873),
.A2(n_879),
.B1(n_912),
.B2(n_928),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_971),
.B(n_1010),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_962),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_995),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_918),
.A2(n_961),
.B(n_980),
.C(n_988),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1005),
.A2(n_1014),
.B(n_964),
.C(n_990),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_SL g1141 ( 
.A(n_1027),
.B(n_1008),
.C(n_1001),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_914),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_881),
.A2(n_1029),
.B1(n_868),
.B2(n_971),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_920),
.A2(n_906),
.B(n_866),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_897),
.A2(n_915),
.B(n_964),
.C(n_1018),
.Y(n_1145)
);

O2A1O1Ixp5_ASAP7_75t_L g1146 ( 
.A1(n_1006),
.A2(n_902),
.B(n_849),
.C(n_957),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_881),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_976),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_897),
.B(n_955),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_863),
.A2(n_877),
.B(n_895),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_955),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_974),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_859),
.A2(n_923),
.B(n_927),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_915),
.B(n_1033),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_976),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_976),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1026),
.A2(n_1028),
.B(n_983),
.C(n_911),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_968),
.B(n_934),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_L g1159 ( 
.A(n_976),
.B(n_969),
.Y(n_1159)
);

AND2x2_ASAP7_75t_SL g1160 ( 
.A(n_938),
.B(n_930),
.Y(n_1160)
);

BUFx4f_ASAP7_75t_L g1161 ( 
.A(n_998),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_934),
.B(n_998),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_965),
.A2(n_892),
.B1(n_953),
.B2(n_929),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_909),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_972),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_931),
.A2(n_967),
.B(n_952),
.Y(n_1166)
);

NAND2x1_ASAP7_75t_L g1167 ( 
.A(n_963),
.B(n_954),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_959),
.A2(n_960),
.B(n_942),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_848),
.A2(n_950),
.B(n_944),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_973),
.A2(n_977),
.B(n_970),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_1032),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1019),
.A2(n_1020),
.B(n_1024),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_982),
.B(n_985),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_999),
.B(n_1000),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1015),
.B(n_1023),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1030),
.A2(n_1013),
.B1(n_886),
.B2(n_689),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_943),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_874),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1011),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_883),
.B(n_709),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_869),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_861),
.B(n_779),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_867),
.B(n_709),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_907),
.B(n_709),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_886),
.A2(n_709),
.B(n_757),
.C(n_530),
.Y(n_1185)
);

NOR2x1_ASAP7_75t_L g1186 ( 
.A(n_938),
.B(n_886),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_853),
.A2(n_937),
.B(n_689),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_SL g1188 ( 
.A1(n_886),
.A2(n_802),
.B(n_986),
.C(n_896),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_874),
.Y(n_1189)
);

BUFx10_ASAP7_75t_L g1190 ( 
.A(n_1103),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1161),
.Y(n_1191)
);

OAI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1133),
.A2(n_1143),
.B1(n_1106),
.B2(n_1085),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1137),
.B(n_1180),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1105),
.A2(n_1146),
.B(n_1073),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1185),
.A2(n_1146),
.B(n_1187),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1187),
.A2(n_1153),
.B(n_1172),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1153),
.A2(n_1172),
.B(n_1175),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1189),
.B(n_1036),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_SL g1200 ( 
.A(n_1131),
.B(n_1114),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1176),
.A2(n_1154),
.B(n_1144),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1056),
.A2(n_1121),
.B(n_1168),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1144),
.A2(n_1158),
.B(n_1188),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1183),
.A2(n_1051),
.B1(n_1100),
.B2(n_1116),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_1071),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1115),
.B(n_1081),
.C(n_1128),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_1036),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1080),
.B(n_1091),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_1049),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1168),
.A2(n_1166),
.B(n_1118),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_L g1211 ( 
.A1(n_1096),
.A2(n_1081),
.B1(n_1087),
.B2(n_1063),
.C(n_1115),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1101),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1167),
.A2(n_1053),
.B(n_1054),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1125),
.A2(n_1130),
.B(n_1123),
.C(n_1045),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1098),
.A2(n_1079),
.B(n_1046),
.Y(n_1215)
);

AO21x2_ASAP7_75t_L g1216 ( 
.A1(n_1126),
.A2(n_1162),
.B(n_1042),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1126),
.A2(n_1145),
.B(n_1052),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1039),
.A2(n_1140),
.B(n_1037),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1035),
.B(n_1184),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1069),
.B(n_1049),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_1178),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1066),
.B(n_1161),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1039),
.A2(n_1037),
.B(n_1170),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1058),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1136),
.A2(n_1052),
.B(n_1157),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1038),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1127),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1119),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1095),
.A2(n_1084),
.B(n_1086),
.C(n_1141),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1139),
.A2(n_1076),
.B(n_1048),
.C(n_1149),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1157),
.A2(n_1163),
.B(n_1145),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1068),
.B(n_1074),
.Y(n_1232)
);

OR2x6_ASAP7_75t_L g1233 ( 
.A(n_1182),
.B(n_1062),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1053),
.A2(n_1054),
.B(n_1055),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1165),
.B(n_1040),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1040),
.B(n_1152),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1043),
.B(n_1050),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1060),
.A2(n_1186),
.B(n_1159),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1124),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1050),
.B(n_1147),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_SL g1241 ( 
.A1(n_1141),
.A2(n_1046),
.B(n_1094),
.C(n_1086),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1093),
.B(n_1082),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1109),
.A2(n_1075),
.B(n_1111),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1147),
.B(n_1061),
.Y(n_1244)
);

OAI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1128),
.A2(n_1092),
.B(n_1042),
.Y(n_1245)
);

BUFx4f_ASAP7_75t_L g1246 ( 
.A(n_1093),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1060),
.A2(n_1174),
.B(n_1164),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1041),
.A2(n_1090),
.B1(n_1110),
.B2(n_1065),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1122),
.B(n_1088),
.Y(n_1249)
);

AOI21xp33_ASAP7_75t_L g1250 ( 
.A1(n_1063),
.A2(n_1047),
.B(n_1135),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1047),
.A2(n_1089),
.B(n_1092),
.C(n_1072),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1164),
.A2(n_1055),
.B(n_1160),
.Y(n_1252)
);

INVxp67_ASAP7_75t_SL g1253 ( 
.A(n_1034),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1129),
.B(n_1102),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_SL g1255 ( 
.A(n_1089),
.B(n_1072),
.C(n_1142),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1120),
.A2(n_1078),
.A3(n_1113),
.B(n_1117),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1044),
.A2(n_1179),
.A3(n_1057),
.B(n_1067),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1041),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1151),
.B(n_1112),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1041),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1173),
.A2(n_1132),
.B(n_1181),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1034),
.A2(n_1181),
.B(n_1097),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1097),
.A2(n_1099),
.B(n_1083),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1064),
.A2(n_1155),
.B(n_1077),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_SL g1265 ( 
.A1(n_1090),
.A2(n_1059),
.B(n_1070),
.C(n_1066),
.Y(n_1265)
);

NOR2xp67_ASAP7_75t_L g1266 ( 
.A(n_1108),
.B(n_1138),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1090),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1182),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1104),
.B(n_1148),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1182),
.B(n_1134),
.C(n_1156),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1104),
.B(n_1148),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1104),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1059),
.A2(n_1070),
.A3(n_1107),
.B(n_1134),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1107),
.A2(n_1134),
.B(n_1148),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1107),
.B(n_1156),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1059),
.A2(n_1070),
.B1(n_1156),
.B2(n_1177),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1177),
.B(n_1171),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1177),
.A2(n_1105),
.B(n_1146),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1171),
.B(n_358),
.Y(n_1279)
);

BUFx8_ASAP7_75t_SL g1280 ( 
.A(n_1058),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1180),
.B(n_1183),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1127),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1180),
.B(n_1183),
.Y(n_1287)
);

CKINVDCx6p67_ASAP7_75t_R g1288 ( 
.A(n_1093),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1180),
.B(n_875),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1127),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1133),
.A2(n_1185),
.B(n_886),
.C(n_1116),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1108),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1104),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1182),
.B(n_1041),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1302)
);

CKINVDCx11_ASAP7_75t_R g1303 ( 
.A(n_1093),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1183),
.B(n_358),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1133),
.A2(n_1185),
.B(n_886),
.C(n_1116),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1104),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1185),
.A2(n_757),
.B(n_886),
.C(n_709),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_1058),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_SL g1315 ( 
.A1(n_1185),
.A2(n_886),
.B(n_1133),
.C(n_802),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1183),
.B(n_358),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1127),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1161),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1127),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1185),
.A2(n_757),
.B(n_886),
.C(n_709),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1133),
.A2(n_1114),
.B1(n_1183),
.B2(n_872),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1185),
.A2(n_886),
.B(n_1096),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1133),
.A2(n_1185),
.B(n_886),
.C(n_1116),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1187),
.A2(n_886),
.B(n_1185),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1127),
.Y(n_1333)
);

AO21x1_ASAP7_75t_L g1334 ( 
.A1(n_1081),
.A2(n_1086),
.B(n_1096),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1176),
.A2(n_1144),
.A3(n_849),
.B(n_902),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1137),
.B(n_1180),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1133),
.A2(n_1185),
.B(n_886),
.C(n_1116),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1108),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1056),
.A2(n_1169),
.B(n_1150),
.Y(n_1340)
);

NAND3xp33_ASAP7_75t_L g1341 ( 
.A(n_1185),
.B(n_1133),
.C(n_757),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1104),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1180),
.B(n_875),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1133),
.A2(n_747),
.B1(n_593),
.B2(n_524),
.C(n_393),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1185),
.A2(n_886),
.B(n_1096),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1180),
.B(n_875),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1133),
.A2(n_1114),
.B1(n_757),
.B2(n_872),
.Y(n_1347)
);

AO32x2_ASAP7_75t_L g1348 ( 
.A1(n_1114),
.A2(n_1087),
.A3(n_1176),
.B1(n_1135),
.B2(n_1120),
.Y(n_1348)
);

INVxp67_ASAP7_75t_SL g1349 ( 
.A(n_1036),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1144),
.A2(n_1105),
.B(n_1073),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1347),
.A2(n_1192),
.B1(n_1344),
.B2(n_1321),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1246),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1208),
.B(n_1214),
.Y(n_1353)
);

INVx6_ASAP7_75t_L g1354 ( 
.A(n_1342),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1301),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1303),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1286),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1235),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1321),
.A2(n_1211),
.B1(n_1206),
.B2(n_1304),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1226),
.Y(n_1360)
);

CKINVDCx6p67_ASAP7_75t_R g1361 ( 
.A(n_1288),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1280),
.Y(n_1362)
);

CKINVDCx6p67_ASAP7_75t_R g1363 ( 
.A(n_1212),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1208),
.B(n_1194),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1206),
.A2(n_1316),
.B1(n_1204),
.B2(n_1245),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1312),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1204),
.A2(n_1245),
.B1(n_1341),
.B2(n_1334),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1292),
.Y(n_1368)
);

INVx11_ASAP7_75t_L g1369 ( 
.A(n_1312),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1195),
.A2(n_1219),
.B1(n_1350),
.B2(n_1341),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1191),
.Y(n_1371)
);

BUFx4_ASAP7_75t_SL g1372 ( 
.A(n_1224),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1283),
.A2(n_1287),
.B1(n_1343),
.B2(n_1289),
.Y(n_1373)
);

BUFx4_ASAP7_75t_R g1374 ( 
.A(n_1190),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1195),
.A2(n_1350),
.B1(n_1205),
.B2(n_1232),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1346),
.A2(n_1215),
.B1(n_1337),
.B2(n_1194),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1267),
.A2(n_1337),
.B1(n_1248),
.B2(n_1258),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1342),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1205),
.A2(n_1248),
.B1(n_1231),
.B2(n_1217),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1318),
.Y(n_1380)
);

CKINVDCx11_ASAP7_75t_R g1381 ( 
.A(n_1190),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1317),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1327),
.A2(n_1345),
.B1(n_1215),
.B2(n_1305),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1319),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1333),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1293),
.A2(n_1330),
.B1(n_1338),
.B2(n_1235),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1200),
.A2(n_1250),
.B1(n_1264),
.B2(n_1255),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1217),
.A2(n_1278),
.B1(n_1196),
.B2(n_1264),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1246),
.A2(n_1199),
.B1(n_1233),
.B2(n_1318),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1222),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1207),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1228),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1342),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1236),
.A2(n_1250),
.B1(n_1270),
.B2(n_1320),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1296),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1339),
.Y(n_1396)
);

BUFx8_ASAP7_75t_SL g1397 ( 
.A(n_1233),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1220),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1239),
.Y(n_1399)
);

INVx8_ASAP7_75t_L g1400 ( 
.A(n_1233),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_SL g1401 ( 
.A(n_1268),
.Y(n_1401)
);

BUFx4_ASAP7_75t_R g1402 ( 
.A(n_1242),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1221),
.A2(n_1349),
.B1(n_1260),
.B2(n_1236),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1257),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1257),
.Y(n_1405)
);

INVxp33_ASAP7_75t_L g1406 ( 
.A(n_1237),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1259),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1240),
.A2(n_1279),
.B1(n_1307),
.B2(n_1294),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1209),
.B(n_1244),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1271),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1244),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1254),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1270),
.A2(n_1311),
.B1(n_1251),
.B2(n_1278),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1272),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1297),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1297),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1256),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_R g1418 ( 
.A1(n_1277),
.A2(n_1275),
.B1(n_1249),
.B2(n_1348),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1229),
.A2(n_1196),
.B1(n_1243),
.B2(n_1223),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_SL g1420 ( 
.A1(n_1281),
.A2(n_1282),
.B(n_1284),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1285),
.A2(n_1328),
.B1(n_1300),
.B2(n_1302),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1261),
.A2(n_1266),
.B1(n_1332),
.B2(n_1331),
.Y(n_1422)
);

BUFx4f_ASAP7_75t_SL g1423 ( 
.A(n_1297),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1306),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1253),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1306),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1306),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1265),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1291),
.A2(n_1313),
.B1(n_1329),
.B2(n_1218),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1216),
.A2(n_1252),
.B1(n_1238),
.B2(n_1225),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1269),
.Y(n_1431)
);

BUFx2_ASAP7_75t_R g1432 ( 
.A(n_1216),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1201),
.A2(n_1247),
.B1(n_1263),
.B2(n_1203),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1348),
.A2(n_1262),
.B1(n_1274),
.B2(n_1197),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1276),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1348),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1198),
.A2(n_1241),
.B1(n_1315),
.B2(n_1230),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1273),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1234),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1213),
.Y(n_1440)
);

INVx4_ASAP7_75t_SL g1441 ( 
.A(n_1290),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1290),
.A2(n_1335),
.B1(n_1314),
.B2(n_1309),
.Y(n_1442)
);

INVxp67_ASAP7_75t_SL g1443 ( 
.A(n_1210),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1202),
.A2(n_1193),
.B1(n_1336),
.B2(n_1324),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1290),
.A2(n_1295),
.B1(n_1335),
.B2(n_1326),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1295),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1295),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1309),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1309),
.Y(n_1449)
);

INVx4_ASAP7_75t_L g1450 ( 
.A(n_1298),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

INVx8_ASAP7_75t_L g1452 ( 
.A(n_1299),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1308),
.A2(n_1310),
.B1(n_1340),
.B2(n_1322),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1323),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1323),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1323),
.A2(n_1325),
.B1(n_1326),
.B2(n_1335),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1325),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1325),
.A2(n_1204),
.B1(n_1287),
.B2(n_1283),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1326),
.B(n_1208),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1204),
.A2(n_511),
.B1(n_1321),
.B2(n_698),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1347),
.A2(n_1133),
.B1(n_1114),
.B2(n_1192),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1204),
.A2(n_1283),
.B1(n_1287),
.B2(n_1194),
.Y(n_1462)
);

OAI21xp33_ASAP7_75t_L g1463 ( 
.A1(n_1344),
.A2(n_757),
.B(n_511),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1304),
.A2(n_1114),
.B1(n_511),
.B2(n_1022),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1226),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1204),
.A2(n_1283),
.B1(n_1287),
.B2(n_1194),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1227),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1204),
.A2(n_511),
.B1(n_1321),
.B2(n_698),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1304),
.A2(n_1114),
.B1(n_511),
.B2(n_1022),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1199),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1204),
.A2(n_1283),
.B1(n_1287),
.B2(n_1194),
.Y(n_1471)
);

BUFx2_ASAP7_75t_SL g1472 ( 
.A(n_1266),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1347),
.A2(n_1133),
.B1(n_1114),
.B2(n_1192),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1304),
.A2(n_872),
.B1(n_1316),
.B2(n_682),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1303),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1226),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1204),
.A2(n_511),
.B1(n_1321),
.B2(n_698),
.Y(n_1477)
);

OAI22x1_ASAP7_75t_L g1478 ( 
.A1(n_1321),
.A2(n_1204),
.B1(n_1206),
.B2(n_1133),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1226),
.Y(n_1479)
);

INVx6_ASAP7_75t_L g1480 ( 
.A(n_1342),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1246),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1227),
.Y(n_1482)
);

INVx6_ASAP7_75t_L g1483 ( 
.A(n_1342),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1204),
.A2(n_1283),
.B1(n_1287),
.B2(n_1194),
.Y(n_1484)
);

INVx6_ASAP7_75t_L g1485 ( 
.A(n_1342),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1304),
.A2(n_872),
.B1(n_1316),
.B2(n_682),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1404),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1364),
.B(n_1373),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1405),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1434),
.A2(n_1419),
.B(n_1437),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1449),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1451),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1454),
.Y(n_1493)
);

NAND2x1_ASAP7_75t_L g1494 ( 
.A(n_1421),
.B(n_1429),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1459),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1459),
.Y(n_1496)
);

INVxp33_ASAP7_75t_L g1497 ( 
.A(n_1470),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1417),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1452),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1444),
.A2(n_1453),
.B(n_1440),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1440),
.A2(n_1433),
.B(n_1439),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1383),
.A2(n_1353),
.B1(n_1386),
.B2(n_1462),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1383),
.A2(n_1419),
.B1(n_1386),
.B2(n_1436),
.Y(n_1503)
);

AND2x4_ASAP7_75t_SL g1504 ( 
.A(n_1409),
.B(n_1387),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1439),
.A2(n_1430),
.B(n_1413),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1360),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1391),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1420),
.A2(n_1367),
.B(n_1448),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1436),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1441),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1452),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1464),
.A2(n_1469),
.B1(n_1477),
.B2(n_1460),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1443),
.A2(n_1445),
.B(n_1442),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1413),
.A2(n_1443),
.B(n_1456),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1364),
.B(n_1462),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1474),
.B(n_1486),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1455),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1358),
.Y(n_1518)
);

AND2x4_ASAP7_75t_SL g1519 ( 
.A(n_1438),
.B(n_1390),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1442),
.A2(n_1445),
.B(n_1456),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1464),
.A2(n_1469),
.B1(n_1359),
.B2(n_1463),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1370),
.B(n_1478),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1358),
.Y(n_1523)
);

AO21x1_ASAP7_75t_L g1524 ( 
.A1(n_1468),
.A2(n_1394),
.B(n_1376),
.Y(n_1524)
);

CKINVDCx6p67_ASAP7_75t_R g1525 ( 
.A(n_1395),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1351),
.A2(n_1365),
.B1(n_1461),
.B2(n_1473),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1446),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1457),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1403),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1370),
.B(n_1375),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1466),
.B(n_1471),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1400),
.B(n_1394),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1465),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_R g1534 ( 
.A(n_1356),
.B(n_1354),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1396),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1422),
.A2(n_1458),
.B(n_1353),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1355),
.B(n_1411),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1398),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1466),
.A2(n_1484),
.B1(n_1471),
.B2(n_1418),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1431),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1476),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1377),
.B(n_1450),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1479),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1450),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1388),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1400),
.B(n_1458),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1388),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1375),
.B(n_1379),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1447),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1354),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1432),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1432),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1392),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1399),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1379),
.B(n_1408),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1425),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1382),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1384),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1385),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1484),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1397),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1357),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1407),
.B(n_1389),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1368),
.B(n_1482),
.Y(n_1564)
);

BUFx10_ASAP7_75t_L g1565 ( 
.A(n_1401),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1467),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1410),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1412),
.B(n_1406),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1371),
.A2(n_1380),
.B(n_1416),
.Y(n_1569)
);

NOR2x1_ASAP7_75t_R g1570 ( 
.A(n_1362),
.B(n_1381),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1435),
.B(n_1472),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1378),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1378),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1485),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1485),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1393),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1393),
.Y(n_1577)
);

AO21x1_ASAP7_75t_SL g1578 ( 
.A1(n_1428),
.A2(n_1374),
.B(n_1480),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1483),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1527),
.B(n_1352),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1515),
.B(n_1481),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1527),
.B(n_1528),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1506),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1518),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1488),
.B(n_1415),
.Y(n_1585)
);

INVx5_ASAP7_75t_L g1586 ( 
.A(n_1532),
.Y(n_1586)
);

AND2x2_ASAP7_75t_SL g1587 ( 
.A(n_1519),
.B(n_1402),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1568),
.B(n_1426),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1568),
.B(n_1424),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1516),
.A2(n_1401),
.B1(n_1366),
.B2(n_1475),
.C(n_1372),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1526),
.A2(n_1361),
.B(n_1363),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1414),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1570),
.B(n_1423),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1552),
.B(n_1414),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1512),
.A2(n_1369),
.B1(n_1414),
.B2(n_1427),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1565),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1525),
.Y(n_1598)
);

O2A1O1Ixp5_ASAP7_75t_L g1599 ( 
.A1(n_1524),
.A2(n_1531),
.B(n_1494),
.C(n_1522),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1512),
.A2(n_1521),
.B(n_1539),
.Y(n_1600)
);

BUFx4f_ASAP7_75t_SL g1601 ( 
.A(n_1525),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1570),
.B(n_1561),
.Y(n_1602)
);

OR2x6_ASAP7_75t_L g1603 ( 
.A(n_1546),
.B(n_1532),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_SL g1604 ( 
.A1(n_1549),
.A2(n_1494),
.B(n_1571),
.C(n_1563),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1503),
.A2(n_1555),
.B(n_1548),
.C(n_1560),
.Y(n_1605)
);

BUFx5_ASAP7_75t_L g1606 ( 
.A(n_1498),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1555),
.A2(n_1548),
.B(n_1560),
.C(n_1504),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1565),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1502),
.A2(n_1529),
.B(n_1505),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1524),
.A2(n_1502),
.B1(n_1532),
.B2(n_1546),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1565),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1530),
.A2(n_1490),
.B(n_1520),
.C(n_1545),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1545),
.A2(n_1547),
.B1(n_1530),
.B2(n_1536),
.C(n_1538),
.Y(n_1614)
);

AO21x2_ASAP7_75t_L g1615 ( 
.A1(n_1500),
.A2(n_1505),
.B(n_1514),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1564),
.B(n_1537),
.Y(n_1616)
);

BUFx4f_ASAP7_75t_SL g1617 ( 
.A(n_1561),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1497),
.B(n_1556),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1564),
.B(n_1554),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1514),
.A2(n_1520),
.B(n_1547),
.Y(n_1620)
);

O2A1O1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1567),
.A2(n_1490),
.B(n_1536),
.C(n_1546),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1490),
.A2(n_1523),
.B(n_1536),
.C(n_1496),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1554),
.B(n_1557),
.Y(n_1623)
);

AO32x2_ASAP7_75t_L g1624 ( 
.A1(n_1550),
.A2(n_1573),
.A3(n_1496),
.B1(n_1495),
.B2(n_1509),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1557),
.B(n_1553),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1495),
.A2(n_1541),
.B(n_1543),
.C(n_1533),
.Y(n_1626)
);

INVx5_ASAP7_75t_L g1627 ( 
.A(n_1544),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1501),
.A2(n_1569),
.B(n_1500),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1542),
.B(n_1499),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1584),
.B(n_1508),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1629),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1598),
.Y(n_1632)
);

NOR2xp67_ASAP7_75t_L g1633 ( 
.A(n_1586),
.B(n_1499),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1620),
.B(n_1513),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1613),
.B(n_1517),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1583),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1613),
.B(n_1513),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1629),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1600),
.A2(n_1508),
.B1(n_1574),
.B2(n_1575),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1609),
.B(n_1513),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1620),
.B(n_1491),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1624),
.B(n_1493),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1599),
.A2(n_1558),
.B1(n_1559),
.B2(n_1566),
.C(n_1562),
.Y(n_1644)
);

NAND2x1_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1511),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1586),
.B(n_1510),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1624),
.B(n_1492),
.Y(n_1647)
);

NAND2x1p5_ASAP7_75t_L g1648 ( 
.A(n_1627),
.B(n_1501),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1624),
.B(n_1492),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1622),
.B(n_1544),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1624),
.B(n_1493),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1487),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1625),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1623),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1628),
.B(n_1489),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1543),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1581),
.B(n_1565),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1619),
.B(n_1626),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1634),
.B(n_1622),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1643),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1642),
.Y(n_1661)
);

AOI33xp33_ASAP7_75t_L g1662 ( 
.A1(n_1640),
.A2(n_1621),
.A3(n_1604),
.B1(n_1611),
.B2(n_1591),
.B3(n_1618),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_R g1663 ( 
.A(n_1632),
.B(n_1598),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1634),
.B(n_1603),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1645),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1643),
.B(n_1626),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1644),
.A2(n_1599),
.B1(n_1605),
.B2(n_1610),
.C(n_1604),
.Y(n_1667)
);

NAND4xp25_ASAP7_75t_SL g1668 ( 
.A(n_1644),
.B(n_1605),
.C(n_1607),
.D(n_1590),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1634),
.Y(n_1669)
);

AO21x2_ASAP7_75t_L g1670 ( 
.A1(n_1638),
.A2(n_1607),
.B(n_1498),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1582),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1643),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1647),
.B(n_1603),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1646),
.Y(n_1674)
);

NAND2x1p5_ASAP7_75t_L g1675 ( 
.A(n_1650),
.B(n_1627),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1630),
.B(n_1616),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_SL g1677 ( 
.A(n_1657),
.B(n_1535),
.C(n_1592),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1645),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1656),
.A2(n_1596),
.B1(n_1587),
.B2(n_1601),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1656),
.B(n_1587),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1649),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1649),
.B(n_1651),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1651),
.B(n_1606),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1651),
.Y(n_1684)
);

INVx5_ASAP7_75t_SL g1685 ( 
.A(n_1646),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1652),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1648),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1636),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1666),
.B(n_1671),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1635),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1671),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1674),
.B(n_1633),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1661),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1682),
.B(n_1641),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1660),
.B(n_1635),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1666),
.B(n_1658),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1650),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1671),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1675),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1666),
.B(n_1671),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1688),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1682),
.B(n_1641),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1655),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1633),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1688),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1676),
.B(n_1658),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1655),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1672),
.B(n_1655),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1676),
.B(n_1653),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1681),
.B(n_1684),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1665),
.B(n_1637),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1681),
.B(n_1631),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1661),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1682),
.B(n_1681),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1676),
.B(n_1653),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1688),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1683),
.B(n_1639),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1683),
.B(n_1639),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1686),
.Y(n_1719)
);

INVx2_ASAP7_75t_SL g1720 ( 
.A(n_1675),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1661),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1676),
.B(n_1654),
.Y(n_1722)
);

NAND2x1_ASAP7_75t_L g1723 ( 
.A(n_1711),
.B(n_1674),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1710),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1696),
.B(n_1662),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1701),
.Y(n_1726)
);

OAI21xp33_ASAP7_75t_L g1727 ( 
.A1(n_1696),
.A2(n_1662),
.B(n_1668),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1701),
.Y(n_1728)
);

NAND2x1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.B(n_1674),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1701),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1706),
.B(n_1680),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1717),
.B(n_1718),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1717),
.B(n_1674),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1717),
.B(n_1674),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1689),
.B(n_1686),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1710),
.Y(n_1736)
);

AND2x2_ASAP7_75t_SL g1737 ( 
.A(n_1692),
.B(n_1667),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1691),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1710),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1718),
.B(n_1674),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1718),
.B(n_1685),
.Y(n_1741)
);

INVx4_ASAP7_75t_L g1742 ( 
.A(n_1692),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1689),
.B(n_1686),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1706),
.B(n_1680),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1700),
.B(n_1667),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1716),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1700),
.A2(n_1668),
.B1(n_1667),
.B2(n_1670),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1716),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1716),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1699),
.B(n_1665),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1709),
.B(n_1659),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1705),
.Y(n_1752)
);

AND2x4_ASAP7_75t_SL g1753 ( 
.A(n_1692),
.B(n_1677),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1709),
.B(n_1659),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1705),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1715),
.B(n_1659),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1691),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1690),
.B(n_1685),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1692),
.B(n_1668),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1722),
.B(n_1602),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1692),
.B(n_1665),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1698),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1715),
.B(n_1659),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1698),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1694),
.B(n_1686),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1738),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1732),
.B(n_1704),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1751),
.B(n_1694),
.Y(n_1768)
);

OAI31xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1759),
.A2(n_1727),
.A3(n_1760),
.B(n_1741),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1725),
.B(n_1722),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1732),
.B(n_1704),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1723),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1745),
.B(n_1617),
.Y(n_1773)
);

NAND2xp33_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1663),
.Y(n_1774)
);

NOR2x1_ASAP7_75t_L g1775 ( 
.A(n_1723),
.B(n_1665),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1729),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1737),
.B(n_1679),
.C(n_1677),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1762),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1754),
.B(n_1694),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1737),
.B(n_1704),
.Y(n_1780)
);

NOR2x1p5_ASAP7_75t_L g1781 ( 
.A(n_1731),
.B(n_1665),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1724),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1753),
.B(n_1704),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1744),
.B(n_1690),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1756),
.B(n_1702),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1763),
.B(n_1690),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1757),
.B(n_1702),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1752),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1753),
.B(n_1741),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1757),
.B(n_1764),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1764),
.B(n_1695),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1758),
.A2(n_1679),
.B(n_1675),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1758),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1742),
.B(n_1704),
.Y(n_1794)
);

NAND2x1_ASAP7_75t_L g1795 ( 
.A(n_1742),
.B(n_1697),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1761),
.A2(n_1670),
.B1(n_1677),
.B2(n_1664),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1742),
.B(n_1697),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1761),
.B(n_1617),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1724),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1735),
.B(n_1702),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1761),
.B(n_1697),
.Y(n_1801)
);

OAI21xp33_ASAP7_75t_L g1802 ( 
.A1(n_1769),
.A2(n_1743),
.B(n_1735),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1790),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1777),
.A2(n_1675),
.B1(n_1729),
.B2(n_1685),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1770),
.B(n_1695),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1766),
.B(n_1695),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1774),
.A2(n_1675),
.B(n_1750),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1797),
.Y(n_1808)
);

AOI32xp33_ASAP7_75t_L g1809 ( 
.A1(n_1774),
.A2(n_1740),
.A3(n_1733),
.B1(n_1734),
.B2(n_1699),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1790),
.Y(n_1810)
);

OAI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1792),
.A2(n_1675),
.B(n_1750),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1796),
.A2(n_1685),
.B1(n_1750),
.B2(n_1678),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1780),
.B(n_1733),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1778),
.B(n_1734),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1780),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1788),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_SL g1817 ( 
.A1(n_1789),
.A2(n_1670),
.B1(n_1663),
.B2(n_1740),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1799),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1787),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1773),
.B(n_1793),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1784),
.B(n_1712),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1797),
.Y(n_1822)
);

OAI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1795),
.A2(n_1699),
.B1(n_1720),
.B2(n_1678),
.C(n_1743),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1787),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1791),
.Y(n_1825)
);

AOI322xp5_ASAP7_75t_L g1826 ( 
.A1(n_1786),
.A2(n_1669),
.A3(n_1708),
.B1(n_1707),
.B2(n_1703),
.C1(n_1686),
.C2(n_1673),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1782),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1815),
.A2(n_1781),
.B1(n_1775),
.B2(n_1798),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1818),
.B(n_1801),
.Y(n_1829)
);

AOI211xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1804),
.A2(n_1789),
.B(n_1783),
.C(n_1794),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1803),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1803),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1813),
.Y(n_1833)
);

AOI32xp33_ASAP7_75t_L g1834 ( 
.A1(n_1817),
.A2(n_1783),
.A3(n_1801),
.B1(n_1794),
.B2(n_1771),
.Y(n_1834)
);

NOR4xp25_ASAP7_75t_SL g1835 ( 
.A(n_1819),
.B(n_1824),
.C(n_1810),
.D(n_1802),
.Y(n_1835)
);

INVxp67_ASAP7_75t_SL g1836 ( 
.A(n_1819),
.Y(n_1836)
);

AOI222xp33_ASAP7_75t_L g1837 ( 
.A1(n_1807),
.A2(n_1767),
.B1(n_1771),
.B2(n_1772),
.C1(n_1776),
.C2(n_1782),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1813),
.Y(n_1838)
);

NAND2x1_ASAP7_75t_L g1839 ( 
.A(n_1824),
.B(n_1772),
.Y(n_1839)
);

NAND3xp33_ASAP7_75t_L g1840 ( 
.A(n_1809),
.B(n_1795),
.C(n_1776),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1808),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1820),
.A2(n_1534),
.B(n_1720),
.Y(n_1842)
);

OAI21xp33_ASAP7_75t_L g1843 ( 
.A1(n_1814),
.A2(n_1779),
.B(n_1768),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1825),
.B(n_1601),
.Y(n_1844)
);

OAI221xp5_ASAP7_75t_SL g1845 ( 
.A1(n_1826),
.A2(n_1785),
.B1(n_1779),
.B2(n_1768),
.C(n_1800),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1808),
.A2(n_1767),
.B1(n_1670),
.B2(n_1720),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1822),
.B(n_1785),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1833),
.A2(n_1822),
.B1(n_1806),
.B2(n_1811),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1836),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1832),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1845),
.A2(n_1812),
.B1(n_1816),
.B2(n_1823),
.C(n_1827),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1841),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1841),
.Y(n_1853)
);

NAND2xp33_ASAP7_75t_L g1854 ( 
.A(n_1834),
.B(n_1805),
.Y(n_1854)
);

NAND3xp33_ASAP7_75t_L g1855 ( 
.A(n_1835),
.B(n_1821),
.C(n_1594),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1844),
.B(n_1800),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1847),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1837),
.A2(n_1728),
.B(n_1726),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1838),
.B(n_1765),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1839),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1855),
.A2(n_1840),
.B(n_1830),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1852),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1857),
.B(n_1829),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1855),
.A2(n_1828),
.B(n_1842),
.Y(n_1864)
);

NOR3xp33_ASAP7_75t_L g1865 ( 
.A(n_1856),
.B(n_1831),
.C(n_1843),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1860),
.B(n_1835),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_SL g1867 ( 
.A(n_1849),
.B(n_1846),
.C(n_1589),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1848),
.B(n_1678),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1851),
.B(n_1728),
.C(n_1726),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1853),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1850),
.B(n_1736),
.Y(n_1871)
);

NAND4xp75_ASAP7_75t_L g1872 ( 
.A(n_1858),
.B(n_1746),
.C(n_1748),
.D(n_1730),
.Y(n_1872)
);

AOI222xp33_ASAP7_75t_L g1873 ( 
.A1(n_1861),
.A2(n_1854),
.B1(n_1859),
.B2(n_1669),
.C1(n_1687),
.C2(n_1749),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1869),
.A2(n_1678),
.B1(n_1714),
.B2(n_1685),
.Y(n_1874)
);

A2O1A1Ixp33_ASAP7_75t_L g1875 ( 
.A1(n_1866),
.A2(n_1678),
.B(n_1687),
.C(n_1765),
.Y(n_1875)
);

OAI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1864),
.A2(n_1687),
.B(n_1612),
.C(n_1608),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1865),
.A2(n_1749),
.B1(n_1748),
.B2(n_1746),
.C(n_1730),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1873),
.B(n_1862),
.Y(n_1878)
);

NOR3xp33_ASAP7_75t_L g1879 ( 
.A(n_1876),
.B(n_1863),
.C(n_1870),
.Y(n_1879)
);

O2A1O1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1875),
.A2(n_1868),
.B(n_1867),
.C(n_1871),
.Y(n_1880)
);

OAI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1874),
.A2(n_1867),
.B1(n_1872),
.B2(n_1597),
.C(n_1608),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1877),
.B(n_1755),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1874),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1883),
.Y(n_1884)
);

A2O1A1Ixp33_ASAP7_75t_L g1885 ( 
.A1(n_1880),
.A2(n_1752),
.B(n_1739),
.C(n_1736),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1878),
.B(n_1739),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1882),
.Y(n_1887)
);

NAND4xp75_ASAP7_75t_L g1888 ( 
.A(n_1879),
.B(n_1593),
.C(n_1595),
.D(n_1588),
.Y(n_1888)
);

NAND3xp33_ASAP7_75t_L g1889 ( 
.A(n_1884),
.B(n_1881),
.C(n_1612),
.Y(n_1889)
);

AOI211xp5_ASAP7_75t_L g1890 ( 
.A1(n_1886),
.A2(n_1580),
.B(n_1687),
.C(n_1719),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1888),
.B(n_1712),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1891),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1892),
.A2(n_1889),
.B1(n_1887),
.B2(n_1885),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1893),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1893),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1894),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_1895),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1890),
.B1(n_1714),
.B2(n_1693),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1896),
.A2(n_1714),
.B1(n_1693),
.B2(n_1713),
.Y(n_1899)
);

OAI21xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1898),
.A2(n_1578),
.B(n_1572),
.Y(n_1900)
);

AND3x1_ASAP7_75t_L g1901 ( 
.A(n_1900),
.B(n_1899),
.C(n_1572),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1901),
.Y(n_1902)
);

OAI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1585),
.B1(n_1719),
.B2(n_1721),
.C(n_1693),
.Y(n_1903)
);

AOI211xp5_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1577),
.B(n_1576),
.C(n_1579),
.Y(n_1904)
);


endmodule