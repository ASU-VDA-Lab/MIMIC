module fake_jpeg_2442_n_591 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_591);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_591;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_55),
.B(n_59),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_68),
.Y(n_113)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_72),
.Y(n_117)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_23),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_54),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_24),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_102),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_34),
.B(n_0),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_2),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_35),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_26),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_92),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_97),
.Y(n_132)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_1),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_1),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_53),
.B(n_51),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_24),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_55),
.B(n_27),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_139),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_59),
.A2(n_50),
.B1(n_22),
.B2(n_29),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_123),
.A2(n_143),
.B1(n_152),
.B2(n_174),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_27),
.B1(n_52),
.B2(n_44),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_126),
.A2(n_141),
.B1(n_156),
.B2(n_88),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_85),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_65),
.A2(n_28),
.B1(n_36),
.B2(n_48),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_138),
.A2(n_37),
.B1(n_32),
.B2(n_57),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_53),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_66),
.A2(n_22),
.B1(n_29),
.B2(n_28),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_75),
.A2(n_50),
.B1(n_29),
.B2(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_42),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_44),
.B1(n_52),
.B2(n_39),
.Y(n_147)
);

AOI22x1_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_149),
.B1(n_61),
.B2(n_85),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_93),
.A2(n_39),
.B1(n_48),
.B2(n_28),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_75),
.A2(n_50),
.B1(n_29),
.B2(n_36),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_58),
.A2(n_53),
.B1(n_51),
.B2(n_49),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_51),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_159),
.B(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_97),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_67),
.B(n_49),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_80),
.A2(n_49),
.B1(n_37),
.B2(n_32),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_80),
.A2(n_37),
.B1(n_32),
.B2(n_47),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_175),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_232)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_178),
.A2(n_183),
.B1(n_204),
.B2(n_218),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_179),
.B(n_219),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_R g272 ( 
.A(n_180),
.B(n_190),
.Y(n_272)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_96),
.B1(n_81),
.B2(n_62),
.Y(n_183)
);

INVx6_ASAP7_75t_SL g184 ( 
.A(n_163),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_184),
.Y(n_289)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_139),
.A2(n_89),
.B1(n_64),
.B2(n_77),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_186),
.A2(n_202),
.B1(n_217),
.B2(n_124),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_76),
.B(n_85),
.C(n_61),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_187),
.B(n_203),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_117),
.B(n_121),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_189),
.B(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_73),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_136),
.B(n_94),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_193),
.B(n_196),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_97),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_194),
.B(n_195),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_122),
.B(n_47),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_113),
.B(n_100),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_197),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_198),
.A2(n_234),
.B1(n_150),
.B2(n_169),
.Y(n_245)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_142),
.B(n_99),
.Y(n_201)
);

NAND2xp67_ASAP7_75t_L g266 ( 
.A(n_201),
.B(n_10),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_120),
.A2(n_91),
.B1(n_79),
.B2(n_78),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_163),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_141),
.A2(n_101),
.B1(n_95),
.B2(n_74),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_132),
.B(n_83),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_206),
.B(n_225),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_142),
.B(n_63),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_207),
.B(n_215),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_110),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_155),
.B(n_171),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_235),
.Y(n_267)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_114),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_110),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_120),
.A2(n_104),
.B1(n_103),
.B2(n_86),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_120),
.A2(n_92),
.B1(n_87),
.B2(n_70),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_137),
.B(n_86),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_161),
.B(n_4),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_154),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_233),
.Y(n_288)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g241 ( 
.A(n_227),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

AO22x1_ASAP7_75t_L g229 ( 
.A1(n_125),
.A2(n_82),
.B1(n_69),
.B2(n_98),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_230),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_125),
.B(n_98),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_167),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_232),
.A2(n_154),
.B1(n_169),
.B2(n_129),
.Y(n_252)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_112),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_118),
.A2(n_5),
.B(n_7),
.C(n_10),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_168),
.B(n_10),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_238),
.Y(n_274)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_118),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_237),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_129),
.B(n_10),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_240),
.B(n_243),
.Y(n_302)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_127),
.B1(n_140),
.B2(n_144),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_266),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_190),
.B(n_140),
.C(n_153),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_260),
.C(n_277),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_252),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_179),
.A2(n_111),
.B1(n_170),
.B2(n_116),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_255),
.A2(n_263),
.B1(n_265),
.B2(n_269),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_203),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_224),
.A2(n_173),
.B1(n_167),
.B2(n_153),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_259),
.A2(n_184),
.B1(n_230),
.B2(n_201),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_195),
.B(n_131),
.C(n_145),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_204),
.A2(n_170),
.B1(n_116),
.B2(n_115),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_186),
.A2(n_150),
.B1(n_158),
.B2(n_145),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_271),
.B1(n_286),
.B2(n_178),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_208),
.A2(n_158),
.B1(n_11),
.B2(n_12),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_178),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_183),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_194),
.A2(n_19),
.B1(n_12),
.B2(n_13),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_275),
.A2(n_216),
.B1(n_199),
.B2(n_222),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_206),
.B(n_191),
.C(n_181),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_11),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_285),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_14),
.C(n_15),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_283),
.B(n_279),
.C(n_291),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_180),
.B(n_15),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_202),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_187),
.B(n_229),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_295),
.A2(n_328),
.B(n_343),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_297),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_238),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_310),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_289),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_304),
.Y(n_386)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_288),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_305),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_247),
.A2(n_224),
.B1(n_180),
.B2(n_218),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_247),
.A2(n_267),
.B1(n_240),
.B2(n_268),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_247),
.A2(n_236),
.B1(n_182),
.B2(n_176),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_176),
.Y(n_310)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_262),
.A2(n_217),
.B1(n_235),
.B2(n_229),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_312),
.A2(n_321),
.B1(n_329),
.B2(n_336),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_313),
.A2(n_318),
.B(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_201),
.B(n_230),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_315),
.A2(n_341),
.B(n_278),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_182),
.B1(n_197),
.B2(n_210),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_320),
.B1(n_323),
.B2(n_327),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_317),
.B(n_339),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_257),
.A2(n_219),
.B(n_209),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_254),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_322),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_257),
.A2(n_197),
.B1(n_219),
.B2(n_216),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_255),
.A2(n_209),
.B1(n_221),
.B2(n_223),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_244),
.B(n_273),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_245),
.A2(n_292),
.B1(n_264),
.B2(n_274),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_242),
.Y(n_324)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_324),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_237),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_326),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_244),
.B(n_226),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_272),
.A2(n_233),
.B1(n_221),
.B2(n_227),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_291),
.A2(n_231),
.B(n_211),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_263),
.A2(n_185),
.B1(n_205),
.B2(n_177),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_228),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_242),
.B(n_220),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_200),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_272),
.B(n_213),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_340),
.C(n_293),
.Y(n_349)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_250),
.Y(n_335)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_248),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_265),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_251),
.B(n_19),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_256),
.A2(n_260),
.B(n_246),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_287),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_342),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_251),
.B(n_287),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_246),
.A2(n_282),
.B(n_285),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_266),
.B(n_293),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_275),
.B(n_283),
.Y(n_345)
);

NOR4xp25_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_294),
.C(n_241),
.D(n_249),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_312),
.A2(n_302),
.B1(n_300),
.B2(n_298),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_347),
.A2(n_369),
.B1(n_371),
.B2(n_373),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_349),
.B(n_381),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_378),
.Y(n_404)
);

OAI32xp33_ASAP7_75t_L g359 ( 
.A1(n_308),
.A2(n_282),
.A3(n_243),
.B1(n_294),
.B2(n_253),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_365),
.Y(n_395)
);

A2O1A1O1Ixp25_ASAP7_75t_L g426 ( 
.A1(n_360),
.A2(n_364),
.B(n_354),
.C(n_372),
.D(n_389),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_297),
.A2(n_271),
.B1(n_286),
.B2(n_243),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_362),
.A2(n_372),
.B1(n_379),
.B2(n_382),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_341),
.A2(n_276),
.B(n_280),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_364),
.A2(n_366),
.B(n_367),
.Y(n_410)
);

AO22x1_ASAP7_75t_SL g365 ( 
.A1(n_302),
.A2(n_243),
.B1(n_249),
.B2(n_253),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_307),
.A2(n_302),
.B1(n_323),
.B2(n_334),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_312),
.A2(n_302),
.B1(n_300),
.B2(n_307),
.Y(n_369)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_342),
.Y(n_370)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_299),
.A2(n_290),
.B1(n_270),
.B2(n_278),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_306),
.A2(n_261),
.B1(n_270),
.B2(n_307),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_299),
.A2(n_261),
.B1(n_325),
.B2(n_295),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_261),
.C(n_330),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_318),
.C(n_328),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_295),
.A2(n_261),
.B(n_307),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_309),
.A2(n_304),
.B1(n_344),
.B2(n_320),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_344),
.A2(n_328),
.B1(n_340),
.B2(n_321),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_381),
.A2(n_369),
.B1(n_373),
.B2(n_347),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_345),
.A2(n_327),
.B1(n_340),
.B2(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_303),
.Y(n_387)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_313),
.A2(n_315),
.B(n_305),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_389),
.A2(n_366),
.B(n_346),
.Y(n_422)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_333),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_405),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_386),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_393),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_386),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_301),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g456 ( 
.A(n_396),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_310),
.Y(n_397)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_378),
.Y(n_398)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_398),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_375),
.B(n_348),
.Y(n_401)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_401),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_322),
.Y(n_402)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_339),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_412),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_333),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_407),
.A2(n_406),
.B1(n_415),
.B2(n_424),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_417),
.C(n_428),
.Y(n_446)
);

OAI22x1_ASAP7_75t_L g411 ( 
.A1(n_367),
.A2(n_313),
.B1(n_332),
.B2(n_336),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_411),
.A2(n_363),
.B1(n_360),
.B2(n_378),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_374),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_358),
.B(n_343),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_418),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_356),
.A2(n_324),
.B1(n_335),
.B2(n_338),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_415),
.A2(n_420),
.B1(n_350),
.B2(n_390),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_353),
.A2(n_337),
.B1(n_317),
.B2(n_329),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_416),
.A2(n_421),
.B1(n_365),
.B2(n_368),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_348),
.B(n_296),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_358),
.B(n_296),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_382),
.B(n_379),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_419),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_356),
.A2(n_316),
.B1(n_319),
.B2(n_311),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_353),
.A2(n_311),
.B1(n_362),
.B2(n_361),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_422),
.A2(n_426),
.B(n_423),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_384),
.B(n_355),
.Y(n_423)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_355),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_424),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_370),
.Y(n_425)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_425),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_370),
.B(n_371),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_427),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_350),
.B(n_368),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_429),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_378),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_448),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_433),
.A2(n_443),
.B1(n_458),
.B2(n_421),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_434),
.B(n_438),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_398),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_441),
.A2(n_442),
.B1(n_447),
.B2(n_395),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_407),
.A2(n_361),
.B1(n_363),
.B2(n_359),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_380),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_380),
.C(n_383),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_451),
.C(n_453),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_383),
.C(n_385),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_385),
.C(n_387),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_365),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_414),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_406),
.B(n_365),
.C(n_352),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_461),
.C(n_409),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_395),
.A2(n_352),
.B1(n_420),
.B2(n_394),
.Y(n_458)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_399),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_460),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_394),
.B(n_422),
.C(n_418),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_439),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_465),
.B(n_486),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_466),
.A2(n_472),
.B1(n_461),
.B2(n_453),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_468),
.A2(n_493),
.B1(n_449),
.B2(n_444),
.Y(n_507)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_439),
.Y(n_469)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_469),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_447),
.A2(n_401),
.B1(n_393),
.B2(n_392),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_SL g497 ( 
.A(n_470),
.B(n_490),
.C(n_454),
.Y(n_497)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_471),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_456),
.A2(n_412),
.B1(n_413),
.B2(n_403),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_440),
.Y(n_473)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_473),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_434),
.A2(n_404),
.B(n_410),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_475),
.A2(n_480),
.B(n_484),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_451),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_404),
.C(n_409),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_479),
.C(n_444),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_446),
.B(n_404),
.C(n_410),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_438),
.A2(n_426),
.B(n_411),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_445),
.B(n_400),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_481),
.B(n_488),
.Y(n_499)
);

BUFx5_ASAP7_75t_L g482 ( 
.A(n_442),
.Y(n_482)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_487),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_416),
.B(n_400),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_436),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_414),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_489),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_435),
.A2(n_463),
.B1(n_430),
.B2(n_459),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_433),
.A2(n_458),
.B1(n_443),
.B2(n_455),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_430),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_494),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_495),
.A2(n_473),
.B1(n_482),
.B2(n_491),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_448),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_496),
.B(n_501),
.Y(n_539)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_497),
.Y(n_530)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_494),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_509),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_475),
.A2(n_432),
.B(n_450),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_503),
.A2(n_505),
.B(n_502),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_437),
.Y(n_505)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_505),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_507),
.A2(n_484),
.B1(n_469),
.B2(n_480),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_460),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_510),
.B(n_513),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_476),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_470),
.B(n_452),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_493),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_467),
.B(n_477),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_518),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_483),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_492),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_479),
.B(n_474),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_520),
.B(n_497),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_474),
.C(n_489),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_524),
.Y(n_542)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_525),
.B(n_526),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_498),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_492),
.C(n_468),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_531),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_504),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_533),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_499),
.B(n_478),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_499),
.B(n_478),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_506),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_534),
.A2(n_512),
.B1(n_508),
.B2(n_504),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_535),
.B(n_519),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_502),
.A2(n_491),
.B(n_503),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_536),
.A2(n_537),
.B(n_514),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_540),
.A2(n_548),
.B1(n_551),
.B2(n_528),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_543),
.B(n_544),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_547),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_520),
.B(n_518),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_534),
.A2(n_512),
.B1(n_508),
.B2(n_516),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_507),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_552),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_530),
.A2(n_519),
.B1(n_516),
.B2(n_498),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_521),
.B(n_496),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_535),
.A2(n_510),
.B1(n_511),
.B2(n_530),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_554),
.B(n_555),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_536),
.A2(n_537),
.B(n_532),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_526),
.A2(n_511),
.B(n_532),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_556),
.A2(n_522),
.B(n_525),
.Y(n_566)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_557),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_549),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_558),
.B(n_559),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_552),
.B(n_539),
.C(n_529),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_550),
.B(n_539),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_560),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_554),
.B(n_527),
.C(n_529),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_564),
.B(n_567),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_566),
.B(n_545),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_547),
.B(n_523),
.C(n_528),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_522),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_568),
.B(n_569),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_543),
.B(n_551),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_571),
.B(n_573),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_563),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_561),
.A2(n_544),
.B1(n_541),
.B2(n_556),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_574),
.B(n_565),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_566),
.B(n_541),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_575),
.Y(n_580)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_579),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_570),
.B(n_562),
.C(n_559),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_582),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_578),
.B(n_565),
.C(n_567),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_583),
.A2(n_577),
.B(n_571),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_581),
.Y(n_587)
);

O2A1O1Ixp33_ASAP7_75t_SL g589 ( 
.A1(n_587),
.A2(n_588),
.B(n_585),
.C(n_572),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_586),
.B(n_580),
.C(n_576),
.Y(n_588)
);

O2A1O1Ixp33_ASAP7_75t_L g590 ( 
.A1(n_589),
.A2(n_575),
.B(n_574),
.C(n_561),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_546),
.Y(n_591)
);


endmodule