module fake_jpeg_10239_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_71;
wire n_52;
wire n_68;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx2_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_13),
.B(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_25),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_3),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_23),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_23),
.B1(n_11),
.B2(n_19),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_16),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_21),
.B1(n_11),
.B2(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_43),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_12),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_45),
.B(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_51),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_9),
.B(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_40),
.B(n_36),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_55),
.B(n_18),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_34),
.B(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_9),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_9),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_61),
.C(n_58),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_18),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_52),
.B1(n_17),
.B2(n_15),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_41),
.B1(n_62),
.B2(n_31),
.Y(n_69)
);

OAI321xp33_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_62),
.A3(n_15),
.B1(n_32),
.B2(n_33),
.C(n_7),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_41),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_69),
.B(n_68),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);


endmodule