module fake_jpeg_1911_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_35),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_4),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_28),
.A2(n_26),
.B1(n_17),
.B2(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_71),
.Y(n_88)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx2_ASAP7_75t_SL g102 ( 
.A(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_85),
.Y(n_99)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_28),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_19),
.Y(n_85)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_50),
.B1(n_29),
.B2(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_66),
.A2(n_17),
.B1(n_22),
.B2(n_4),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_58),
.B1(n_55),
.B2(n_73),
.Y(n_109)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_98),
.Y(n_121)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_5),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_78),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_63),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_64),
.Y(n_119)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_68),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_57),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_58),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_55),
.B(n_69),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_89),
.B(n_93),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_60),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_125),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_67),
.B1(n_62),
.B2(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_56),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_133),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_139),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_138),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_105),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_139),
.B(n_140),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_143),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_112),
.B(n_116),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_149),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_150),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_118),
.B1(n_100),
.B2(n_122),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_141),
.B1(n_117),
.B2(n_121),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_117),
.B(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

NAND4xp25_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_153),
.C(n_141),
.D(n_98),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_137),
.C(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_159),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_157),
.A2(n_141),
.B1(n_154),
.B2(n_156),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_137),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_146),
.C(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_101),
.B(n_90),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_121),
.C(n_122),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_159),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_167),
.B(n_166),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_154),
.B(n_101),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_171),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_91),
.B(n_87),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_92),
.C(n_95),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_173),
.B(n_100),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_102),
.Y(n_176)
);


endmodule