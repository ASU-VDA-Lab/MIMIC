module fake_jpeg_4264_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_25),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

OR2x4_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_20),
.Y(n_47)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_20),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_43),
.Y(n_68)
);

NAND2x1_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_27),
.A2(n_13),
.B1(n_23),
.B2(n_19),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_24),
.B1(n_21),
.B2(n_12),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_62),
.B1(n_3),
.B2(n_6),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_60),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_20),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_42),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_29),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_69),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_34),
.B1(n_29),
.B2(n_38),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_13),
.B1(n_19),
.B2(n_17),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_17),
.B1(n_37),
.B2(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_16),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_40),
.B1(n_39),
.B2(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_77),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_8),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_52),
.B1(n_67),
.B2(n_59),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_68),
.B(n_65),
.C(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_51),
.B(n_54),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_71),
.B(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_69),
.B1(n_64),
.B2(n_75),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_85),
.B(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_52),
.B1(n_59),
.B2(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_80),
.B1(n_83),
.B2(n_81),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_68),
.C(n_76),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_89),
.C(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_101),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_108),
.B(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_100),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_93),
.C(n_89),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_101),
.A3(n_102),
.B1(n_103),
.B2(n_96),
.C1(n_99),
.C2(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_114),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_110),
.B1(n_109),
.B2(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_91),
.C(n_53),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_112),
.C(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_120),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_118),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_116),
.C(n_10),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_121),
.C(n_8),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_58),
.Y(n_125)
);


endmodule