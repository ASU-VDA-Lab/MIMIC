module fake_netlist_6_1598_n_2088 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2088);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2088;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_292;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_79),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_24),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_148),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_27),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_71),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_126),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_84),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_138),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_89),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_140),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_10),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_103),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_119),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_69),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_42),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_129),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_41),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_14),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_45),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_84),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_123),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_19),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_150),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_39),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_56),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_132),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_141),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_67),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_35),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_178),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_79),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_86),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_81),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_73),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_192),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_120),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_164),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_18),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_80),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_70),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_156),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_92),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_133),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_149),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_20),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_60),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_73),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_155),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_107),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_173),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_89),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_161),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_196),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_24),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_99),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_101),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_162),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_66),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_124),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_65),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_11),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_135),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_80),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_17),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_166),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_83),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_35),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_55),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_122),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_47),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_105),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_60),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_151),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_66),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_88),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_20),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_113),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_17),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_58),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_94),
.Y(n_294)
);

BUFx2_ASAP7_75t_SL g295 ( 
.A(n_98),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_97),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_186),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_44),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_152),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_23),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_159),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_54),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_56),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_47),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_1),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_183),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_108),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_62),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_49),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_33),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_130),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_74),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_172),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_8),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_96),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_8),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_58),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_147),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_116),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_4),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_21),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_76),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_131),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_184),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_36),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_16),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_16),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_181),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_49),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_40),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_0),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_22),
.Y(n_333)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_179),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_69),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_59),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_90),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_88),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_127),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_23),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_19),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_72),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_9),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_44),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_194),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_174),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_191),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_54),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_154),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_93),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_100),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_48),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_187),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_182),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_52),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_144),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_117),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_45),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_75),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_11),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_15),
.Y(n_361)
);

HB1xp67_ASAP7_75t_SL g362 ( 
.A(n_21),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_77),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_77),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_115),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_165),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_40),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_50),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_82),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_163),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_1),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_175),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_171),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_7),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_139),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_137),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_18),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_46),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_146),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_50),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_71),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_95),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_180),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_114),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_36),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_9),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_86),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_10),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_169),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_102),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_81),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_91),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_205),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_230),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_290),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_197),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_201),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_257),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_263),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_202),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_222),
.B(n_0),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_257),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_226),
.B(n_2),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_303),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_257),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_248),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_253),
.B(n_3),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_303),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_248),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_208),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_264),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_248),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_279),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_279),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_237),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_279),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_210),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_353),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_312),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_388),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_366),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_200),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_375),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_222),
.B(n_3),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_200),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_211),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_214),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_226),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_275),
.B(n_4),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_215),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_229),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_229),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_203),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_322),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_198),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_292),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_253),
.B(n_5),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_219),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_232),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_232),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_227),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_242),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_203),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_242),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_231),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_247),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_247),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_243),
.B(n_5),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_240),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_236),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_249),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_249),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_246),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_252),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_204),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_265),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_259),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_266),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_268),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_265),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_269),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_271),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_274),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_267),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_277),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_283),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_267),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_272),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_272),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_278),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_392),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_392),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_285),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_300),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_308),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_316),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_320),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_278),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_281),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_325),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_337),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_281),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_204),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_345),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_286),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_326),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_286),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_289),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_289),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_396),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_397),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_400),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_393),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_410),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_430),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_R g499 ( 
.A(n_417),
.B(n_346),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_430),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_428),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_429),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_421),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_394),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_431),
.B(n_245),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_433),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_398),
.A2(n_244),
.B(n_234),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_433),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_432),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_441),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_453),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_461),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_462),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_464),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_476),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_398),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_409),
.B(n_243),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_402),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_405),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_R g530 ( 
.A(n_477),
.B(n_347),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_409),
.B(n_280),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_479),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_412),
.B(n_296),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_492),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_412),
.B(n_280),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_480),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_445),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_447),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_399),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_447),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_439),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_449),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_449),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_403),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_450),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_450),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_454),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_411),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_419),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_458),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_454),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_455),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_440),
.B(n_451),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_444),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_459),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_448),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_456),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_459),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_457),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_460),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_463),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_465),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_R g568 ( 
.A(n_466),
.B(n_349),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_463),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_424),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_531),
.B(n_280),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_514),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_545),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_545),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_514),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_504),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_557),
.B(n_413),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_503),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_557),
.B(n_407),
.C(n_548),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_504),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_548),
.B(n_437),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_572),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_498),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_498),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_531),
.B(n_287),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_552),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_552),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_500),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_548),
.B(n_531),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_506),
.B(n_468),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_548),
.B(n_458),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_500),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_506),
.B(n_469),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_507),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_531),
.B(n_287),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_503),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_507),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_510),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_510),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_548),
.A2(n_475),
.B1(n_474),
.B2(n_452),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_504),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_568),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_537),
.B(n_478),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_572),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_568),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_512),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_537),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_503),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_493),
.A2(n_415),
.B1(n_484),
.B2(n_483),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_531),
.B(n_287),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

INVx6_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_553),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_534),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_508),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_535),
.B(n_296),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_553),
.B(n_423),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_508),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_559),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_535),
.B(n_339),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_508),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_526),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_512),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_519),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_535),
.B(n_234),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_535),
.B(n_225),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_534),
.B(n_234),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_494),
.B(n_487),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_495),
.B(n_489),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_554),
.B(n_436),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_519),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_569),
.B(n_225),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_525),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_534),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_534),
.B(n_258),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_497),
.B(n_489),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_569),
.B(n_244),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_496),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_525),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_501),
.B(n_427),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_527),
.B(n_339),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_534),
.B(n_244),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_R g654 ( 
.A(n_561),
.B(n_425),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_527),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_534),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_526),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_536),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_526),
.Y(n_659)
);

INVx4_ASAP7_75t_SL g660 ( 
.A(n_526),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_526),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_569),
.B(n_319),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_502),
.B(n_427),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_509),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_562),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_526),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_536),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_538),
.Y(n_668)
);

NAND3x1_ASAP7_75t_L g669 ( 
.A(n_524),
.B(n_451),
.C(n_321),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_538),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_541),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_541),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_511),
.B(n_435),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_542),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_554),
.B(n_436),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_505),
.Y(n_677)
);

AND3x4_ASAP7_75t_L g678 ( 
.A(n_564),
.B(n_426),
.C(n_401),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_542),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_546),
.Y(n_680)
);

AND2x6_ASAP7_75t_L g681 ( 
.A(n_569),
.B(n_258),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_569),
.B(n_319),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_509),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_546),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_522),
.B(n_350),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_547),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_499),
.B(n_258),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_499),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_522),
.B(n_350),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_547),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_550),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_529),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_529),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_550),
.B(n_258),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_522),
.B(n_382),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_513),
.B(n_446),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_509),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_555),
.Y(n_698)
);

INVx6_ASAP7_75t_L g699 ( 
.A(n_529),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_524),
.B(n_403),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_529),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_515),
.B(n_516),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_529),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_558),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_558),
.B(n_258),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_522),
.B(n_382),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_529),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_560),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_530),
.B(n_258),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_560),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_563),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_563),
.B(n_339),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_570),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_509),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_570),
.B(n_413),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_571),
.B(n_414),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_565),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_517),
.B(n_486),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_571),
.B(n_414),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_509),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_540),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_540),
.Y(n_723)
);

INVx4_ASAP7_75t_SL g724 ( 
.A(n_522),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_518),
.B(n_521),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_622),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_581),
.B(n_532),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_581),
.B(n_539),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_697),
.A2(n_533),
.B(n_206),
.Y(n_729)
);

AND2x2_ASAP7_75t_SL g730 ( 
.A(n_598),
.B(n_601),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_716),
.B(n_199),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_683),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_588),
.B(n_395),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_583),
.B(n_533),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_635),
.A2(n_206),
.B1(n_212),
.B2(n_199),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_716),
.B(n_212),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_573),
.B(n_530),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_622),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_688),
.B(n_567),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_599),
.B(n_404),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_622),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_575),
.B(n_578),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_597),
.A2(n_544),
.B(n_540),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_640),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_580),
.B(n_544),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_622),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_584),
.B(n_544),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_579),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_L g749 ( 
.A1(n_664),
.A2(n_235),
.B(n_260),
.C(n_254),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_599),
.B(n_408),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_635),
.A2(n_235),
.B1(n_260),
.B2(n_254),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_587),
.B(n_683),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_669),
.A2(n_216),
.B1(n_426),
.B2(n_401),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_SL g754 ( 
.A(n_688),
.B(n_245),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_579),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_654),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_683),
.B(n_549),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_697),
.A2(n_551),
.B(n_549),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_683),
.B(n_549),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_635),
.A2(n_314),
.B1(n_291),
.B2(n_294),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_586),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_586),
.Y(n_762)
);

O2A1O1Ixp5_ASAP7_75t_L g763 ( 
.A1(n_664),
.A2(n_365),
.B(n_351),
.C(n_329),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_683),
.B(n_551),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_636),
.A2(n_389),
.B1(n_291),
.B2(n_294),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_715),
.B(n_551),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_651),
.B(n_543),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_635),
.A2(n_324),
.B1(n_351),
.B2(n_297),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_715),
.B(n_556),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_640),
.B(n_676),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_715),
.B(n_556),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_715),
.B(n_556),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_676),
.B(n_322),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_617),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_635),
.A2(n_297),
.B1(n_329),
.B2(n_383),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_641),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_715),
.B(n_566),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_635),
.A2(n_376),
.B1(n_314),
.B2(n_383),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_701),
.A2(n_365),
.B1(n_307),
.B2(n_324),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_611),
.B(n_354),
.Y(n_780)
);

OR2x6_ASAP7_75t_L g781 ( 
.A(n_701),
.B(n_295),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_701),
.A2(n_376),
.B1(n_307),
.B2(n_295),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_590),
.B(n_566),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_591),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_610),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_617),
.B(n_368),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_663),
.B(n_368),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_669),
.A2(n_276),
.B1(n_220),
.B2(n_282),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_611),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_614),
.B(n_356),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_614),
.B(n_357),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_701),
.A2(n_313),
.B1(n_340),
.B2(n_364),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_589),
.B(n_416),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_648),
.B(n_312),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_596),
.B(n_566),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_716),
.B(n_416),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_673),
.B(n_207),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_642),
.B(n_302),
.C(n_370),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_610),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_613),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_600),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_628),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_648),
.B(n_312),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_602),
.B(n_528),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_606),
.B(n_528),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_629),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_664),
.A2(n_302),
.B1(n_312),
.B2(n_334),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_574),
.B(n_418),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_628),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_607),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_608),
.B(n_528),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_616),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_609),
.B(n_372),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_574),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_619),
.B(n_373),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_662),
.A2(n_682),
.B1(n_626),
.B2(n_721),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_721),
.A2(n_302),
.B1(n_312),
.B2(n_334),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_696),
.B(n_209),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_719),
.B(n_379),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_641),
.B(n_213),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_633),
.B(n_523),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_658),
.B(n_384),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_574),
.A2(n_284),
.B1(n_390),
.B2(n_228),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_717),
.B(n_418),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_721),
.A2(n_302),
.B1(n_312),
.B2(n_334),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_593),
.A2(n_302),
.B1(n_312),
.B2(n_334),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_625),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_634),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_643),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_650),
.B(n_523),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_655),
.B(n_667),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_668),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_625),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_671),
.B(n_523),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_672),
.B(n_302),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_658),
.B(n_245),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_674),
.B(n_312),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_679),
.B(n_312),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_670),
.B(n_245),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_684),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_625),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_686),
.B(n_334),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_690),
.B(n_334),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_670),
.A2(n_250),
.B1(n_224),
.B2(n_223),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_717),
.B(n_420),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_680),
.B(n_217),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_593),
.A2(n_334),
.B1(n_228),
.B2(n_330),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_680),
.B(n_218),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_691),
.B(n_334),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_698),
.B(n_334),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_720),
.B(n_420),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_700),
.B(n_422),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_705),
.B(n_422),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_709),
.B(n_470),
.Y(n_855)
);

O2A1O1Ixp5_ASAP7_75t_L g856 ( 
.A1(n_593),
.A2(n_492),
.B(n_491),
.C(n_490),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_711),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_631),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_712),
.B(n_470),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_604),
.A2(n_620),
.B1(n_630),
.B2(n_714),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_639),
.B(n_221),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_722),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_685),
.B(n_471),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_647),
.B(n_251),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_689),
.B(n_471),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_723),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_695),
.B(n_472),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_707),
.B(n_472),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_604),
.A2(n_336),
.B1(n_391),
.B2(n_310),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_SL g870 ( 
.A1(n_612),
.A2(n_251),
.B1(n_361),
.B2(n_360),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_631),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_604),
.A2(n_371),
.B(n_321),
.C(n_330),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_620),
.B(n_473),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_620),
.B(n_630),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_720),
.B(n_473),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_652),
.B(n_251),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_630),
.B(n_481),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_678),
.B(n_233),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_618),
.B(n_481),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_678),
.B(n_238),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_631),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_652),
.B(n_482),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_687),
.A2(n_239),
.B1(n_241),
.B2(n_387),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_637),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_687),
.A2(n_336),
.B(n_310),
.C(n_342),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_703),
.B(n_255),
.Y(n_886)
);

INVx8_ASAP7_75t_L g887 ( 
.A(n_648),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_652),
.A2(n_338),
.B1(n_256),
.B2(n_261),
.Y(n_888)
);

NOR3x1_ASAP7_75t_L g889 ( 
.A(n_710),
.B(n_342),
.C(n_348),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_618),
.B(n_482),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_618),
.B(n_713),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_725),
.B(n_262),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_713),
.B(n_251),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_713),
.B(n_485),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_710),
.B(n_638),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_632),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_649),
.B(n_270),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_774),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_774),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_727),
.B(n_677),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_808),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_808),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_SL g903 ( 
.A(n_878),
.B(n_288),
.C(n_273),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_824),
.B(n_629),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_734),
.B(n_656),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_734),
.B(n_656),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_770),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_732),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_732),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_732),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_732),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_800),
.Y(n_912)
);

BUFx4f_ASAP7_75t_SL g913 ( 
.A(n_739),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_808),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_732),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_728),
.B(n_724),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_887),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_776),
.B(n_724),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_863),
.B(n_656),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_800),
.Y(n_920)
);

AND2x2_ASAP7_75t_SL g921 ( 
.A(n_730),
.B(n_348),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_887),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_865),
.B(n_867),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_808),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_748),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_SL g926 ( 
.A(n_787),
.B(n_577),
.C(n_576),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_744),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_862),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_862),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_866),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_806),
.Y(n_931)
);

INVx3_ASAP7_75t_SL g932 ( 
.A(n_806),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_776),
.B(n_724),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_868),
.B(n_784),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_866),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_880),
.B(n_298),
.C(n_293),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_784),
.B(n_801),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_726),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_748),
.Y(n_939)
);

BUFx4_ASAP7_75t_SL g940 ( 
.A(n_756),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_887),
.Y(n_941)
);

BUFx8_ASAP7_75t_L g942 ( 
.A(n_744),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_801),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_810),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_726),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_810),
.B(n_582),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_824),
.B(n_665),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_730),
.A2(n_359),
.B(n_369),
.C(n_371),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_812),
.B(n_582),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_852),
.B(n_724),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_730),
.B(n_582),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_845),
.B(n_665),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_812),
.B(n_582),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_887),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_887),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_833),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_755),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_833),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_828),
.Y(n_959)
);

AND2x2_ASAP7_75t_SL g960 ( 
.A(n_754),
.B(n_359),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_SL g961 ( 
.A(n_895),
.B(n_718),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_860),
.B(n_582),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_755),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_828),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_814),
.B(n_585),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_829),
.B(n_585),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_829),
.B(n_585),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_886),
.B(n_595),
.C(n_594),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_832),
.B(n_585),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_814),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_833),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_832),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_738),
.B(n_585),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_738),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_874),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_SL g976 ( 
.A(n_789),
.B(n_301),
.C(n_299),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_L g977 ( 
.A(n_892),
.B(n_623),
.C(n_718),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_840),
.B(n_603),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_875),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_797),
.A2(n_648),
.B1(n_621),
.B2(n_624),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_840),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_852),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_857),
.Y(n_983)
);

OR2x6_ASAP7_75t_SL g984 ( 
.A(n_789),
.B(n_304),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_882),
.B(n_648),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_818),
.B(n_627),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_875),
.Y(n_987)
);

BUFx4f_ASAP7_75t_L g988 ( 
.A(n_781),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_741),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_857),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_752),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_745),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_882),
.B(n_796),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_754),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_SL g995 ( 
.A(n_782),
.B(n_645),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_756),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_845),
.B(n_603),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_851),
.B(n_796),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_747),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_851),
.B(n_603),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_761),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_731),
.A2(n_648),
.B1(n_637),
.B2(n_653),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_882),
.B(n_603),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_742),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_770),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_873),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_877),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_882),
.B(n_603),
.Y(n_1008)
);

NOR2xp67_ASAP7_75t_L g1009 ( 
.A(n_798),
.B(n_897),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_731),
.A2(n_653),
.B1(n_621),
.B2(n_624),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_741),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_761),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_879),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_SL g1014 ( 
.A(n_737),
.B(n_645),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_746),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_746),
.B(n_592),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_890),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_762),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_757),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_762),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_759),
.B(n_605),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_764),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_816),
.B(n_605),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_896),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_766),
.B(n_605),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_785),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_769),
.B(n_605),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_785),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_731),
.B(n_632),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_799),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_896),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_781),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_799),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_733),
.A2(n_592),
.B1(n_661),
.B2(n_675),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_802),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_773),
.B(n_627),
.Y(n_1036)
);

BUFx12f_ASAP7_75t_L g1037 ( 
.A(n_786),
.Y(n_1037)
);

AO22x1_ASAP7_75t_L g1038 ( 
.A1(n_889),
.A2(n_861),
.B1(n_750),
.B2(n_740),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_781),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_729),
.B(n_605),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_767),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_786),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_771),
.B(n_615),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_802),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_809),
.Y(n_1045)
);

INVx8_ASAP7_75t_L g1046 ( 
.A(n_781),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_772),
.B(n_615),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_777),
.B(n_615),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_809),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_773),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_SL g1051 ( 
.A(n_844),
.B(n_311),
.C(n_381),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_871),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_884),
.B(n_615),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_827),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_SL g1055 ( 
.A(n_815),
.B(n_309),
.C(n_358),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_731),
.B(n_644),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_736),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_792),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_793),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_827),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_L g1061 ( 
.A(n_780),
.B(n_661),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_793),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_871),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_841),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_819),
.B(n_592),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_779),
.B(n_306),
.C(n_305),
.Y(n_1066)
);

CKINVDCx6p67_ASAP7_75t_R g1067 ( 
.A(n_790),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_891),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_792),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_841),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_881),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_831),
.B(n_615),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_881),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_SL g1074 ( 
.A(n_883),
.B(n_315),
.C(n_355),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_783),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_791),
.B(n_820),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_894),
.B(n_661),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_736),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_884),
.B(n_645),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_846),
.B(n_317),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_743),
.B(n_645),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_736),
.B(n_675),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_736),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_753),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_788),
.B(n_485),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_788),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_848),
.B(n_675),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_795),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_804),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_805),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_811),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1081),
.A2(n_758),
.B(n_821),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_991),
.B(n_830),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1086),
.A2(n_870),
.B1(n_765),
.B2(n_823),
.C(n_753),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_923),
.B(n_855),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_948),
.A2(n_872),
.A3(n_835),
.B(n_838),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1052),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_912),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_951),
.A2(n_763),
.B(n_749),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_951),
.A2(n_817),
.B(n_807),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_986),
.B(n_900),
.C(n_1086),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1021),
.A2(n_858),
.B(n_803),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1004),
.B(n_859),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_904),
.B(n_888),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_948),
.A2(n_1027),
.A3(n_1043),
.B(n_1025),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1063),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_898),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1081),
.A2(n_834),
.B(n_837),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1040),
.A2(n_843),
.B(n_842),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_SL g1110 ( 
.A1(n_921),
.A2(n_825),
.B(n_876),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_SL g1111 ( 
.A(n_1041),
.B(n_864),
.C(n_888),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_997),
.A2(n_856),
.B(n_798),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1047),
.A2(n_803),
.B(n_794),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_998),
.B(n_853),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_904),
.B(n_823),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_998),
.B(n_854),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_979),
.B(n_869),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1084),
.A2(n_760),
.B1(n_735),
.B2(n_751),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1048),
.A2(n_794),
.B(n_768),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_898),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_905),
.A2(n_849),
.A3(n_850),
.B(n_693),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1000),
.A2(n_813),
.B(n_826),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_907),
.B(n_893),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_925),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_921),
.A2(n_775),
.B1(n_778),
.B2(n_847),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_SL g1126 ( 
.A(n_931),
.B(n_326),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_979),
.B(n_836),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_947),
.B(n_889),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_906),
.A2(n_666),
.A3(n_659),
.B(n_657),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1042),
.B(n_839),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_937),
.A2(n_659),
.A3(n_666),
.B(n_657),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_987),
.B(n_822),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1071),
.A2(n_693),
.B(n_704),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1041),
.B(n_885),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_947),
.B(n_326),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_991),
.A2(n_699),
.B1(n_644),
.B2(n_704),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_993),
.B(n_1057),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_917),
.A2(n_645),
.B(n_646),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1005),
.B(n_318),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_987),
.B(n_692),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_919),
.A2(n_369),
.A3(n_380),
.B(n_391),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_960),
.A2(n_380),
.B(n_488),
.C(n_490),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_SL g1143 ( 
.A(n_917),
.B(n_488),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_917),
.A2(n_646),
.B(n_702),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_SL g1145 ( 
.A1(n_908),
.A2(n_491),
.B(n_109),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_917),
.A2(n_702),
.B(n_708),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_932),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1040),
.A2(n_708),
.B(n_692),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1071),
.A2(n_692),
.B(n_708),
.Y(n_1149)
);

AOI221x1_ASAP7_75t_L g1150 ( 
.A1(n_1014),
.A2(n_694),
.B1(n_706),
.B2(n_699),
.C(n_681),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_934),
.B(n_323),
.Y(n_1151)
);

OAI21xp33_ASAP7_75t_L g1152 ( 
.A1(n_1080),
.A2(n_1069),
.B(n_1058),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_917),
.A2(n_702),
.B(n_660),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_928),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_952),
.B(n_326),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_954),
.A2(n_955),
.B(n_908),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_929),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1071),
.A2(n_660),
.B(n_699),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_910),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_930),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1073),
.A2(n_660),
.B(n_699),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_1023),
.A2(n_660),
.B(n_681),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_918),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_L g1164 ( 
.A(n_926),
.B(n_386),
.C(n_385),
.Y(n_1164)
);

AOI21x1_ASAP7_75t_SL g1165 ( 
.A1(n_1087),
.A2(n_706),
.B(n_694),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1006),
.B(n_327),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_932),
.Y(n_1167)
);

AOI211x1_ASAP7_75t_L g1168 ( 
.A1(n_1038),
.A2(n_360),
.B(n_361),
.C(n_374),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_962),
.A2(n_681),
.B(n_694),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_954),
.A2(n_702),
.B(n_681),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1076),
.A2(n_681),
.B1(n_706),
.B2(n_694),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_SL g1172 ( 
.A(n_931),
.B(n_360),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_SL g1173 ( 
.A(n_977),
.B(n_378),
.C(n_377),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1073),
.A2(n_702),
.B(n_681),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_899),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1007),
.B(n_328),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_935),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_920),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_942),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1088),
.B(n_331),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1073),
.A2(n_706),
.B(n_694),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_954),
.A2(n_955),
.B(n_908),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1090),
.B(n_1091),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_925),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_992),
.B(n_332),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_962),
.A2(n_706),
.B(n_694),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_973),
.A2(n_706),
.B(n_195),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1075),
.A2(n_6),
.A3(n_12),
.B(n_13),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_952),
.B(n_360),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1050),
.B(n_333),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_1014),
.A2(n_6),
.B(n_12),
.Y(n_1191)
);

NAND3x1_ASAP7_75t_L g1192 ( 
.A(n_968),
.B(n_361),
.C(n_363),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_999),
.B(n_335),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1053),
.A2(n_193),
.B(n_190),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1075),
.B(n_367),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_954),
.A2(n_143),
.B(n_106),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1089),
.B(n_352),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_918),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_991),
.B(n_344),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_954),
.A2(n_955),
.B(n_1072),
.Y(n_1200)
);

AOI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1053),
.A2(n_188),
.B(n_170),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_SL g1202 ( 
.A1(n_1077),
.A2(n_361),
.B(n_22),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_973),
.A2(n_158),
.B(n_157),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_940),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1037),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1023),
.A2(n_343),
.B(n_341),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_993),
.B(n_1057),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1089),
.B(n_13),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_SL g1209 ( 
.A1(n_1079),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_943),
.B(n_25),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1016),
.A2(n_145),
.B(n_142),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_944),
.B(n_28),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_955),
.A2(n_136),
.B(n_121),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1016),
.A2(n_118),
.B(n_111),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_959),
.B(n_28),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_946),
.A2(n_110),
.B(n_104),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1046),
.B(n_29),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_955),
.A2(n_87),
.B(n_30),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_949),
.A2(n_966),
.B(n_953),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_910),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_910),
.A2(n_87),
.B(n_30),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_964),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_910),
.A2(n_85),
.B(n_31),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_991),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_991),
.B(n_32),
.Y(n_1225)
);

AOI21xp33_ASAP7_75t_L g1226 ( 
.A1(n_1058),
.A2(n_33),
.B(n_34),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_967),
.A2(n_978),
.B(n_969),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1065),
.A2(n_34),
.A3(n_37),
.B(n_38),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_972),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_993),
.B(n_37),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_985),
.B(n_38),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1013),
.A2(n_39),
.A3(n_41),
.B(n_42),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_SL g1233 ( 
.A(n_910),
.B(n_43),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_939),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1024),
.A2(n_43),
.B(n_46),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_994),
.B(n_48),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_981),
.Y(n_1237)
);

OAI22x1_ASAP7_75t_L g1238 ( 
.A1(n_1069),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_983),
.B(n_51),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1019),
.A2(n_53),
.B1(n_57),
.B2(n_59),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1017),
.A2(n_61),
.A3(n_62),
.B(n_63),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_SL g1242 ( 
.A1(n_956),
.A2(n_61),
.B(n_63),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1009),
.A2(n_961),
.B1(n_960),
.B2(n_1067),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_996),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_975),
.B(n_64),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_990),
.B(n_1019),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1018),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1003),
.A2(n_85),
.B(n_65),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1054),
.A2(n_64),
.A3(n_67),
.B(n_68),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1019),
.B(n_68),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1019),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1008),
.A2(n_83),
.B(n_76),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_980),
.A2(n_75),
.B(n_78),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_975),
.B(n_78),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1019),
.B(n_82),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1022),
.B(n_1078),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1024),
.A2(n_1031),
.B(n_965),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1085),
.A2(n_1062),
.B(n_1066),
.C(n_1074),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1101),
.B(n_1036),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1178),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1137),
.B(n_901),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1115),
.B(n_1059),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1126),
.A2(n_1036),
.B1(n_1037),
.B2(n_913),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1099),
.A2(n_1079),
.B(n_1020),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1178),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1133),
.A2(n_916),
.B(n_965),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1107),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1092),
.A2(n_916),
.B(n_1082),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1191),
.A2(n_1035),
.A3(n_1044),
.B(n_1045),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1149),
.A2(n_1060),
.B(n_1064),
.Y(n_1270)
);

OR2x4_ASAP7_75t_L g1271 ( 
.A(n_1111),
.B(n_1085),
.Y(n_1271)
);

OAI22x1_ASAP7_75t_L g1272 ( 
.A1(n_1243),
.A2(n_1032),
.B1(n_1039),
.B2(n_996),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1110),
.A2(n_995),
.B(n_1002),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1108),
.A2(n_1064),
.B(n_1054),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1147),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1137),
.B(n_902),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1124),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1137),
.B(n_924),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1095),
.A2(n_1183),
.B1(n_1103),
.B2(n_1094),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1184),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1145),
.A2(n_1011),
.B(n_1061),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1184),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1114),
.B(n_1022),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1234),
.Y(n_1284)
);

O2A1O1Ixp5_ASAP7_75t_SL g1285 ( 
.A1(n_1245),
.A2(n_1028),
.B(n_1031),
.C(n_1024),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1234),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1097),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1104),
.B(n_914),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1200),
.A2(n_1227),
.B(n_1219),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1111),
.A2(n_961),
.B1(n_1083),
.B2(n_1067),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1109),
.A2(n_1257),
.B(n_1161),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1172),
.A2(n_942),
.B1(n_988),
.B2(n_1046),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_SL g1293 ( 
.A1(n_1253),
.A2(n_1030),
.B(n_1033),
.C(n_939),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1158),
.A2(n_1060),
.B(n_1031),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1258),
.A2(n_903),
.B(n_936),
.C(n_1051),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1116),
.B(n_1022),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1113),
.A2(n_995),
.B(n_922),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1165),
.A2(n_1049),
.B(n_1001),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1164),
.A2(n_1083),
.B1(n_988),
.B2(n_975),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1119),
.A2(n_941),
.B(n_922),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1154),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1165),
.A2(n_1049),
.B(n_1001),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1157),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1236),
.A2(n_942),
.B1(n_988),
.B2(n_1046),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1160),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1236),
.A2(n_1046),
.B1(n_927),
.B2(n_1083),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1151),
.B(n_1022),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1093),
.A2(n_1012),
.B(n_1026),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1246),
.A2(n_982),
.B1(n_1083),
.B2(n_1022),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1106),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1128),
.B(n_985),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1152),
.A2(n_1055),
.B1(n_1083),
.B2(n_975),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1244),
.A2(n_984),
.B1(n_982),
.B2(n_945),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1098),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1177),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1156),
.A2(n_963),
.B(n_1012),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1163),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1134),
.A2(n_975),
.B1(n_985),
.B2(n_982),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1222),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1182),
.A2(n_957),
.B(n_1033),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1231),
.B(n_1056),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1229),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1148),
.A2(n_957),
.B(n_1030),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1163),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1134),
.A2(n_1029),
.B(n_1056),
.C(n_976),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1122),
.A2(n_1010),
.B(n_1034),
.Y(n_1326)
);

AOI21xp33_ASAP7_75t_L g1327 ( 
.A1(n_1190),
.A2(n_1056),
.B(n_1029),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1237),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1216),
.A2(n_1214),
.B(n_1211),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1180),
.B(n_982),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1102),
.A2(n_963),
.B(n_1026),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1175),
.B(n_982),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1247),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1140),
.Y(n_1334)
);

OR2x6_ASAP7_75t_SL g1335 ( 
.A(n_1224),
.B(n_984),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1231),
.B(n_1029),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1130),
.B(n_945),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1107),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1112),
.A2(n_918),
.B(n_950),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1187),
.A2(n_1015),
.B(n_974),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1256),
.B(n_1068),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_SL g1342 ( 
.A(n_1204),
.B(n_950),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_SL g1343 ( 
.A1(n_1233),
.A2(n_1011),
.B(n_956),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1131),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1159),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1203),
.A2(n_1015),
.B(n_974),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_R g1347 ( 
.A(n_1244),
.B(n_938),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1130),
.B(n_938),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1235),
.A2(n_1015),
.B(n_974),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1127),
.A2(n_945),
.B1(n_938),
.B2(n_970),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1231),
.B(n_1230),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1093),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1208),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1250),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1120),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1131),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1173),
.A2(n_989),
.B(n_971),
.C(n_958),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1131),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1174),
.A2(n_989),
.B(n_958),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1159),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1199),
.B(n_1068),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1100),
.A2(n_950),
.B(n_933),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1164),
.B(n_1068),
.C(n_1011),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1168),
.B(n_1068),
.C(n_970),
.Y(n_1364)
);

CKINVDCx8_ASAP7_75t_R g1365 ( 
.A(n_1204),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1207),
.B(n_933),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1138),
.A2(n_1194),
.B(n_1201),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1146),
.A2(n_989),
.B(n_958),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1144),
.A2(n_1153),
.B(n_1202),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1118),
.A2(n_941),
.B(n_922),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1226),
.A2(n_1068),
.B1(n_970),
.B2(n_945),
.C(n_938),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1159),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1159),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1199),
.A2(n_933),
.B(n_956),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1136),
.A2(n_1070),
.B(n_970),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1220),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1150),
.A2(n_1070),
.B(n_971),
.Y(n_1377)
);

OAI21xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1210),
.A2(n_971),
.B(n_911),
.Y(n_1378)
);

OAI221xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1135),
.A2(n_909),
.B1(n_911),
.B2(n_915),
.C(n_970),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1198),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1202),
.A2(n_909),
.B(n_911),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1170),
.A2(n_909),
.B(n_915),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1255),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1181),
.A2(n_915),
.B(n_922),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1125),
.A2(n_1070),
.B(n_922),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1198),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1230),
.B(n_1070),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1212),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1196),
.A2(n_941),
.B(n_1070),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1205),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1215),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1213),
.A2(n_941),
.B(n_1186),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_R g1393 ( 
.A(n_1167),
.B(n_941),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1123),
.B(n_1193),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1169),
.A2(n_1209),
.B(n_1254),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1245),
.A2(n_1254),
.B(n_1225),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1123),
.B(n_1185),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1206),
.A2(n_1132),
.B(n_1117),
.C(n_1142),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1190),
.Y(n_1399)
);

BUFx12f_ASAP7_75t_L g1400 ( 
.A(n_1217),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1220),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1173),
.A2(n_1189),
.B1(n_1155),
.B2(n_1139),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1230),
.B(n_1207),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1195),
.A2(n_1197),
.B(n_1162),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1220),
.B(n_1225),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1166),
.A2(n_1176),
.B(n_1171),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1220),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1131),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1207),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1142),
.B(n_1105),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1147),
.Y(n_1411)
);

OAI211xp5_ASAP7_75t_L g1412 ( 
.A1(n_1139),
.A2(n_1252),
.B(n_1248),
.C(n_1221),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1167),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1239),
.B(n_1105),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1141),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1238),
.A2(n_1217),
.B1(n_1251),
.B2(n_1240),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1129),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1141),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1217),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1223),
.A2(n_1218),
.B1(n_1242),
.B2(n_1179),
.C(n_1192),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1129),
.A2(n_1121),
.B(n_1162),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1129),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1141),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1129),
.A2(n_1121),
.B(n_1096),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1141),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1121),
.A2(n_1096),
.B(n_1105),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1105),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_SL g1428 ( 
.A1(n_1096),
.A2(n_1121),
.B(n_1249),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1179),
.B(n_1143),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1096),
.A2(n_1228),
.B1(n_1232),
.B2(n_1241),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1394),
.A2(n_1228),
.B1(n_1232),
.B2(n_1241),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1347),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1366),
.Y(n_1433)
);

NAND2xp33_ASAP7_75t_SL g1434 ( 
.A(n_1393),
.B(n_1228),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1411),
.Y(n_1435)
);

AO221x2_ASAP7_75t_L g1436 ( 
.A1(n_1272),
.A2(n_1273),
.B1(n_1313),
.B2(n_1279),
.C(n_1263),
.Y(n_1436)
);

AO31x2_ASAP7_75t_L g1437 ( 
.A1(n_1344),
.A2(n_1228),
.A3(n_1188),
.B(n_1249),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1397),
.A2(n_1232),
.B1(n_1241),
.B2(n_1188),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1411),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1314),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1399),
.A2(n_1232),
.B1(n_1241),
.B2(n_1188),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1259),
.A2(n_1416),
.B1(n_1388),
.B2(n_1391),
.C(n_1402),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1405),
.B(n_1249),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1411),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1262),
.B(n_1260),
.Y(n_1445)
);

CKINVDCx12_ASAP7_75t_R g1446 ( 
.A(n_1262),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1412),
.B(n_1188),
.C(n_1249),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1300),
.A2(n_1297),
.B(n_1349),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1265),
.B(n_1288),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1277),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1379),
.A2(n_1318),
.B1(n_1271),
.B2(n_1290),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1351),
.B(n_1409),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1365),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1337),
.A2(n_1348),
.B1(n_1272),
.B2(n_1288),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1354),
.B(n_1383),
.Y(n_1455)
);

AO32x2_ASAP7_75t_L g1456 ( 
.A1(n_1430),
.A2(n_1428),
.A3(n_1338),
.B1(n_1267),
.B2(n_1309),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1353),
.A2(n_1326),
.B1(n_1406),
.B2(n_1400),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1271),
.A2(n_1371),
.B1(n_1312),
.B2(n_1306),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1267),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1351),
.B(n_1409),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1400),
.A2(n_1419),
.B1(n_1335),
.B2(n_1413),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1325),
.A2(n_1295),
.B(n_1398),
.C(n_1327),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1345),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1370),
.A2(n_1293),
.B(n_1385),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1366),
.Y(n_1465)
);

CKINVDCx11_ASAP7_75t_R g1466 ( 
.A(n_1365),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1420),
.A2(n_1410),
.B1(n_1413),
.B2(n_1396),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1428),
.A2(n_1289),
.B(n_1375),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1410),
.A2(n_1396),
.B1(n_1296),
.B2(n_1283),
.Y(n_1469)
);

BUFx12f_ASAP7_75t_L g1470 ( 
.A(n_1390),
.Y(n_1470)
);

AOI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1307),
.A2(n_1330),
.B(n_1361),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1310),
.A2(n_1319),
.B1(n_1352),
.B2(n_1304),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1335),
.A2(n_1271),
.B1(n_1342),
.B2(n_1361),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1411),
.A2(n_1405),
.B1(n_1311),
.B2(n_1332),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1409),
.B(n_1403),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1319),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1315),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1338),
.B(n_1403),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1405),
.A2(n_1311),
.B1(n_1363),
.B2(n_1275),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1280),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1352),
.A2(n_1364),
.B1(n_1333),
.B2(n_1414),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1355),
.A2(n_1390),
.B1(n_1341),
.B2(n_1315),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1292),
.A2(n_1299),
.B1(n_1355),
.B2(n_1322),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_1341),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1322),
.A2(n_1328),
.B1(n_1301),
.B2(n_1303),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1334),
.B(n_1261),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1366),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1387),
.B(n_1321),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1333),
.A2(n_1305),
.B1(n_1328),
.B2(n_1321),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1345),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1336),
.A2(n_1387),
.B1(n_1261),
.B2(n_1278),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1282),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1349),
.A2(n_1329),
.B(n_1289),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1336),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1282),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1334),
.A2(n_1261),
.B1(n_1278),
.B2(n_1276),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1404),
.A2(n_1418),
.B1(n_1425),
.B2(n_1415),
.C(n_1423),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1276),
.A2(n_1278),
.B1(n_1429),
.B2(n_1350),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1329),
.A2(n_1367),
.B(n_1291),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1276),
.B(n_1380),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1415),
.A2(n_1425),
.B1(n_1423),
.B2(n_1427),
.Y(n_1501)
);

INVx4_ASAP7_75t_SL g1502 ( 
.A(n_1345),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1317),
.B(n_1380),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1284),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1317),
.B(n_1380),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1317),
.B(n_1324),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1427),
.A2(n_1395),
.B1(n_1362),
.B2(n_1286),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1284),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1372),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1286),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1324),
.B(n_1386),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1372),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1324),
.B(n_1386),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1395),
.A2(n_1362),
.B1(n_1339),
.B2(n_1386),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1373),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1373),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1376),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1362),
.B(n_1339),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1339),
.A2(n_1374),
.B1(n_1264),
.B2(n_1358),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1374),
.A2(n_1264),
.B1(n_1358),
.B2(n_1408),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1376),
.Y(n_1521)
);

NAND2x1_ASAP7_75t_L g1522 ( 
.A(n_1343),
.B(n_1281),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1407),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1407),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1360),
.B(n_1401),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1345),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1401),
.Y(n_1527)
);

NOR2xp67_ASAP7_75t_SL g1528 ( 
.A(n_1401),
.B(n_1264),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1401),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1269),
.B(n_1374),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1308),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1269),
.B(n_1357),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1344),
.A2(n_1356),
.B1(n_1408),
.B2(n_1417),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_R g1534 ( 
.A(n_1377),
.B(n_1392),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1308),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1356),
.A2(n_1417),
.B1(n_1422),
.B2(n_1281),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_SL g1537 ( 
.A1(n_1343),
.A2(n_1375),
.B(n_1422),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1426),
.A2(n_1424),
.B1(n_1378),
.B2(n_1331),
.Y(n_1538)
);

CKINVDCx11_ASAP7_75t_R g1539 ( 
.A(n_1269),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1377),
.A2(n_1285),
.B1(n_1269),
.B2(n_1381),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1389),
.A2(n_1392),
.B(n_1377),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1285),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1298),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1367),
.A2(n_1389),
.B1(n_1381),
.B2(n_1346),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1269),
.B(n_1426),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1424),
.B(n_1331),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1298),
.B(n_1302),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1302),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1274),
.Y(n_1549)
);

OR2x6_ASAP7_75t_L g1550 ( 
.A(n_1340),
.B(n_1346),
.Y(n_1550)
);

INVx4_ASAP7_75t_L g1551 ( 
.A(n_1384),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1323),
.A2(n_1268),
.B1(n_1421),
.B2(n_1274),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1268),
.A2(n_1266),
.B(n_1369),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1340),
.A2(n_1368),
.B1(n_1323),
.B2(n_1266),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1369),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1368),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1421),
.B(n_1320),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1384),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1382),
.Y(n_1559)
);

NOR3xp33_ASAP7_75t_SL g1560 ( 
.A(n_1382),
.B(n_1316),
.C(n_1320),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1316),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1270),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1359),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1359),
.A2(n_1291),
.B1(n_1270),
.B2(n_1294),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1294),
.A2(n_730),
.B1(n_1094),
.B2(n_960),
.Y(n_1565)
);

AOI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1394),
.A2(n_787),
.B1(n_797),
.B2(n_818),
.C(n_1397),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1394),
.A2(n_730),
.B1(n_1094),
.B2(n_960),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1366),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1275),
.Y(n_1569)
);

AO32x2_ASAP7_75t_L g1570 ( 
.A1(n_1279),
.A2(n_1251),
.A3(n_1240),
.B1(n_1224),
.B2(n_1430),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1394),
.B(n_730),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1424),
.A2(n_1426),
.B(n_1421),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1394),
.B(n_1397),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1394),
.A2(n_730),
.B1(n_1094),
.B2(n_960),
.Y(n_1574)
);

INVx4_ASAP7_75t_L g1575 ( 
.A(n_1411),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1262),
.B(n_1288),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1262),
.B(n_1288),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1394),
.B(n_730),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1411),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1262),
.B(n_1288),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1277),
.Y(n_1581)
);

NAND3x1_ASAP7_75t_L g1582 ( 
.A(n_1402),
.B(n_1243),
.C(n_1394),
.Y(n_1582)
);

CKINVDCx16_ASAP7_75t_R g1583 ( 
.A(n_1347),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1287),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1277),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1277),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1399),
.A2(n_730),
.B1(n_994),
.B2(n_1101),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1394),
.A2(n_730),
.B1(n_1094),
.B2(n_960),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1394),
.B(n_1397),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1493),
.A2(n_1499),
.B(n_1448),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1566),
.A2(n_1567),
.B1(n_1588),
.B2(n_1574),
.C(n_1442),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1573),
.A2(n_1589),
.B1(n_1583),
.B2(n_1571),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1567),
.A2(n_1588),
.B1(n_1574),
.B2(n_1571),
.Y(n_1593)
);

OAI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1457),
.A2(n_1578),
.B1(n_1462),
.B2(n_1587),
.C(n_1461),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1464),
.A2(n_1565),
.B(n_1578),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1576),
.B(n_1577),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1436),
.A2(n_1457),
.B1(n_1473),
.B2(n_1458),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1459),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1436),
.A2(n_1451),
.B1(n_1483),
.B2(n_1460),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1580),
.B(n_1469),
.Y(n_1600)
);

OAI211xp5_ASAP7_75t_L g1601 ( 
.A1(n_1431),
.A2(n_1565),
.B(n_1454),
.C(n_1467),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1553),
.A2(n_1564),
.B(n_1447),
.Y(n_1602)
);

OR2x6_ASAP7_75t_L g1603 ( 
.A(n_1522),
.B(n_1443),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1436),
.A2(n_1460),
.B1(n_1452),
.B2(n_1475),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1532),
.B(n_1484),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1455),
.B(n_1486),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1440),
.B(n_1446),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1582),
.A2(n_1482),
.B1(n_1432),
.B2(n_1498),
.Y(n_1608)
);

INVxp33_ASAP7_75t_L g1609 ( 
.A(n_1445),
.Y(n_1609)
);

OAI211xp5_ASAP7_75t_L g1610 ( 
.A1(n_1431),
.A2(n_1467),
.B(n_1438),
.C(n_1472),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1452),
.A2(n_1475),
.B1(n_1488),
.B2(n_1491),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1469),
.B(n_1488),
.Y(n_1612)
);

AO31x2_ASAP7_75t_L g1613 ( 
.A1(n_1540),
.A2(n_1441),
.A3(n_1561),
.B(n_1518),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1479),
.A2(n_1474),
.B1(n_1471),
.B2(n_1494),
.C(n_1496),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1488),
.A2(n_1433),
.B1(n_1568),
.B2(n_1465),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1489),
.B(n_1438),
.C(n_1496),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1476),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1466),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1435),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1434),
.A2(n_1489),
.B1(n_1485),
.B2(n_1481),
.C(n_1542),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1518),
.A2(n_1541),
.B(n_1556),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1582),
.A2(n_1487),
.B1(n_1516),
.B2(n_1470),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1449),
.B(n_1478),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1434),
.A2(n_1481),
.B1(n_1497),
.B2(n_1530),
.C(n_1507),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1437),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1539),
.A2(n_1516),
.B1(n_1500),
.B2(n_1470),
.Y(n_1626)
);

OAI211xp5_ASAP7_75t_L g1627 ( 
.A1(n_1539),
.A2(n_1466),
.B(n_1524),
.C(n_1584),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1443),
.B(n_1456),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1506),
.A2(n_1569),
.B1(n_1503),
.B2(n_1505),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1506),
.A2(n_1569),
.B1(n_1579),
.B2(n_1439),
.Y(n_1630)
);

AOI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1507),
.A2(n_1514),
.B1(n_1501),
.B2(n_1545),
.C(n_1521),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1443),
.B(n_1456),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1435),
.A2(n_1439),
.B1(n_1444),
.B2(n_1575),
.Y(n_1633)
);

OAI211xp5_ASAP7_75t_L g1634 ( 
.A1(n_1511),
.A2(n_1514),
.B(n_1523),
.C(n_1512),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1435),
.A2(n_1579),
.B1(n_1439),
.B2(n_1444),
.Y(n_1635)
);

OAI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1544),
.A2(n_1579),
.B1(n_1575),
.B2(n_1513),
.C(n_1554),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_L g1637 ( 
.A1(n_1515),
.A2(n_1517),
.B(n_1495),
.C(n_1492),
.Y(n_1637)
);

OAI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1509),
.A2(n_1548),
.B1(n_1480),
.B2(n_1508),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1504),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_SL g1640 ( 
.A(n_1555),
.B(n_1550),
.Y(n_1640)
);

NAND2xp33_ASAP7_75t_R g1641 ( 
.A(n_1548),
.B(n_1525),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1555),
.A2(n_1510),
.B1(n_1529),
.B2(n_1527),
.Y(n_1642)
);

AO31x2_ASAP7_75t_L g1643 ( 
.A1(n_1543),
.A2(n_1546),
.A3(n_1549),
.B(n_1535),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1490),
.B(n_1502),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1537),
.A2(n_1586),
.B1(n_1450),
.B2(n_1585),
.Y(n_1645)
);

OAI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1538),
.A2(n_1536),
.B1(n_1519),
.B2(n_1552),
.C(n_1560),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1501),
.A2(n_1533),
.B1(n_1519),
.B2(n_1536),
.C(n_1520),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1437),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1551),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1528),
.B(n_1552),
.C(n_1531),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1570),
.A2(n_1526),
.B1(n_1463),
.B2(n_1581),
.Y(n_1651)
);

INVx3_ASAP7_75t_SL g1652 ( 
.A(n_1502),
.Y(n_1652)
);

AO21x2_ASAP7_75t_L g1653 ( 
.A1(n_1562),
.A2(n_1468),
.B(n_1557),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1463),
.A2(n_1526),
.B1(n_1550),
.B2(n_1551),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1550),
.A2(n_1551),
.B1(n_1558),
.B2(n_1547),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1563),
.A2(n_1559),
.B1(n_1570),
.B2(n_1502),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1563),
.A2(n_1570),
.B1(n_1572),
.B2(n_1456),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1570),
.A2(n_1534),
.B1(n_1563),
.B2(n_1572),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1572),
.A2(n_730),
.B1(n_1566),
.B2(n_1436),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1534),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1437),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1576),
.B(n_1577),
.Y(n_1664)
);

OAI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1566),
.A2(n_870),
.B(n_787),
.C(n_788),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1566),
.A2(n_994),
.B1(n_1574),
.B2(n_1567),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1566),
.A2(n_994),
.B1(n_1574),
.B2(n_1567),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1566),
.A2(n_787),
.B1(n_1588),
.B2(n_1574),
.C(n_1567),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1459),
.Y(n_1670)
);

OAI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1566),
.A2(n_994),
.B1(n_754),
.B2(n_1573),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1436),
.A2(n_730),
.B1(n_994),
.B2(n_960),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1674)
);

BUFx4_ASAP7_75t_R g1675 ( 
.A(n_1569),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1436),
.A2(n_730),
.B1(n_994),
.B2(n_960),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1576),
.B(n_1577),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1477),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1461),
.A2(n_1041),
.B1(n_994),
.B2(n_1573),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1555),
.Y(n_1683)
);

NOR3xp33_ASAP7_75t_L g1684 ( 
.A(n_1566),
.B(n_986),
.C(n_601),
.Y(n_1684)
);

OAI22x1_ASAP7_75t_L g1685 ( 
.A1(n_1454),
.A2(n_1571),
.B1(n_1578),
.B2(n_1402),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1477),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1477),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1566),
.A2(n_986),
.B1(n_598),
.B2(n_601),
.C(n_870),
.Y(n_1689)
);

NAND5xp2_ASAP7_75t_L g1690 ( 
.A(n_1566),
.B(n_1567),
.C(n_1588),
.D(n_1574),
.E(n_1094),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1566),
.A2(n_994),
.B1(n_1574),
.B2(n_1567),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1436),
.A2(n_730),
.B1(n_994),
.B2(n_960),
.Y(n_1693)
);

BUFx8_ASAP7_75t_L g1694 ( 
.A(n_1470),
.Y(n_1694)
);

AOI222xp33_ASAP7_75t_L g1695 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1567),
.B2(n_1588),
.C1(n_1574),
.C2(n_1094),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1532),
.B(n_1427),
.Y(n_1696)
);

AOI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1566),
.A2(n_730),
.B(n_1462),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1566),
.A2(n_787),
.B1(n_1588),
.B2(n_1574),
.C(n_1567),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1566),
.A2(n_986),
.B1(n_730),
.B2(n_1041),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1566),
.A2(n_994),
.B1(n_1574),
.B2(n_1567),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1461),
.A2(n_1041),
.B1(n_994),
.B2(n_1573),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_R g1702 ( 
.A(n_1453),
.B(n_654),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1522),
.B(n_1443),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1566),
.A2(n_787),
.B1(n_1588),
.B2(n_1574),
.C(n_1567),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1566),
.A2(n_730),
.B(n_787),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1576),
.B(n_1577),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1566),
.A2(n_994),
.B1(n_1574),
.B2(n_1567),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1566),
.A2(n_730),
.B1(n_1436),
.B2(n_1567),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1689),
.A2(n_1684),
.B1(n_1708),
.B2(n_1690),
.C(n_1591),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1628),
.B(n_1632),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_SL g1715 ( 
.A(n_1603),
.B(n_1703),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1628),
.B(n_1632),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1613),
.B(n_1605),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1643),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1605),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1656),
.B(n_1658),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1656),
.B(n_1653),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1653),
.B(n_1613),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1696),
.B(n_1606),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1696),
.B(n_1639),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1613),
.B(n_1602),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1613),
.B(n_1625),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1613),
.B(n_1648),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1662),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1603),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1612),
.B(n_1602),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1655),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1602),
.B(n_1621),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1612),
.B(n_1600),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1649),
.B(n_1661),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1603),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1661),
.B(n_1631),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1703),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1647),
.B(n_1657),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1659),
.B(n_1650),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1703),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1624),
.B(n_1595),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1646),
.B(n_1651),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1680),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1592),
.B(n_1697),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1590),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1640),
.B(n_1683),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1686),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1668),
.A2(n_1698),
.B1(n_1707),
.B2(n_1695),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1590),
.Y(n_1749)
);

INVxp67_ASAP7_75t_SL g1750 ( 
.A(n_1687),
.Y(n_1750)
);

NOR2x1p5_ASAP7_75t_L g1751 ( 
.A(n_1616),
.B(n_1683),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1670),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1620),
.B(n_1617),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1637),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1660),
.B(n_1654),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1623),
.B(n_1609),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1598),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1596),
.B(n_1664),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1645),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1598),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1634),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1636),
.Y(n_1762)
);

OAI21xp33_ASAP7_75t_L g1763 ( 
.A1(n_1665),
.A2(n_1712),
.B(n_1663),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1685),
.B(n_1638),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1685),
.B(n_1609),
.Y(n_1765)
);

OAI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1713),
.A2(n_1597),
.B1(n_1699),
.B2(n_1693),
.C(n_1676),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1745),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1719),
.B(n_1601),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1713),
.B(n_1671),
.C(n_1594),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1718),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1741),
.A2(n_1711),
.B1(n_1667),
.B2(n_1666),
.C(n_1691),
.Y(n_1771)
);

NOR4xp25_ASAP7_75t_SL g1772 ( 
.A(n_1761),
.B(n_1641),
.C(n_1702),
.D(n_1618),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_SL g1773 ( 
.A(n_1744),
.B(n_1741),
.C(n_1748),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_R g1774 ( 
.A(n_1762),
.B(n_1618),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1719),
.B(n_1709),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1743),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1760),
.Y(n_1777)
);

OR2x6_ASAP7_75t_L g1778 ( 
.A(n_1729),
.B(n_1610),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1743),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1741),
.A2(n_1700),
.B1(n_1706),
.B2(n_1705),
.C(n_1704),
.Y(n_1780)
);

OAI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1741),
.A2(n_1673),
.B(n_1677),
.C(n_1692),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1763),
.A2(n_1710),
.B1(n_1672),
.B2(n_1669),
.C(n_1678),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1744),
.A2(n_1674),
.B1(n_1682),
.B2(n_1688),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1763),
.A2(n_1593),
.B1(n_1701),
.B2(n_1681),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1714),
.B(n_1709),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1760),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1763),
.A2(n_1599),
.B1(n_1614),
.B2(n_1608),
.Y(n_1787)
);

OAI211xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1765),
.A2(n_1622),
.B(n_1642),
.C(n_1627),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1714),
.B(n_1679),
.Y(n_1789)
);

AOI21xp33_ASAP7_75t_L g1790 ( 
.A1(n_1754),
.A2(n_1629),
.B(n_1626),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1729),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

NAND4xp25_ASAP7_75t_L g1793 ( 
.A(n_1748),
.B(n_1753),
.C(n_1761),
.D(n_1762),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1718),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1743),
.Y(n_1795)
);

AOI211xp5_ASAP7_75t_L g1796 ( 
.A1(n_1748),
.A2(n_1607),
.B(n_1652),
.C(n_1679),
.Y(n_1796)
);

AOI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1736),
.A2(n_1604),
.B1(n_1611),
.B2(n_1615),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1717),
.B(n_1630),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1723),
.B(n_1635),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1746),
.Y(n_1800)
);

OAI21xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1736),
.A2(n_1675),
.B(n_1633),
.Y(n_1801)
);

AO21x2_ASAP7_75t_L g1802 ( 
.A1(n_1749),
.A2(n_1644),
.B(n_1675),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1747),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1729),
.Y(n_1804)
);

OAI31xp33_ASAP7_75t_L g1805 ( 
.A1(n_1751),
.A2(n_1644),
.A3(n_1694),
.B(n_1652),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1723),
.B(n_1619),
.Y(n_1806)
);

INVxp67_ASAP7_75t_SL g1807 ( 
.A(n_1754),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1747),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1714),
.B(n_1644),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1716),
.B(n_1694),
.Y(n_1810)
);

AOI33xp33_ASAP7_75t_L g1811 ( 
.A1(n_1736),
.A2(n_1761),
.A3(n_1762),
.B1(n_1738),
.B2(n_1730),
.B3(n_1722),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1736),
.A2(n_1764),
.B1(n_1738),
.B2(n_1753),
.C(n_1765),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1738),
.A2(n_1751),
.B1(n_1764),
.B2(n_1755),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1716),
.B(n_1733),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1738),
.A2(n_1751),
.B1(n_1755),
.B2(n_1742),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1732),
.B(n_1739),
.C(n_1742),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1755),
.A2(n_1742),
.B1(n_1759),
.B2(n_1756),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1792),
.B(n_1717),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1773),
.A2(n_1755),
.B1(n_1739),
.B2(n_1730),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1814),
.B(n_1730),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1807),
.B(n_1717),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1816),
.B(n_1752),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1800),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1776),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1785),
.B(n_1730),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1776),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1798),
.B(n_1721),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1816),
.B(n_1752),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1779),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1785),
.B(n_1721),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1789),
.B(n_1721),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1811),
.B(n_1733),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1800),
.B(n_1733),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1770),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1770),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1798),
.B(n_1733),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1775),
.B(n_1732),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1779),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1795),
.B(n_1750),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1775),
.B(n_1732),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1795),
.B(n_1750),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1791),
.B(n_1725),
.Y(n_1842)
);

INVx2_ASAP7_75t_SL g1843 ( 
.A(n_1800),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1803),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1804),
.B(n_1720),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1804),
.B(n_1720),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1804),
.B(n_1725),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1803),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1804),
.B(n_1720),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1804),
.B(n_1725),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1808),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1804),
.B(n_1720),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1809),
.B(n_1722),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1806),
.B(n_1756),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1768),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1768),
.B(n_1727),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1806),
.B(n_1756),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1767),
.B(n_1722),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1802),
.B(n_1724),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1824),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1855),
.B(n_1812),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1834),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1845),
.B(n_1802),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1824),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1855),
.B(n_1726),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1822),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1826),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1832),
.B(n_1793),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1826),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1829),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1856),
.B(n_1726),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1829),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1838),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1838),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1844),
.Y(n_1875)
);

OAI31xp33_ASAP7_75t_L g1876 ( 
.A1(n_1819),
.A2(n_1769),
.A3(n_1766),
.B(n_1781),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1818),
.Y(n_1877)
);

O2A1O1Ixp5_ASAP7_75t_L g1878 ( 
.A1(n_1822),
.A2(n_1828),
.B(n_1782),
.C(n_1832),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1856),
.B(n_1726),
.Y(n_1879)
);

INVxp67_ASAP7_75t_SL g1880 ( 
.A(n_1828),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1844),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1827),
.B(n_1794),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1821),
.B(n_1726),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1845),
.B(n_1802),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1802),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1848),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1834),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1846),
.B(n_1767),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1848),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1834),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1835),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1846),
.B(n_1767),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1821),
.B(n_1727),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1823),
.B(n_1767),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1835),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1846),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1823),
.B(n_1843),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1851),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1851),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1823),
.B(n_1715),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1849),
.B(n_1722),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1896),
.B(n_1849),
.Y(n_1902)
);

AOI32xp33_ASAP7_75t_L g1903 ( 
.A1(n_1868),
.A2(n_1784),
.A3(n_1813),
.B1(n_1815),
.B2(n_1787),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_L g1904 ( 
.A(n_1878),
.B(n_1793),
.C(n_1788),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1868),
.B(n_1827),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1866),
.B(n_1837),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1896),
.B(n_1849),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1866),
.B(n_1880),
.Y(n_1908)
);

CKINVDCx16_ASAP7_75t_R g1909 ( 
.A(n_1861),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1880),
.B(n_1837),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1860),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1896),
.B(n_1852),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1861),
.B(n_1801),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1865),
.B(n_1840),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1863),
.B(n_1852),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1900),
.B(n_1852),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1877),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1871),
.B(n_1810),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1863),
.B(n_1825),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_R g1920 ( 
.A(n_1876),
.B(n_1810),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1865),
.B(n_1840),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1890),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1860),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1863),
.B(n_1825),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1876),
.B(n_1836),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1871),
.B(n_1836),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1877),
.B(n_1825),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1890),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1879),
.B(n_1854),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1879),
.B(n_1830),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1884),
.B(n_1820),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1864),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1864),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1867),
.B(n_1830),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1884),
.B(n_1820),
.Y(n_1935)
);

NAND5xp2_ASAP7_75t_L g1936 ( 
.A(n_1884),
.B(n_1796),
.C(n_1805),
.D(n_1801),
.E(n_1771),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1867),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1869),
.B(n_1830),
.Y(n_1938)
);

NOR3xp33_ASAP7_75t_L g1939 ( 
.A(n_1878),
.B(n_1790),
.C(n_1796),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1885),
.B(n_1820),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1869),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1885),
.B(n_1901),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1885),
.B(n_1853),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1883),
.B(n_1859),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1870),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1870),
.B(n_1831),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1920),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1909),
.A2(n_1778),
.B(n_1715),
.Y(n_1948)
);

XOR2xp5_ASAP7_75t_L g1949 ( 
.A(n_1909),
.B(n_1817),
.Y(n_1949)
);

O2A1O1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1904),
.A2(n_1739),
.B(n_1778),
.C(n_1790),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1913),
.B(n_1939),
.Y(n_1951)
);

AO21x1_ASAP7_75t_L g1952 ( 
.A1(n_1925),
.A2(n_1897),
.B(n_1894),
.Y(n_1952)
);

CKINVDCx16_ASAP7_75t_R g1953 ( 
.A(n_1913),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1937),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1903),
.A2(n_1783),
.B1(n_1778),
.B2(n_1772),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1902),
.B(n_1900),
.Y(n_1956)
);

OAI32xp33_ASAP7_75t_L g1957 ( 
.A1(n_1908),
.A2(n_1728),
.A3(n_1883),
.B1(n_1893),
.B2(n_1850),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1903),
.B(n_1853),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1911),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1902),
.B(n_1900),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1907),
.Y(n_1961)
);

NAND4xp25_ASAP7_75t_L g1962 ( 
.A(n_1936),
.B(n_1908),
.C(n_1905),
.D(n_1917),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1907),
.B(n_1900),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1936),
.A2(n_1780),
.B1(n_1778),
.B2(n_1735),
.Y(n_1964)
);

AOI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1905),
.A2(n_1778),
.B1(n_1900),
.B2(n_1729),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1912),
.Y(n_1966)
);

OAI222xp33_ASAP7_75t_L g1967 ( 
.A1(n_1927),
.A2(n_1859),
.B1(n_1893),
.B2(n_1888),
.C1(n_1892),
.C2(n_1797),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1918),
.B(n_1853),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1910),
.A2(n_1772),
.B(n_1805),
.Y(n_1969)
);

INVxp67_ASAP7_75t_SL g1970 ( 
.A(n_1910),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1927),
.A2(n_1797),
.B1(n_1729),
.B2(n_1735),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1911),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1916),
.A2(n_1729),
.B1(n_1735),
.B2(n_1737),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1906),
.B(n_1854),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1912),
.Y(n_1975)
);

A2O1A1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1929),
.A2(n_1901),
.B(n_1897),
.C(n_1847),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1916),
.B(n_1901),
.Y(n_1977)
);

OAI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1926),
.A2(n_1729),
.B1(n_1735),
.B2(n_1728),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1906),
.B(n_1758),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1923),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1923),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1932),
.A2(n_1799),
.B(n_1897),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1934),
.B(n_1882),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1951),
.A2(n_1774),
.B(n_1915),
.C(n_1944),
.Y(n_1984)
);

OAI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1953),
.A2(n_1916),
.B1(n_1930),
.B2(n_1926),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1962),
.A2(n_1915),
.B1(n_1941),
.B2(n_1945),
.C(n_1933),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1959),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1949),
.A2(n_1964),
.B1(n_1955),
.B2(n_1958),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1959),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1967),
.A2(n_1933),
.B1(n_1941),
.B2(n_1945),
.C(n_1932),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1947),
.B(n_1916),
.Y(n_1991)
);

NOR2x1_ASAP7_75t_L g1992 ( 
.A(n_1949),
.B(n_1897),
.Y(n_1992)
);

AOI222xp33_ASAP7_75t_L g1993 ( 
.A1(n_1970),
.A2(n_1759),
.B1(n_1914),
.B2(n_1921),
.C1(n_1946),
.C2(n_1934),
.Y(n_1993)
);

XOR2x2_ASAP7_75t_L g1994 ( 
.A(n_1969),
.B(n_1715),
.Y(n_1994)
);

OAI22xp33_ASAP7_75t_SL g1995 ( 
.A1(n_1966),
.A2(n_1946),
.B1(n_1938),
.B2(n_1944),
.Y(n_1995)
);

AOI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1950),
.A2(n_1921),
.B(n_1914),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1954),
.B(n_1943),
.Y(n_1997)
);

OAI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1965),
.A2(n_1938),
.B1(n_1930),
.B2(n_1735),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1954),
.B(n_1943),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1948),
.A2(n_1942),
.B1(n_1924),
.B2(n_1919),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1948),
.A2(n_1942),
.B1(n_1924),
.B2(n_1919),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1952),
.A2(n_1735),
.B1(n_1729),
.B2(n_1740),
.Y(n_2002)
);

INVx2_ASAP7_75t_SL g2003 ( 
.A(n_1961),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1977),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1972),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1952),
.A2(n_1735),
.B1(n_1729),
.B2(n_1740),
.Y(n_2006)
);

NAND3x2_ASAP7_75t_L g2007 ( 
.A(n_1956),
.B(n_1940),
.C(n_1935),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1982),
.A2(n_1897),
.B(n_1888),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1971),
.A2(n_1735),
.B1(n_1740),
.B2(n_1737),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1974),
.B(n_1940),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_2003),
.B(n_1961),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1987),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1989),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2005),
.Y(n_2014)
);

OAI21xp33_ASAP7_75t_L g2015 ( 
.A1(n_1986),
.A2(n_1976),
.B(n_1975),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1991),
.B(n_1975),
.Y(n_2016)
);

OAI21xp33_ASAP7_75t_SL g2017 ( 
.A1(n_1992),
.A2(n_1977),
.B(n_1956),
.Y(n_2017)
);

AOI221xp5_ASAP7_75t_L g2018 ( 
.A1(n_1988),
.A2(n_1957),
.B1(n_1978),
.B2(n_1972),
.C(n_1981),
.Y(n_2018)
);

NAND2x1_ASAP7_75t_L g2019 ( 
.A(n_2002),
.B(n_1980),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_SL g2020 ( 
.A(n_1984),
.B(n_1957),
.C(n_1980),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_2004),
.B(n_1960),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1997),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2008),
.B(n_1960),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_2008),
.B(n_1963),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1999),
.Y(n_2025)
);

INVx1_ASAP7_75t_SL g2026 ( 
.A(n_1994),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1995),
.Y(n_2027)
);

INVxp67_ASAP7_75t_L g2028 ( 
.A(n_1985),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1996),
.B(n_1968),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_2010),
.Y(n_2030)
);

INVx3_ASAP7_75t_SL g2031 ( 
.A(n_2011),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2019),
.A2(n_1990),
.B(n_2001),
.Y(n_2032)
);

NAND4xp25_ASAP7_75t_L g2033 ( 
.A(n_2026),
.B(n_2006),
.C(n_2000),
.D(n_1993),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2011),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_2011),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2019),
.A2(n_1993),
.B(n_1998),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2016),
.B(n_1963),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_2028),
.B(n_1979),
.Y(n_2038)
);

O2A1O1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_2027),
.A2(n_1981),
.B(n_1973),
.C(n_1983),
.Y(n_2039)
);

OAI221xp5_ASAP7_75t_SL g2040 ( 
.A1(n_2015),
.A2(n_2009),
.B1(n_2007),
.B2(n_1983),
.C(n_1935),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2021),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_2027),
.B(n_2025),
.Y(n_2042)
);

NAND4xp25_ASAP7_75t_SL g2043 ( 
.A(n_2032),
.B(n_2018),
.C(n_2017),
.D(n_2024),
.Y(n_2043)
);

OAI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2033),
.A2(n_2020),
.B1(n_2029),
.B2(n_2022),
.C(n_2030),
.Y(n_2044)
);

NAND2xp33_ASAP7_75t_R g2045 ( 
.A(n_2042),
.B(n_2016),
.Y(n_2045)
);

NAND4xp25_ASAP7_75t_L g2046 ( 
.A(n_2038),
.B(n_2025),
.C(n_2013),
.D(n_2023),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_2036),
.A2(n_2021),
.B(n_2014),
.Y(n_2047)
);

NAND5xp2_ASAP7_75t_L g2048 ( 
.A(n_2039),
.B(n_2024),
.C(n_2023),
.D(n_2014),
.E(n_2012),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_R g2049 ( 
.A(n_2031),
.B(n_2035),
.Y(n_2049)
);

AOI221xp5_ASAP7_75t_L g2050 ( 
.A1(n_2040),
.A2(n_2012),
.B1(n_2021),
.B2(n_1922),
.C(n_1928),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2037),
.A2(n_1931),
.B1(n_1888),
.B2(n_1892),
.Y(n_2051)
);

XNOR2xp5_ASAP7_75t_L g2052 ( 
.A(n_2041),
.B(n_1731),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2034),
.A2(n_1843),
.B1(n_1931),
.B2(n_1894),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2034),
.Y(n_2054)
);

NAND2xp33_ASAP7_75t_R g2055 ( 
.A(n_2049),
.B(n_1777),
.Y(n_2055)
);

AOI221xp5_ASAP7_75t_L g2056 ( 
.A1(n_2043),
.A2(n_1928),
.B1(n_1922),
.B2(n_1892),
.C(n_1899),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2044),
.A2(n_1786),
.B1(n_1894),
.B2(n_1928),
.Y(n_2057)
);

AOI21xp33_ASAP7_75t_L g2058 ( 
.A1(n_2045),
.A2(n_1922),
.B(n_1847),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_2047),
.B(n_2050),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2052),
.A2(n_1843),
.B1(n_1894),
.B2(n_1850),
.Y(n_2060)
);

NAND4xp25_ASAP7_75t_SL g2061 ( 
.A(n_2057),
.B(n_2054),
.C(n_2048),
.D(n_2051),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_L g2062 ( 
.A(n_2059),
.B(n_2046),
.C(n_2053),
.Y(n_2062)
);

NOR3xp33_ASAP7_75t_L g2063 ( 
.A(n_2060),
.B(n_1857),
.C(n_1862),
.Y(n_2063)
);

NOR3x2_ASAP7_75t_L g2064 ( 
.A(n_2055),
.B(n_1882),
.C(n_1857),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2056),
.B(n_1872),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_2058),
.A2(n_1894),
.B(n_1862),
.Y(n_2066)
);

NAND2x1p5_ASAP7_75t_SL g2067 ( 
.A(n_2059),
.B(n_1740),
.Y(n_2067)
);

NAND4xp75_ASAP7_75t_L g2068 ( 
.A(n_2065),
.B(n_1858),
.C(n_1898),
.D(n_1873),
.Y(n_2068)
);

AOI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_2061),
.A2(n_1862),
.B1(n_1895),
.B2(n_1891),
.Y(n_2069)
);

NOR3xp33_ASAP7_75t_L g2070 ( 
.A(n_2062),
.B(n_1839),
.C(n_1841),
.Y(n_2070)
);

AND4x1_ASAP7_75t_L g2071 ( 
.A(n_2063),
.B(n_1858),
.C(n_1734),
.D(n_1833),
.Y(n_2071)
);

NAND3xp33_ASAP7_75t_SL g2072 ( 
.A(n_2066),
.B(n_1842),
.C(n_1818),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2064),
.A2(n_1862),
.B1(n_1895),
.B2(n_1891),
.Y(n_2073)
);

OAI22x1_ASAP7_75t_L g2074 ( 
.A1(n_2069),
.A2(n_2067),
.B1(n_1887),
.B2(n_1895),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2068),
.Y(n_2075)
);

AOI311xp33_ASAP7_75t_L g2076 ( 
.A1(n_2070),
.A2(n_1899),
.A3(n_1898),
.B(n_1874),
.C(n_1872),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_2072),
.A2(n_2073),
.B(n_2071),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2075),
.B(n_1882),
.Y(n_2078)
);

NOR2xp67_ASAP7_75t_L g2079 ( 
.A(n_2078),
.B(n_2077),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2079),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2079),
.A2(n_2074),
.B1(n_2076),
.B2(n_1891),
.Y(n_2081)
);

AOI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2080),
.A2(n_1890),
.B1(n_1874),
.B2(n_1889),
.Y(n_2082)
);

NAND3xp33_ASAP7_75t_L g2083 ( 
.A(n_2081),
.B(n_1881),
.C(n_1889),
.Y(n_2083)
);

INVxp67_ASAP7_75t_SL g2084 ( 
.A(n_2083),
.Y(n_2084)
);

AOI221xp5_ASAP7_75t_L g2085 ( 
.A1(n_2082),
.A2(n_1886),
.B1(n_1881),
.B2(n_1875),
.C(n_1873),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2084),
.A2(n_1887),
.B1(n_1890),
.B2(n_1875),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_2086),
.A2(n_2085),
.B1(n_1887),
.B2(n_1890),
.Y(n_2087)
);

AOI211xp5_ASAP7_75t_L g2088 ( 
.A1(n_2087),
.A2(n_1886),
.B(n_1839),
.C(n_1841),
.Y(n_2088)
);


endmodule