module real_jpeg_15667_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_306),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_0),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_3),
.B(n_49),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

NAND2x1_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_3),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_138),
.Y(n_137)
);

NAND2x1_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_4),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_4),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_4),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_4),
.B(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_5),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_5),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_5),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_5),
.B(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_8),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_9),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_10),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_10),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_10),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_10),
.B(n_187),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g129 ( 
.A(n_12),
.Y(n_129)
);

BUFx8_ASAP7_75t_L g187 ( 
.A(n_13),
.Y(n_187)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_13),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_273),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_234),
.B(n_267),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_200),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_163),
.B(n_199),
.Y(n_20)
);

AOI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_115),
.B(n_162),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_23),
.B(n_76),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.C(n_62),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_25),
.Y(n_153)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_26),
.A2(n_38),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_27),
.A2(n_28),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_41),
.B(n_43),
.Y(n_40)
);

NAND2x1p5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_41),
.Y(n_43)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_31),
.Y(n_142)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_32),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_32),
.Y(n_144)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_R g136 ( 
.A1(n_38),
.A2(n_137),
.B(n_139),
.C(n_145),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_38),
.B(n_137),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_38),
.A2(n_44),
.B1(n_137),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_40),
.A2(n_45),
.B1(n_86),
.B2(n_87),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_41),
.A2(n_126),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_41),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_41),
.B(n_140),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_41),
.A2(n_132),
.B1(n_140),
.B2(n_143),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_41),
.A2(n_140),
.B(n_242),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_43),
.B(n_81),
.C(n_87),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_46),
.A2(n_62),
.B1(n_63),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_52),
.C(n_57),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_47),
.A2(n_48),
.B1(n_57),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_47),
.A2(n_48),
.B1(n_175),
.B2(n_179),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_48),
.B(n_212),
.Y(n_211)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_48),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_48),
.B(n_64),
.C(n_175),
.Y(n_287)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_53),
.B1(n_94),
.B2(n_104),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_52),
.A2(n_53),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_53),
.A2(n_96),
.B(n_98),
.C(n_145),
.Y(n_170)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_56),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_57),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_57),
.A2(n_81),
.B1(n_89),
.B2(n_123),
.Y(n_208)
);

XNOR2x2_ASAP7_75t_L g296 ( 
.A(n_57),
.B(n_297),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_112),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_58),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_75),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_64),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_69),
.C(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_69),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_69),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_69),
.B(n_259),
.C(n_262),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_69),
.B(n_222),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_71),
.Y(n_196)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_72),
.A2(n_108),
.B1(n_174),
.B2(n_180),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_75),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_92),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_90),
.B2(n_91),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_79),
.B(n_90),
.C(n_92),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_89),
.B(n_123),
.C(n_207),
.Y(n_255)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_105),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_93),
.B(n_106),
.C(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_103),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_95),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_152),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_95),
.B(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_96),
.B(n_137),
.C(n_186),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_97),
.Y(n_260)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g297 ( 
.A1(n_98),
.A2(n_103),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_108),
.B(n_140),
.C(n_175),
.Y(n_231)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_111),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_111),
.A2(n_114),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_111),
.B(n_223),
.C(n_226),
.Y(n_262)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_114),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_125),
.B(n_126),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_134),
.B(n_161),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.C(n_130),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_130),
.B1(n_131),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_149),
.B(n_160),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_146),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_137),
.A2(n_158),
.B1(n_211),
.B2(n_216),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_137),
.B(n_213),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_143),
.B1(n_175),
.B2(n_179),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_156),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_155),
.B(n_159),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_158),
.B(n_212),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_165),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_181),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_168),
.C(n_181),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_173),
.C(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_172),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_198),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_189),
.C(n_198),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B(n_197),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_194),
.Y(n_197)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_201),
.B(n_202),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_219),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_203),
.B(n_220),
.C(n_233),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_217),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_209),
.C(n_217),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_233),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_231),
.C(n_232),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_266),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_266),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_238),
.C(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_253),
.Y(n_237)
);

XOR2x2_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_251),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_247),
.B2(n_248),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_248),
.C(n_251),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_253),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_263),
.B2(n_264),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_264),
.C(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_259),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_304),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NAND2x1p5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_278),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_293),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_290),
.B2(n_291),
.Y(n_283)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

XOR2x1_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_302),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);


endmodule