module fake_netlist_1_11650_n_48 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_48);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_48;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
BUFx6f_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_10), .B(n_4), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_1), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_6), .A2(n_14), .B1(n_2), .B2(n_1), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_17), .B(n_2), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_19), .B(n_3), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_18), .B(n_20), .Y(n_25) );
OA21x2_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_18), .B(n_20), .Y(n_26) );
INVx2_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_26), .B1(n_22), .B2(n_24), .Y(n_30) );
CKINVDCx14_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
OAI221xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_26), .B1(n_16), .B2(n_15), .C(n_8), .Y(n_32) );
XNOR2x1_ASAP7_75t_L g33 ( .A(n_31), .B(n_26), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_30), .A2(n_16), .B1(n_15), .B2(n_7), .Y(n_34) );
NAND2xp33_ASAP7_75t_R g35 ( .A(n_32), .B(n_3), .Y(n_35) );
AOI21xp5_ASAP7_75t_L g36 ( .A1(n_32), .A2(n_16), .B(n_15), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_33), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_37) );
AOI21xp33_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_5), .B(n_9), .Y(n_38) );
NOR2xp33_ASAP7_75t_R g39 ( .A(n_36), .B(n_11), .Y(n_39) );
INVx2_ASAP7_75t_L g40 ( .A(n_34), .Y(n_40) );
INVxp67_ASAP7_75t_L g41 ( .A(n_33), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g42 ( .A(n_37), .Y(n_42) );
AO22x2_ASAP7_75t_L g43 ( .A1(n_41), .A2(n_12), .B1(n_13), .B2(n_40), .Y(n_43) );
HB1xp67_ASAP7_75t_L g44 ( .A(n_39), .Y(n_44) );
INVx1_ASAP7_75t_L g45 ( .A(n_38), .Y(n_45) );
AOI21xp5_ASAP7_75t_L g46 ( .A1(n_44), .A2(n_43), .B(n_45), .Y(n_46) );
AOI21xp5_ASAP7_75t_L g47 ( .A1(n_44), .A2(n_43), .B(n_42), .Y(n_47) );
AOI21xp5_ASAP7_75t_L g48 ( .A1(n_46), .A2(n_43), .B(n_47), .Y(n_48) );
endmodule