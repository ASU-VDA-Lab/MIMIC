module fake_netlist_6_4359_n_1118 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1118);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1118;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_1015;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_842;
wire n_758;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_989;
wire n_843;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_940;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_981;
wire n_476;
wire n_880;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_71),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_17),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_37),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_42),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_78),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_180),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_56),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_126),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_183),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_124),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_25),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_59),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_55),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_67),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_18),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_63),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_104),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_140),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_110),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_203),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_201),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_107),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_66),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_154),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_9),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_88),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_6),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_72),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_3),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_174),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_48),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_127),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_150),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_64),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_38),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_155),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_45),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_32),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_204),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_161),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_165),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_12),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_208),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_192),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_53),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_132),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_156),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_102),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_31),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_70),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_177),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_24),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_120),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_46),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_233),
.Y(n_283)
);

INVxp33_ASAP7_75t_SL g284 ( 
.A(n_277),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_216),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_213),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_266),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_216),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_217),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_276),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_215),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_218),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_219),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_256),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_229),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_251),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_220),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_256),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_269),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_221),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_287),
.A2(n_225),
.B1(n_232),
.B2(n_236),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_292),
.A2(n_282),
.B1(n_281),
.B2(n_279),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_310),
.B(n_272),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_315),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_222),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_292),
.A2(n_249),
.B1(n_268),
.B2(n_265),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

CKINVDCx8_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_327),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_284),
.A2(n_271),
.B1(n_263),
.B2(n_261),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_290),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_318),
.B(n_223),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_291),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_293),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_228),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_287),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_322),
.B(n_230),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_325),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_298),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_305),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_306),
.B(n_231),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_227),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_294),
.B(n_243),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_311),
.Y(n_372)
);

OAI22x1_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_260),
.B1(n_259),
.B2(n_258),
.Y(n_373)
);

CKINVDCx8_ASAP7_75t_R g374 ( 
.A(n_307),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_255),
.Y(n_375)
);

INVx5_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

CKINVDCx6p67_ASAP7_75t_R g377 ( 
.A(n_294),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_326),
.B(n_244),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_319),
.Y(n_379)
);

OAI22x1_ASAP7_75t_SL g380 ( 
.A1(n_283),
.A2(n_252),
.B1(n_247),
.B2(n_246),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_245),
.Y(n_381)
);

BUFx12f_ASAP7_75t_L g382 ( 
.A(n_302),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_332),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_284),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_379),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_34),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_374),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_354),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_352),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_382),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_320),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_342),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_362),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_362),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_360),
.Y(n_402)
);

CKINVDCx6p67_ASAP7_75t_R g403 ( 
.A(n_377),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_360),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_357),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_357),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_370),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_346),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_386),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_386),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_386),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_386),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_369),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_387),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_387),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_387),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_333),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_387),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_376),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_376),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_376),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_376),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_384),
.B(n_320),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_346),
.Y(n_429)
);

INVxp33_ASAP7_75t_SL g430 ( 
.A(n_350),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_380),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_385),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_337),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_345),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_343),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_336),
.B(n_375),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_385),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_385),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_385),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_346),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_373),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_375),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_378),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_369),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_334),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_378),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_341),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_336),
.B(n_323),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_359),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_339),
.B(n_353),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_355),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_356),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_359),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_334),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_355),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_341),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_381),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_381),
.B(n_323),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_339),
.Y(n_462)
);

INVx4_ASAP7_75t_SL g463 ( 
.A(n_406),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_417),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_391),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_SL g467 ( 
.A(n_461),
.B(n_331),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_403),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_437),
.A2(n_369),
.B1(n_227),
.B2(n_383),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_427),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_369),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_406),
.A2(n_227),
.B1(n_383),
.B2(n_364),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_415),
.B(n_368),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_415),
.A2(n_227),
.B1(n_364),
.B2(n_344),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_462),
.A2(n_227),
.B1(n_358),
.B2(n_368),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_331),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_432),
.B(n_349),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_417),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_366),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_L g490 ( 
.A(n_446),
.B(n_227),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_399),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_408),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_436),
.B(n_366),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_410),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_429),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_442),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_392),
.B(n_361),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_453),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_430),
.A2(n_367),
.B1(n_366),
.B2(n_363),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_446),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_455),
.B(n_400),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_401),
.B(n_283),
.Y(n_505)
);

BUFx6f_ASAP7_75t_SL g506 ( 
.A(n_435),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_435),
.B(n_366),
.Y(n_507)
);

NOR3xp33_ASAP7_75t_SL g508 ( 
.A(n_443),
.B(n_0),
.C(n_1),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_454),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_419),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_449),
.B(n_367),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_458),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_459),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_447),
.B(n_361),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_439),
.B(n_361),
.Y(n_517)
);

NOR3xp33_ASAP7_75t_L g518 ( 
.A(n_451),
.B(n_340),
.C(n_338),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_446),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_459),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_396),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_405),
.B(n_407),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_435),
.B(n_363),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_440),
.B(n_363),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_441),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_367),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_433),
.B(n_340),
.C(n_338),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_456),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_444),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_412),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_413),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_445),
.A2(n_367),
.B1(n_341),
.B2(n_98),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_416),
.B(n_341),
.Y(n_535)
);

NAND3x1_ASAP7_75t_L g536 ( 
.A(n_420),
.B(n_0),
.C(n_1),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_434),
.B(n_35),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_423),
.B(n_36),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

INVx4_ASAP7_75t_SL g540 ( 
.A(n_425),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_426),
.B(n_39),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_395),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_389),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_402),
.B(n_2),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_404),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_424),
.B(n_2),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_509),
.B(n_388),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_517),
.B(n_393),
.Y(n_550)
);

OR2x2_ASAP7_75t_SL g551 ( 
.A(n_530),
.B(n_397),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_466),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_509),
.A2(n_428),
.B1(n_461),
.B2(n_5),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_464),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_517),
.B(n_431),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_479),
.A2(n_476),
.B1(n_488),
.B2(n_471),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_468),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_488),
.B(n_428),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_480),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_464),
.B(n_40),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_493),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_476),
.B(n_41),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_544),
.Y(n_563)
);

OA22x2_ASAP7_75t_L g564 ( 
.A1(n_532),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_524),
.B(n_43),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_524),
.B(n_535),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_472),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_536),
.A2(n_528),
.B1(n_522),
.B2(n_518),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_481),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_482),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_476),
.B(n_44),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_485),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_512),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_493),
.B(n_47),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_531),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_512),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

NAND2x1p5_ASAP7_75t_L g578 ( 
.A(n_542),
.B(n_49),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_476),
.B(n_50),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_515),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_531),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_478),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_465),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

AO22x2_ASAP7_75t_L g585 ( 
.A1(n_528),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_492),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_494),
.Y(n_587)
);

OA22x2_ASAP7_75t_L g588 ( 
.A1(n_533),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_476),
.B(n_51),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_520),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_487),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_513),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_495),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_496),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_502),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_497),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_499),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_484),
.B(n_10),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_518),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_479),
.B(n_52),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_535),
.B(n_54),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_500),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_501),
.B(n_57),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_510),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_514),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_471),
.B(n_507),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_539),
.B(n_58),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_537),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_609)
);

OAI22x1_ASAP7_75t_SL g610 ( 
.A1(n_491),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_465),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_516),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_521),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_516),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_540),
.B(n_60),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_549),
.B(n_504),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_581),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_577),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_558),
.B(n_505),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_561),
.B(n_546),
.Y(n_620)
);

CKINVDCx10_ASAP7_75t_R g621 ( 
.A(n_613),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_566),
.B(n_543),
.Y(n_622)
);

NOR3xp33_ASAP7_75t_L g623 ( 
.A(n_558),
.B(n_467),
.C(n_547),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_548),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_566),
.B(n_543),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_591),
.B(n_546),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_560),
.A2(n_527),
.B(n_523),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_560),
.A2(n_519),
.B(n_503),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_556),
.A2(n_501),
.B1(n_525),
.B2(n_475),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_575),
.B(n_529),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_607),
.A2(n_519),
.B(n_503),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_607),
.A2(n_519),
.B(n_474),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_580),
.Y(n_633)
);

O2A1O1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_601),
.A2(n_545),
.B(n_541),
.C(n_538),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_602),
.B(n_498),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_593),
.B(n_554),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_550),
.B(n_547),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_601),
.A2(n_534),
.B(n_498),
.C(n_538),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_609),
.A2(n_604),
.B(n_586),
.C(n_584),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_582),
.B(n_526),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_581),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_587),
.Y(n_642)
);

AOI21x1_ASAP7_75t_L g643 ( 
.A1(n_562),
.A2(n_527),
.B(n_541),
.Y(n_643)
);

CKINVDCx8_ASAP7_75t_R g644 ( 
.A(n_550),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_562),
.A2(n_475),
.B(n_477),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_602),
.B(n_565),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_551),
.B(n_511),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_590),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_599),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_571),
.A2(n_519),
.B(n_486),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_SL g651 ( 
.A1(n_574),
.A2(n_477),
.B(n_508),
.C(n_490),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_565),
.A2(n_508),
.B(n_470),
.C(n_489),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_594),
.B(n_463),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_595),
.B(n_463),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_597),
.B(n_463),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_598),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_568),
.A2(n_506),
.B1(n_540),
.B2(n_489),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_606),
.B(n_540),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_571),
.A2(n_469),
.B(n_489),
.Y(n_659)
);

AOI21xp33_ASAP7_75t_L g660 ( 
.A1(n_575),
.A2(n_470),
.B(n_469),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_548),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_579),
.A2(n_469),
.B(n_486),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_579),
.A2(n_486),
.B(n_112),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_596),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_605),
.B(n_506),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_589),
.A2(n_123),
.B(n_212),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_548),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_563),
.B(n_521),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_589),
.A2(n_122),
.B(n_209),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_573),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_612),
.A2(n_121),
.B1(n_207),
.B2(n_205),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_583),
.A2(n_118),
.B(n_202),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_592),
.B(n_17),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_583),
.A2(n_119),
.B(n_200),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_567),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_614),
.A2(n_117),
.B1(n_199),
.B2(n_197),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_568),
.B(n_19),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_638),
.A2(n_611),
.B(n_583),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_623),
.A2(n_559),
.B1(n_553),
.B2(n_564),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_619),
.B(n_555),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_618),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_616),
.B(n_553),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_644),
.B(n_615),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_619),
.B(n_555),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_641),
.Y(n_685)
);

O2A1O1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_623),
.A2(n_608),
.B(n_578),
.C(n_603),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_632),
.A2(n_611),
.B(n_578),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_SL g688 ( 
.A(n_652),
.B(n_559),
.C(n_610),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_645),
.A2(n_620),
.B(n_635),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_617),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_634),
.A2(n_569),
.B(n_572),
.C(n_552),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_621),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_L g693 ( 
.A1(n_630),
.A2(n_564),
.B(n_588),
.Y(n_693)
);

AO21x1_ASAP7_75t_L g694 ( 
.A1(n_629),
.A2(n_662),
.B(n_639),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_624),
.Y(n_695)
);

A2O1A1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_646),
.A2(n_557),
.B(n_570),
.C(n_615),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_649),
.A2(n_608),
.B(n_576),
.C(n_585),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_636),
.A2(n_588),
.B1(n_585),
.B2(n_600),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_624),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_637),
.A2(n_600),
.B1(n_611),
.B2(n_21),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_626),
.B(n_19),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_647),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_649),
.B(n_622),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_635),
.A2(n_115),
.B(n_196),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_630),
.B(n_20),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_642),
.B(n_20),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_656),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_657),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_664),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_675),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_664),
.B(n_22),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_661),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_640),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_665),
.B(n_23),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_633),
.B(n_24),
.Y(n_715)
);

BUFx8_ASAP7_75t_L g716 ( 
.A(n_677),
.Y(n_716)
);

NOR2x1_ASAP7_75t_SL g717 ( 
.A(n_658),
.B(n_61),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_653),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_718)
);

AND2x2_ASAP7_75t_SL g719 ( 
.A(n_665),
.B(n_673),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_673),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_628),
.A2(n_650),
.B(n_631),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_625),
.B(n_28),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_667),
.Y(n_723)
);

O2A1O1Ixp5_ASAP7_75t_L g724 ( 
.A1(n_643),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_648),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_668),
.B(n_29),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_663),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_670),
.B(n_33),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_627),
.A2(n_210),
.B(n_65),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_667),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

OAI22x1_ASAP7_75t_L g732 ( 
.A1(n_659),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_666),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_669),
.A2(n_76),
.B(n_77),
.C(n_79),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_660),
.B(n_80),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_654),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_705),
.A2(n_671),
.B1(n_676),
.B2(n_672),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_695),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_681),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_690),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_723),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_685),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_680),
.B(n_655),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_707),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_710),
.Y(n_745)
);

BUFx4_ASAP7_75t_SL g746 ( 
.A(n_692),
.Y(n_746)
);

BUFx12f_ASAP7_75t_L g747 ( 
.A(n_702),
.Y(n_747)
);

BUFx5_ASAP7_75t_L g748 ( 
.A(n_736),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_725),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_716),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_695),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_713),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_715),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_679),
.A2(n_674),
.B1(n_651),
.B2(n_83),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_708),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_709),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_703),
.Y(n_757)
);

BUFx2_ASAP7_75t_SL g758 ( 
.A(n_695),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_716),
.Y(n_759)
);

CKINVDCx11_ASAP7_75t_R g760 ( 
.A(n_699),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_688),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_684),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_731),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_682),
.Y(n_764)
);

BUFx2_ASAP7_75t_SL g765 ( 
.A(n_699),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_730),
.Y(n_766)
);

BUFx12f_ASAP7_75t_L g767 ( 
.A(n_699),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_728),
.Y(n_768)
);

BUFx4f_ASAP7_75t_L g769 ( 
.A(n_719),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_712),
.Y(n_770)
);

BUFx4_ASAP7_75t_SL g771 ( 
.A(n_683),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_706),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_712),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_701),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_712),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_735),
.B(n_85),
.Y(n_776)
);

BUFx12f_ASAP7_75t_L g777 ( 
.A(n_683),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_724),
.Y(n_778)
);

INVx5_ASAP7_75t_L g779 ( 
.A(n_732),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_722),
.Y(n_780)
);

BUFx2_ASAP7_75t_SL g781 ( 
.A(n_714),
.Y(n_781)
);

BUFx5_ASAP7_75t_L g782 ( 
.A(n_721),
.Y(n_782)
);

BUFx8_ASAP7_75t_L g783 ( 
.A(n_711),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_691),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_694),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_689),
.B(n_86),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_726),
.Y(n_787)
);

INVx6_ASAP7_75t_L g788 ( 
.A(n_696),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_717),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_700),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_693),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_698),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_698),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_708),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_678),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_687),
.B(n_87),
.Y(n_796)
);

CKINVDCx6p67_ASAP7_75t_R g797 ( 
.A(n_720),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_793),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_766),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_SL g801 ( 
.A1(n_790),
.A2(n_769),
.B1(n_787),
.B2(n_794),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_769),
.A2(n_727),
.B1(n_697),
.B2(n_686),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_774),
.B(n_704),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_792),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_785),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_767),
.Y(n_806)
);

AO22x2_ASAP7_75t_L g807 ( 
.A1(n_785),
.A2(n_729),
.B1(n_734),
.B2(n_733),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_766),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_757),
.B(n_89),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_742),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_744),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_752),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_795),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_780),
.B(n_90),
.Y(n_814)
);

BUFx8_ASAP7_75t_L g815 ( 
.A(n_787),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_739),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_786),
.A2(n_91),
.B(n_92),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_754),
.B(n_755),
.C(n_790),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_762),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_789),
.A2(n_96),
.B(n_97),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_784),
.A2(n_99),
.B(n_100),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_797),
.A2(n_195),
.B1(n_103),
.B2(n_105),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_772),
.B(n_101),
.Y(n_823)
);

AOI221xp5_ASAP7_75t_L g824 ( 
.A1(n_755),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.C(n_114),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_754),
.A2(n_125),
.B(n_128),
.C(n_130),
.Y(n_825)
);

AOI221xp5_ASAP7_75t_L g826 ( 
.A1(n_798),
.A2(n_787),
.B1(n_737),
.B2(n_768),
.C(n_753),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_779),
.B(n_131),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_787),
.A2(n_194),
.B1(n_135),
.B2(n_136),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_R g830 ( 
.A(n_760),
.B(n_134),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_745),
.Y(n_831)
);

AOI221xp5_ASAP7_75t_L g832 ( 
.A1(n_737),
.A2(n_137),
.B1(n_139),
.B2(n_141),
.C(n_142),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_749),
.Y(n_833)
);

AO21x2_ASAP7_75t_L g834 ( 
.A1(n_778),
.A2(n_796),
.B(n_782),
.Y(n_834)
);

BUFx2_ASAP7_75t_SL g835 ( 
.A(n_750),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_776),
.A2(n_143),
.B(n_144),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_741),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_748),
.Y(n_838)
);

AO21x2_ASAP7_75t_L g839 ( 
.A1(n_796),
.A2(n_782),
.B(n_743),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_742),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_748),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_746),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_776),
.A2(n_145),
.B(n_147),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_780),
.A2(n_193),
.B1(n_151),
.B2(n_152),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_748),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_747),
.B(n_148),
.Y(n_846)
);

AO21x2_ASAP7_75t_L g847 ( 
.A1(n_782),
.A2(n_157),
.B(n_158),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_748),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_760),
.Y(n_849)
);

INVx5_ASAP7_75t_L g850 ( 
.A(n_788),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_791),
.A2(n_160),
.B(n_162),
.Y(n_851)
);

AO31x2_ASAP7_75t_L g852 ( 
.A1(n_782),
.A2(n_163),
.A3(n_164),
.B(n_166),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_799),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_799),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_815),
.Y(n_855)
);

AOI21x1_ASAP7_75t_L g856 ( 
.A1(n_802),
.A2(n_763),
.B(n_756),
.Y(n_856)
);

AND2x6_ASAP7_75t_L g857 ( 
.A(n_827),
.B(n_780),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_800),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_813),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_813),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_840),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_808),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_805),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_811),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_839),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_841),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_805),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_841),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_838),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_845),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_848),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_815),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_834),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_833),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_804),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_812),
.B(n_780),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_804),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_816),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_837),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_831),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_850),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_834),
.Y(n_882)
);

BUFx4f_ASAP7_75t_SL g883 ( 
.A(n_849),
.Y(n_883)
);

CKINVDCx11_ASAP7_75t_R g884 ( 
.A(n_849),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_839),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_810),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_852),
.Y(n_887)
);

CKINVDCx8_ASAP7_75t_R g888 ( 
.A(n_835),
.Y(n_888)
);

NAND2x1p5_ASAP7_75t_L g889 ( 
.A(n_850),
.B(n_779),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_852),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_852),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_852),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_818),
.A2(n_781),
.B1(n_788),
.B2(n_762),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_826),
.A2(n_764),
.B1(n_761),
.B2(n_777),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_817),
.A2(n_782),
.B(n_738),
.Y(n_895)
);

AO21x2_ASAP7_75t_L g896 ( 
.A1(n_825),
.A2(n_803),
.B(n_851),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_842),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_864),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_893),
.A2(n_824),
.B1(n_788),
.B2(n_801),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_894),
.A2(n_801),
.B1(n_832),
.B2(n_819),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_859),
.B(n_740),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_889),
.B(n_828),
.Y(n_902)
);

BUFx4f_ASAP7_75t_L g903 ( 
.A(n_897),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_889),
.B(n_828),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_SL g905 ( 
.A(n_876),
.B(n_759),
.C(n_825),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_884),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_864),
.Y(n_907)
);

NAND4xp25_ASAP7_75t_L g908 ( 
.A(n_894),
.B(n_823),
.C(n_741),
.D(n_822),
.Y(n_908)
);

AO31x2_ASAP7_75t_L g909 ( 
.A1(n_887),
.A2(n_807),
.A3(n_779),
.B(n_751),
.Y(n_909)
);

OR2x4_ASAP7_75t_L g910 ( 
.A(n_883),
.B(n_814),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_896),
.A2(n_822),
.B1(n_807),
.B2(n_783),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_874),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_860),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_879),
.B(n_748),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_861),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_865),
.A2(n_820),
.B(n_821),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_SL g917 ( 
.A(n_890),
.B(n_746),
.C(n_771),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_SL g918 ( 
.A(n_855),
.B(n_830),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_896),
.A2(n_807),
.B1(n_783),
.B2(n_850),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_878),
.B(n_850),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_863),
.B(n_867),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_874),
.B(n_806),
.Y(n_922)
);

NAND3xp33_ASAP7_75t_SL g923 ( 
.A(n_888),
.B(n_830),
.C(n_844),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_888),
.A2(n_779),
.B1(n_844),
.B2(n_829),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_886),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_878),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_R g927 ( 
.A(n_897),
.B(n_750),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_SL g928 ( 
.A(n_890),
.B(n_771),
.C(n_761),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_898),
.B(n_865),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_909),
.B(n_873),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_921),
.B(n_853),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_926),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_921),
.B(n_882),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_907),
.B(n_885),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_912),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_923),
.A2(n_896),
.B1(n_829),
.B2(n_857),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_909),
.B(n_873),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_909),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_922),
.B(n_873),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_920),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_906),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_914),
.B(n_882),
.Y(n_942)
);

NOR2xp67_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_873),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_916),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_916),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_919),
.B(n_868),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_901),
.B(n_853),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_915),
.B(n_855),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_925),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_911),
.B(n_866),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_902),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_945),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_951),
.B(n_902),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_936),
.A2(n_900),
.B1(n_905),
.B2(n_924),
.Y(n_954)
);

BUFx4f_ASAP7_75t_L g955 ( 
.A(n_949),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_932),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_950),
.A2(n_908),
.B1(n_899),
.B2(n_918),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_950),
.A2(n_951),
.B1(n_946),
.B2(n_949),
.Y(n_958)
);

OAI221xp5_ASAP7_75t_L g959 ( 
.A1(n_948),
.A2(n_903),
.B1(n_917),
.B2(n_928),
.C(n_872),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_932),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_935),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_951),
.Y(n_962)
);

OAI221xp5_ASAP7_75t_L g963 ( 
.A1(n_940),
.A2(n_903),
.B1(n_902),
.B2(n_904),
.C(n_872),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_947),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_950),
.A2(n_856),
.B(n_904),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_934),
.B(n_854),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_954),
.A2(n_946),
.B1(n_904),
.B2(n_940),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_957),
.A2(n_946),
.B1(n_940),
.B2(n_941),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_956),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_962),
.B(n_939),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_961),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_953),
.B(n_939),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_955),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_960),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_L g975 ( 
.A1(n_958),
.A2(n_947),
.B(n_931),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_953),
.B(n_939),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_955),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_969),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_972),
.B(n_976),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_977),
.B(n_952),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_969),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_977),
.B(n_965),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_972),
.B(n_964),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_968),
.B(n_966),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_984),
.B(n_975),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_978),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_981),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_979),
.B(n_977),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_983),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_983),
.B(n_974),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_980),
.B(n_967),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_L g992 ( 
.A1(n_985),
.A2(n_982),
.B1(n_980),
.B2(n_973),
.C(n_945),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_988),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_989),
.B(n_980),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_991),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_990),
.B(n_973),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_986),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_987),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_989),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_989),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_988),
.B(n_973),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_988),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_1002),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_1002),
.B(n_976),
.Y(n_1006)
);

OR2x2_ASAP7_75t_L g1007 ( 
.A(n_995),
.B(n_982),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_1002),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_995),
.B(n_971),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_998),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_994),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1005),
.B(n_993),
.Y(n_1012)
);

CKINVDCx14_ASAP7_75t_R g1013 ( 
.A(n_1008),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1003),
.A2(n_993),
.B1(n_996),
.B2(n_992),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_1007),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_1004),
.A2(n_997),
.B(n_1000),
.C(n_999),
.Y(n_1016)
);

OAI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_1011),
.A2(n_963),
.B1(n_959),
.B2(n_982),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1010),
.B(n_1001),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_1009),
.A2(n_941),
.B(n_959),
.Y(n_1019)
);

OAI22xp33_ASAP7_75t_SL g1020 ( 
.A1(n_1009),
.A2(n_941),
.B1(n_945),
.B2(n_971),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_1015),
.B(n_1006),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1012),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1016),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1018),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1014),
.B(n_970),
.Y(n_1026)
);

AND4x1_ASAP7_75t_L g1027 ( 
.A(n_1019),
.B(n_927),
.C(n_809),
.D(n_970),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_1020),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1017),
.B(n_966),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_1022),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_1021),
.B(n_931),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1028),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1024),
.B(n_945),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1026),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_1025),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1023),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1026),
.B(n_935),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1027),
.B(n_942),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_1029),
.B(n_806),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_1030),
.B(n_910),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1032),
.B(n_944),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_1039),
.B(n_770),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1031),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_1039),
.B(n_944),
.Y(n_1044)
);

AND3x1_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_944),
.C(n_937),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_1035),
.B(n_943),
.Y(n_1046)
);

AOI211xp5_ASAP7_75t_SL g1047 ( 
.A1(n_1033),
.A2(n_846),
.B(n_943),
.C(n_937),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1040),
.B(n_1036),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1043),
.A2(n_1038),
.B1(n_1037),
.B2(n_942),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1041),
.B(n_935),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_1046),
.A2(n_847),
.B(n_889),
.C(n_775),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_1042),
.B(n_751),
.C(n_770),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_1044),
.B(n_167),
.Y(n_1053)
);

AOI221xp5_ASAP7_75t_L g1054 ( 
.A1(n_1045),
.A2(n_942),
.B1(n_930),
.B2(n_934),
.C(n_933),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1048),
.A2(n_1047),
.B1(n_930),
.B2(n_938),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_SL g1056 ( 
.A(n_1050),
.B(n_168),
.C(n_169),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1049),
.B(n_942),
.Y(n_1057)
);

OAI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1052),
.A2(n_938),
.B1(n_881),
.B2(n_937),
.Y(n_1058)
);

AOI211xp5_ASAP7_75t_L g1059 ( 
.A1(n_1053),
.A2(n_836),
.B(n_843),
.C(n_773),
.Y(n_1059)
);

OAI211xp5_ASAP7_75t_L g1060 ( 
.A1(n_1051),
.A2(n_773),
.B(n_856),
.C(n_770),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_SL g1061 ( 
.A1(n_1054),
.A2(n_847),
.B(n_881),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1048),
.A2(n_881),
.B(n_938),
.C(n_930),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1048),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1049),
.B(n_934),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1056),
.B(n_1063),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1064),
.B(n_930),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1058),
.A2(n_930),
.B1(n_765),
.B2(n_758),
.C(n_933),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1057),
.B(n_1055),
.Y(n_1068)
);

AOI221xp5_ASAP7_75t_L g1069 ( 
.A1(n_1061),
.A2(n_933),
.B1(n_770),
.B2(n_929),
.C(n_891),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_L g1070 ( 
.A(n_1060),
.B(n_933),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_1062),
.Y(n_1071)
);

AND3x2_ASAP7_75t_L g1072 ( 
.A(n_1059),
.B(n_929),
.C(n_171),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1063),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_1073),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1068),
.Y(n_1075)
);

NOR2x1_ASAP7_75t_L g1076 ( 
.A(n_1065),
.B(n_764),
.Y(n_1076)
);

AND3x2_ASAP7_75t_L g1077 ( 
.A(n_1069),
.B(n_170),
.C(n_172),
.Y(n_1077)
);

NAND3x1_ASAP7_75t_L g1078 ( 
.A(n_1070),
.B(n_929),
.C(n_891),
.Y(n_1078)
);

NAND4xp75_ASAP7_75t_L g1079 ( 
.A(n_1067),
.B(n_173),
.C(n_175),
.D(n_176),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1071),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_1066),
.Y(n_1081)
);

NAND3x1_ASAP7_75t_L g1082 ( 
.A(n_1072),
.B(n_867),
.C(n_863),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_1073),
.B(n_880),
.C(n_871),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1073),
.B(n_880),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1073),
.A2(n_854),
.B1(n_892),
.B2(n_887),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_SL g1086 ( 
.A(n_1073),
.B(n_178),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1076),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1075),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_1074),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1080),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1082),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_1081),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1086),
.B(n_179),
.Y(n_1093)
);

XOR2xp5_ASAP7_75t_L g1094 ( 
.A(n_1079),
.B(n_181),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1078),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_1091),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1088),
.A2(n_1084),
.B1(n_1077),
.B2(n_1083),
.Y(n_1097)
);

AND3x1_ASAP7_75t_L g1098 ( 
.A(n_1090),
.B(n_1085),
.C(n_185),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1092),
.A2(n_857),
.B1(n_869),
.B2(n_871),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_1089),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1087),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1095),
.Y(n_1102)
);

OAI322xp33_ASAP7_75t_L g1103 ( 
.A1(n_1101),
.A2(n_1094),
.A3(n_1093),
.B1(n_892),
.B2(n_869),
.C1(n_870),
.C2(n_190),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1100),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1098),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1104),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_1106),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1107),
.Y(n_1108)
);

OAI322xp33_ASAP7_75t_L g1109 ( 
.A1(n_1108),
.A2(n_1102),
.A3(n_1096),
.B1(n_1097),
.B2(n_1105),
.C1(n_1100),
.C2(n_1103),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1108),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1110),
.A2(n_1099),
.B1(n_875),
.B2(n_877),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1109),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1112),
.A2(n_857),
.B1(n_186),
.B2(n_187),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_R g1114 ( 
.A1(n_1111),
.A2(n_182),
.B1(n_188),
.B2(n_189),
.Y(n_1114)
);

AOI22x1_ASAP7_75t_L g1115 ( 
.A1(n_1114),
.A2(n_191),
.B1(n_862),
.B2(n_858),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1113),
.A2(n_895),
.B(n_870),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1115),
.A2(n_895),
.B(n_870),
.Y(n_1117)
);

AOI211xp5_ASAP7_75t_L g1118 ( 
.A1(n_1117),
.A2(n_1116),
.B(n_862),
.C(n_875),
.Y(n_1118)
);


endmodule