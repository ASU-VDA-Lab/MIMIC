module fake_jpeg_20395_n_111 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_SL g9 ( 
.A(n_8),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_29),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_15),
.B1(n_9),
.B2(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_38),
.B1(n_28),
.B2(n_29),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_15),
.B1(n_9),
.B2(n_14),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_25),
.A2(n_20),
.B(n_10),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_49),
.B1(n_29),
.B2(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_50),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_33),
.C(n_36),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_11),
.A3(n_10),
.B1(n_13),
.B2(n_15),
.C1(n_39),
.C2(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_49),
.B1(n_29),
.B2(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_70),
.B1(n_18),
.B2(n_1),
.Y(n_81)
);

OAI22x1_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_41),
.B1(n_44),
.B2(n_43),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_52),
.B1(n_57),
.B2(n_14),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_27),
.A3(n_47),
.B1(n_38),
.B2(n_37),
.C1(n_16),
.C2(n_12),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_23),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_47),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_52),
.Y(n_71)
);

OAI21x1_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_6),
.B(n_7),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_11),
.B(n_39),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_30),
.B1(n_31),
.B2(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_13),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_68),
.B(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_13),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_22),
.B1(n_18),
.B2(n_13),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_22),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_86),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_71),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_60),
.B1(n_78),
.B2(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_75),
.B(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_79),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_95),
.C(n_84),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_18),
.C(n_2),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_0),
.C(n_1),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_5),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_106),
.C(n_103),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_109),
.B(n_0),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_107),
.A2(n_0),
.B(n_1),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_0),
.Y(n_111)
);


endmodule