module fake_jpeg_20078_n_43 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_43);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_43;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_21),
.B1(n_19),
.B2(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_32)
);

CKINVDCx12_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_13),
.B(n_18),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.C(n_34),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_37),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_38),
.B(n_1),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_2),
.Y(n_43)
);


endmodule