module fake_jpeg_13349_n_28 (n_3, n_2, n_1, n_0, n_4, n_5, n_28);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx4f_ASAP7_75t_SL g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_8),
.A2(n_0),
.B1(n_2),
.B2(n_1),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_6),
.C(n_7),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_15),
.C(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_0),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_9),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_1),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_16),
.C(n_13),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_26),
.A2(n_20),
.B(n_22),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_26),
.B1(n_18),
.B2(n_19),
.Y(n_28)
);


endmodule