module real_jpeg_6371_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_1),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_1),
.A2(n_34),
.B1(n_72),
.B2(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_2),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_3),
.A2(n_88),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_3),
.Y(n_142)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_5),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_6),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_6),
.B(n_126),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_123),
.B1(n_170),
.B2(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_181),
.C(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_6),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_6),
.B(n_98),
.Y(n_208)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_7),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_70),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_43),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_10),
.A2(n_43),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_165),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_163),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_92),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_14),
.B(n_92),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_56),
.C(n_64),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_15),
.A2(n_16),
.B1(n_56),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_31),
.B(n_38),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_17)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_23),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_27),
.Y(n_141)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_30),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_31),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_47),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_39),
.B(n_98),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_46),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_46),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_47),
.Y(n_96)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_56),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_60),
.Y(n_162)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_64),
.B(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_76),
.B(n_83),
.Y(n_64)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_65),
.Y(n_213)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_76),
.A2(n_83),
.B(n_123),
.Y(n_199)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_77),
.B(n_86),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_77),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_136),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_105),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_96),
.A2(n_169),
.B(n_176),
.Y(n_168)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_118),
.B(n_128),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B1(n_113),
.B2(n_117),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_123),
.B(n_124),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_148),
.A3(n_149),
.B1(n_152),
.B2(n_156),
.Y(n_147)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_143),
.B(n_146),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_202),
.B(n_206),
.Y(n_201)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_188),
.B(n_219),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_185),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_168),
.A2(n_177),
.B1(n_178),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_210),
.B(n_218),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_200),
.B(n_209),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_199),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_208),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_208),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_216),
.Y(n_218)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);


endmodule