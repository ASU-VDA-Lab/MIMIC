module fake_jpeg_20590_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_31),
.Y(n_50)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_24),
.B1(n_22),
.B2(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_24),
.B1(n_32),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_22),
.B1(n_18),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_39),
.B1(n_38),
.B2(n_45),
.Y(n_96)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_25),
.CON(n_59),
.SN(n_59)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_42),
.B(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_26),
.B1(n_32),
.B2(n_16),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_39),
.B1(n_45),
.B2(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2x1_ASAP7_75t_SL g113 ( 
.A(n_66),
.B(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_72),
.B(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_84),
.C(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_42),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_96),
.B1(n_102),
.B2(n_53),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_33),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_99),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_21),
.B1(n_23),
.B2(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_100),
.B1(n_38),
.B2(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_33),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_26),
.C(n_25),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_33),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_37),
.B1(n_25),
.B2(n_32),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_33),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_105),
.CI(n_106),
.CON(n_119),
.SN(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_29),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_29),
.Y(n_106)
);

AO21x2_ASAP7_75t_SL g107 ( 
.A1(n_98),
.A2(n_38),
.B(n_41),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_102),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_45),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_135),
.C(n_89),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_124),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_44),
.B1(n_53),
.B2(n_51),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_86),
.B1(n_97),
.B2(n_91),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_96),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_37),
.C(n_35),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_113),
.B(n_72),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_138),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_76),
.B1(n_81),
.B2(n_71),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_124),
.B(n_108),
.C(n_131),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_75),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_65),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_149),
.B(n_155),
.Y(n_186)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_73),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_153),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_118),
.B(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_152),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_65),
.B1(n_88),
.B2(n_70),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_119),
.B1(n_122),
.B2(n_92),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_73),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_95),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_163),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_21),
.B(n_35),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_111),
.B1(n_16),
.B2(n_17),
.Y(n_190)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_118),
.A2(n_87),
.B(n_77),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_160),
.B(n_16),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_119),
.B(n_21),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_107),
.B(n_80),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_167),
.Y(n_182)
);

NOR2x1_ASAP7_75t_SL g165 ( 
.A(n_107),
.B(n_25),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_20),
.C(n_29),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_74),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_129),
.B1(n_107),
.B2(n_124),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_168),
.A2(n_172),
.B1(n_174),
.B2(n_189),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_170),
.B(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_180),
.B1(n_190),
.B2(n_148),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_161),
.B1(n_141),
.B2(n_144),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_124),
.B1(n_133),
.B2(n_135),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_117),
.B(n_122),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_119),
.C(n_92),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_137),
.C(n_186),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_90),
.B1(n_121),
.B2(n_85),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_111),
.B1(n_117),
.B2(n_121),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_196),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_145),
.A2(n_23),
.B(n_28),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_199),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_29),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_200),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_28),
.B1(n_23),
.B2(n_17),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_143),
.C(n_140),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_202),
.A2(n_211),
.B(n_226),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_219),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_217),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_218),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_181),
.B(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_209),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_146),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_127),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_213),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_167),
.A3(n_138),
.B1(n_149),
.B2(n_157),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_159),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_178),
.B(n_177),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_220),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_183),
.A2(n_78),
.B1(n_103),
.B2(n_20),
.Y(n_221)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_187),
.B1(n_169),
.B2(n_175),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_8),
.C(n_14),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_186),
.C(n_195),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_198),
.B1(n_171),
.B2(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_190),
.B1(n_169),
.B2(n_184),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_177),
.B(n_6),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_193),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_0),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_243),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_230),
.B1(n_226),
.B2(n_205),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_252),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_222),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_184),
.B1(n_185),
.B2(n_174),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_196),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_254),
.A2(n_236),
.B1(n_2),
.B2(n_1),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_218),
.C(n_206),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_263),
.C(n_265),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_260),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_225),
.C(n_229),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_261),
.A2(n_256),
.B1(n_168),
.B2(n_266),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_204),
.C(n_228),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_267),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_216),
.C(n_213),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_217),
.C(n_172),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_272),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_SL g270 ( 
.A(n_239),
.B(n_211),
.C(n_225),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_270),
.A2(n_247),
.B(n_224),
.Y(n_278)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_215),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_248),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_278),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_238),
.B1(n_237),
.B2(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_244),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_283),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_231),
.B(n_242),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_283),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_242),
.B(n_245),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_223),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_294),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_255),
.C(n_263),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_3),
.C(n_4),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_303),
.C(n_276),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_3),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_300),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_3),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_275),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_286),
.C(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_313),
.C(n_6),
.Y(n_318)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_311),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_309),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_301),
.B1(n_280),
.B2(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_287),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_297),
.B(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_285),
.C(n_281),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_4),
.C(n_6),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_318),
.Y(n_322)
);

OA21x2_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_310),
.B(n_312),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_8),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_7),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_10),
.B(n_11),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_315),
.Y(n_321)
);

O2A1O1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_323),
.B(n_324),
.C(n_319),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_317),
.B(n_320),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

AOI221xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_10),
.B1(n_11),
.B2(n_15),
.C(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_10),
.Y(n_331)
);


endmodule