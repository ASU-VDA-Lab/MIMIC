module fake_netlist_5_1577_n_753 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_753);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_753;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_385;
wire n_212;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_509;
wire n_568;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_344;
wire n_287;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_679;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_15),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_44),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_63),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_101),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_55),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_8),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_14),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_L g173 ( 
.A(n_76),
.B(n_10),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_72),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_54),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_1),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_24),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_69),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_73),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_102),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_68),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_117),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_66),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_65),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_98),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_2),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_108),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_104),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_67),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_11),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_123),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_27),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_9),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_86),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_154),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_92),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_131),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_129),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_38),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_20),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_41),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_150),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_64),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_20),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_137),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_50),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_25),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_5),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_94),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_113),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_87),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_40),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_0),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_14),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_19),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_16),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_120),
.B(n_139),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_103),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_89),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_84),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_51),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_4),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_159),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_177),
.A2(n_0),
.B(n_1),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

BUFx8_ASAP7_75t_SL g251 ( 
.A(n_234),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_168),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_2),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_3),
.Y(n_254)
);

BUFx8_ASAP7_75t_SL g255 ( 
.A(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_188),
.B(n_5),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g259 ( 
.A1(n_187),
.A2(n_6),
.B(n_7),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVxp33_ASAP7_75t_SL g261 ( 
.A(n_158),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_95),
.B(n_157),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_167),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_188),
.B(n_196),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_174),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_196),
.A2(n_6),
.B(n_7),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_180),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_21),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_175),
.Y(n_274)
);

OAI22x1_ASAP7_75t_SL g275 ( 
.A1(n_169),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_180),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_162),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_164),
.B(n_12),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_165),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_179),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_183),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_183),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_160),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_170),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_183),
.B(n_13),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_181),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_183),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_161),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_183),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_163),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_215),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_198),
.B(n_13),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_222),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

BUFx8_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

BUFx8_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_173),
.B(n_15),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_172),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_244),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_166),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_252),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_171),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_252),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_251),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_255),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_255),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_280),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_246),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_261),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_248),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_192),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_296),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_195),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_249),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_254),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_297),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_R g330 ( 
.A(n_267),
.B(n_225),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_298),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_248),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_298),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_270),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_270),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_247),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_247),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_266),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_274),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_241),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_279),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_279),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_299),
.B(n_203),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_294),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_253),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_349),
.Y(n_352)
);

AOI21x1_ASAP7_75t_L g353 ( 
.A1(n_338),
.A2(n_265),
.B(n_285),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_299),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_301),
.B(n_258),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_349),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_304),
.C(n_302),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_271),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_307),
.B(n_278),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

BUFx6f_ASAP7_75t_SL g362 ( 
.A(n_300),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_278),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_323),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_337),
.B(n_228),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_243),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_271),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_271),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_309),
.B(n_271),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_339),
.B(n_176),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_317),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_318),
.B(n_258),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_250),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_269),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_330),
.B(n_178),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_340),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_322),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_306),
.B(n_256),
.Y(n_386)
);

NOR3xp33_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_227),
.C(n_207),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_321),
.B(n_328),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_334),
.B(n_282),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_282),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_288),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_182),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_311),
.B(n_269),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_311),
.B(n_284),
.Y(n_395)
);

AOI221xp5_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_275),
.B1(n_233),
.B2(n_236),
.C(n_232),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_L g398 ( 
.A(n_320),
.B(n_273),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_320),
.B(n_288),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_320),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_320),
.B(n_284),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_326),
.B(n_273),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_333),
.B(n_185),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_313),
.B(n_284),
.Y(n_409)
);

OR2x6_ASAP7_75t_L g410 ( 
.A(n_310),
.B(n_257),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_308),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_312),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_314),
.B(n_286),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_315),
.B(n_286),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_300),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_345),
.B(n_286),
.Y(n_416)
);

AND2x6_ASAP7_75t_SL g417 ( 
.A(n_345),
.B(n_260),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_268),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_399),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_367),
.B(n_186),
.Y(n_420)
);

OR2x6_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_268),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_356),
.B(n_268),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_356),
.B(n_245),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_411),
.A2(n_245),
.B1(n_259),
.B2(n_189),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_386),
.A2(n_245),
.B1(n_259),
.B2(n_273),
.Y(n_426)
);

AND2x2_ASAP7_75t_SL g427 ( 
.A(n_396),
.B(n_259),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_360),
.B(n_287),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_366),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_416),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

AND2x2_ASAP7_75t_SL g434 ( 
.A(n_387),
.B(n_287),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_190),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_369),
.B(n_287),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_365),
.A2(n_398),
.B(n_394),
.C(n_415),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_370),
.B(n_382),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_414),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_385),
.B(n_263),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_377),
.B(n_291),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_377),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_291),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_414),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_291),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_407),
.A2(n_210),
.B1(n_240),
.B2(n_239),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_384),
.B(n_191),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_413),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_358),
.B(n_293),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_293),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_409),
.B(n_193),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_406),
.A2(n_273),
.B1(n_293),
.B2(n_281),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_388),
.B(n_194),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_392),
.A2(n_217),
.B1(n_199),
.B2(n_201),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_372),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_391),
.B(n_273),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_375),
.B(n_197),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_376),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_383),
.B(n_202),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_391),
.B(n_205),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_368),
.B(n_208),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_400),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_400),
.B(n_209),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_408),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_352),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_353),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_SL g474 ( 
.A(n_373),
.B(n_226),
.C(n_218),
.Y(n_474)
);

BUFx4f_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_374),
.A2(n_290),
.B1(n_281),
.B2(n_224),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_405),
.B(n_212),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

OR2x2_ASAP7_75t_SL g479 ( 
.A(n_417),
.B(n_16),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_393),
.A2(n_223),
.B(n_219),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_401),
.B(n_281),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_395),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_362),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_441),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_478),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_418),
.A2(n_359),
.B1(n_371),
.B2(n_357),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_432),
.B(n_397),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_422),
.A2(n_402),
.B(n_401),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_420),
.B(n_437),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_441),
.B(n_447),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_425),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_419),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_362),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_422),
.A2(n_290),
.B1(n_100),
.B2(n_155),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_423),
.A2(n_401),
.B(n_99),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_454),
.B(n_17),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_452),
.Y(n_501)
);

NOR2x1_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_401),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_475),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_423),
.A2(n_430),
.B(n_472),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_483),
.Y(n_505)
);

NOR2x1_ASAP7_75t_R g506 ( 
.A(n_462),
.B(n_401),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_444),
.A2(n_18),
.B(n_19),
.C(n_22),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_462),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_471),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_434),
.B(n_23),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_440),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_446),
.A2(n_107),
.B1(n_26),
.B2(n_28),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_427),
.A2(n_110),
.B1(n_29),
.B2(n_30),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_469),
.B(n_18),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_475),
.Y(n_516)
);

AOI221xp5_ASAP7_75t_L g517 ( 
.A1(n_450),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.C(n_36),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_39),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_456),
.B(n_42),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_463),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_479),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_SL g522 ( 
.A1(n_457),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g523 ( 
.A(n_474),
.B(n_52),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_456),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_464),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_468),
.B(n_53),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_473),
.A2(n_56),
.B(n_57),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_467),
.B(n_58),
.Y(n_528)
);

OAI21xp33_ASAP7_75t_L g529 ( 
.A1(n_459),
.A2(n_59),
.B(n_60),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_421),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_436),
.B(n_61),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_477),
.B(n_71),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_465),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_472),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_461),
.A2(n_75),
.B(n_77),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_466),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_SL g538 ( 
.A(n_433),
.B(n_78),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_489),
.A2(n_461),
.B(n_443),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_503),
.B(n_439),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_504),
.A2(n_445),
.B(n_443),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_499),
.A2(n_445),
.B(n_449),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_536),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_492),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_528),
.A2(n_438),
.B(n_470),
.Y(n_545)
);

AO21x2_ASAP7_75t_L g546 ( 
.A1(n_490),
.A2(n_470),
.B(n_467),
.Y(n_546)
);

CKINVDCx6p67_ASAP7_75t_R g547 ( 
.A(n_510),
.Y(n_547)
);

AO21x1_ASAP7_75t_L g548 ( 
.A1(n_526),
.A2(n_442),
.B(n_449),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_502),
.A2(n_455),
.B(n_481),
.Y(n_550)
);

BUFx5_ASAP7_75t_L g551 ( 
.A(n_530),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_509),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_518),
.A2(n_455),
.B(n_481),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_485),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_486),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_536),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_487),
.A2(n_451),
.B(n_428),
.Y(n_557)
);

NAND2x1p5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_428),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_494),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_505),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_484),
.Y(n_561)
);

AO21x2_ASAP7_75t_L g562 ( 
.A1(n_511),
.A2(n_442),
.B(n_480),
.Y(n_562)
);

BUFx2_ASAP7_75t_SL g563 ( 
.A(n_503),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_497),
.Y(n_564)
);

BUFx2_ASAP7_75t_SL g565 ( 
.A(n_516),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_515),
.A2(n_426),
.B(n_424),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_524),
.B(n_421),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_520),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_497),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_491),
.B(n_421),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_L g571 ( 
.A(n_534),
.B(n_79),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_524),
.B(n_537),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_498),
.A2(n_476),
.B(n_426),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_496),
.Y(n_575)
);

BUFx8_ASAP7_75t_L g576 ( 
.A(n_519),
.Y(n_576)
);

AO21x1_ASAP7_75t_L g577 ( 
.A1(n_532),
.A2(n_80),
.B(n_82),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_493),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_500),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_512),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_534),
.B(n_88),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_501),
.B(n_152),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_500),
.B(n_90),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_535),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_534),
.B(n_91),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_548),
.A2(n_522),
.B(n_488),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_570),
.B(n_506),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_559),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_583),
.A2(n_531),
.B1(n_514),
.B2(n_495),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_556),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_544),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_582),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_560),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_578),
.Y(n_595)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_556),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_578),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_574),
.A2(n_533),
.B(n_529),
.Y(n_598)
);

NAND2x1p5_ASAP7_75t_L g599 ( 
.A(n_543),
.B(n_538),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_570),
.B(n_508),
.Y(n_600)
);

BUFx6f_ASAP7_75t_SL g601 ( 
.A(n_564),
.Y(n_601)
);

OA21x2_ASAP7_75t_L g602 ( 
.A1(n_541),
.A2(n_507),
.B(n_517),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_552),
.A2(n_521),
.B1(n_513),
.B2(n_527),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_583),
.A2(n_508),
.B1(n_527),
.B2(n_535),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_568),
.B(n_93),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_563),
.Y(n_606)
);

CKINVDCx11_ASAP7_75t_R g607 ( 
.A(n_560),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_582),
.A2(n_566),
.B1(n_573),
.B2(n_567),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_572),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_564),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_523),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_554),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g613 ( 
.A1(n_541),
.A2(n_539),
.B(n_550),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_97),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_580),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_566),
.A2(n_105),
.B1(n_111),
.B2(n_112),
.Y(n_617)
);

AO21x2_ASAP7_75t_L g618 ( 
.A1(n_550),
.A2(n_115),
.B(n_116),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_573),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_567),
.A2(n_122),
.B1(n_124),
.B2(n_127),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_543),
.B(n_128),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_556),
.B(n_130),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_132),
.Y(n_623)
);

CKINVDCx11_ASAP7_75t_R g624 ( 
.A(n_547),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_R g625 ( 
.A(n_594),
.B(n_547),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_R g626 ( 
.A(n_607),
.B(n_569),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_590),
.A2(n_583),
.B1(n_540),
.B2(n_579),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_609),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_614),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_592),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_619),
.A2(n_585),
.B(n_581),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_SL g632 ( 
.A(n_598),
.B(n_577),
.C(n_581),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_598),
.A2(n_576),
.B1(n_567),
.B2(n_540),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_624),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_612),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_622),
.B(n_585),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_589),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_R g638 ( 
.A(n_596),
.B(n_569),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_593),
.B(n_576),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_587),
.B(n_595),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_597),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_608),
.B(n_546),
.Y(n_642)
);

AND2x2_ASAP7_75t_SL g643 ( 
.A(n_617),
.B(n_542),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_616),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_610),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_622),
.B(n_571),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_603),
.A2(n_565),
.B1(n_571),
.B2(n_558),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_623),
.B(n_611),
.Y(n_648)
);

AOI222xp33_ASAP7_75t_L g649 ( 
.A1(n_600),
.A2(n_576),
.B1(n_574),
.B2(n_549),
.C1(n_555),
.C2(n_557),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_593),
.B(n_546),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_R g651 ( 
.A(n_588),
.B(n_584),
.Y(n_651)
);

OR2x2_ASAP7_75t_SL g652 ( 
.A(n_605),
.B(n_551),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_615),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_R g654 ( 
.A(n_596),
.B(n_549),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_603),
.B(n_551),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_596),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_602),
.B(n_545),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_591),
.B(n_557),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_606),
.Y(n_659)
);

CKINVDCx8_ASAP7_75t_R g660 ( 
.A(n_622),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_602),
.B(n_545),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_R g662 ( 
.A(n_601),
.B(n_551),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_591),
.B(n_551),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_604),
.A2(n_542),
.B(n_562),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_650),
.B(n_648),
.Y(n_665)
);

AND2x2_ASAP7_75t_SL g666 ( 
.A(n_643),
.B(n_642),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_658),
.B(n_618),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_642),
.B(n_613),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_627),
.A2(n_633),
.B1(n_655),
.B2(n_636),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_640),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_657),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_652),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_644),
.B(n_613),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_661),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_637),
.B(n_627),
.Y(n_675)
);

AOI221xp5_ASAP7_75t_L g676 ( 
.A1(n_641),
.A2(n_620),
.B1(n_601),
.B2(n_586),
.C(n_618),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_635),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_630),
.B(n_586),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_636),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_645),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_649),
.B(n_621),
.Y(n_681)
);

OAI211xp5_ASAP7_75t_SL g682 ( 
.A1(n_641),
.A2(n_584),
.B(n_551),
.C(n_599),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_628),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_658),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_659),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_632),
.A2(n_647),
.B1(n_631),
.B2(n_664),
.C(n_653),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_646),
.B(n_542),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_651),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_668),
.B(n_639),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_672),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_672),
.B(n_663),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_672),
.B(n_656),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_670),
.B(n_647),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_665),
.B(n_660),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_678),
.B(n_553),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_683),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_684),
.B(n_634),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_673),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_689),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_675),
.A2(n_681),
.B1(n_669),
.B2(n_666),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_687),
.B(n_625),
.Y(n_702)
);

OAI221xp5_ASAP7_75t_SL g703 ( 
.A1(n_686),
.A2(n_626),
.B1(n_662),
.B2(n_638),
.C(n_654),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_678),
.B(n_551),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_685),
.B(n_558),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_668),
.B(n_134),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_666),
.B(n_136),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_666),
.B(n_140),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_674),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_674),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_699),
.B(n_688),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_691),
.B(n_667),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_692),
.B(n_688),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_692),
.B(n_700),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_697),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_709),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_709),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_694),
.B(n_680),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_690),
.B(n_695),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_701),
.B(n_671),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_710),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_718),
.B(n_682),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_716),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_712),
.B(n_692),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_714),
.B(n_704),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_711),
.B(n_696),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_713),
.B(n_698),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_R g728 ( 
.A1(n_719),
.A2(n_708),
.B(n_707),
.C(n_681),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_719),
.B(n_696),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_703),
.B1(n_720),
.B2(n_679),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_729),
.B(n_676),
.C(n_715),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_724),
.A2(n_708),
.B1(n_707),
.B2(n_693),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_727),
.Y(n_733)
);

AOI21xp33_ASAP7_75t_L g734 ( 
.A1(n_728),
.A2(n_706),
.B(n_702),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_SL g735 ( 
.A1(n_724),
.A2(n_698),
.B(n_693),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_731),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_733),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_730),
.A2(n_734),
.B(n_735),
.C(n_705),
.Y(n_738)
);

XOR2x2_ASAP7_75t_L g739 ( 
.A(n_732),
.B(n_698),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_736),
.B(n_726),
.Y(n_740)
);

OAI211xp5_ASAP7_75t_SL g741 ( 
.A1(n_740),
.A2(n_738),
.B(n_737),
.C(n_739),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_741),
.B(n_723),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_742),
.B(n_725),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_743),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_744),
.B(n_721),
.Y(n_745)
);

OA22x2_ASAP7_75t_L g746 ( 
.A1(n_745),
.A2(n_717),
.B1(n_716),
.B2(n_677),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_746),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_L g748 ( 
.A(n_747),
.B(n_142),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_748),
.Y(n_749)
);

AOI21x1_ASAP7_75t_L g750 ( 
.A1(n_749),
.A2(n_143),
.B(n_144),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_750),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_751),
.B(n_145),
.Y(n_752)
);

AOI211xp5_ASAP7_75t_L g753 ( 
.A1(n_752),
.A2(n_146),
.B(n_148),
.C(n_149),
.Y(n_753)
);


endmodule