module real_jpeg_23401_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_0),
.B(n_38),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_0),
.B(n_48),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_0),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_0),
.B(n_83),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_0),
.B(n_25),
.Y(n_214)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_2),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_2),
.B(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_2),
.B(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_7),
.B(n_27),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_7),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_7),
.B(n_83),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_7),
.B(n_51),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_7),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_8),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_8),
.B(n_48),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_8),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_8),
.B(n_83),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_9),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_9),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_9),
.B(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_9),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_9),
.B(n_51),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_12),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_12),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_12),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_83),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_12),
.B(n_51),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_12),
.B(n_48),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_12),
.B(n_38),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_12),
.B(n_27),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_13),
.B(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_51),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_13),
.B(n_102),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_13),
.B(n_48),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_13),
.B(n_38),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_13),
.B(n_27),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_13),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_13),
.B(n_108),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_14),
.B(n_48),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_14),
.B(n_38),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_14),
.B(n_51),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_14),
.B(n_83),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_14),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_14),
.B(n_27),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_14),
.B(n_25),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_14),
.B(n_108),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_32),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_15),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_155),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_15),
.B(n_83),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_15),
.B(n_51),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_16),
.B(n_51),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_16),
.B(n_48),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_16),
.B(n_83),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_16),
.B(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_16),
.B(n_38),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_16),
.B(n_27),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_16),
.B(n_25),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_16),
.B(n_302),
.Y(n_301)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_17),
.Y(n_146)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_17),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_61),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.C(n_53),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_22),
.B(n_117),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_62),
.Y(n_61)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_26),
.CI(n_30),
.CON(n_23),
.SN(n_23)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.C(n_39),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_35),
.B(n_185),
.Y(n_246)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_35),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_38),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_41),
.B(n_53),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_45),
.C(n_50),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_42),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_43),
.B(n_47),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_44),
.B(n_297),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_57),
.C(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_45),
.A2(n_50),
.B1(n_58),
.B2(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_46),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_47),
.B(n_260),
.Y(n_259)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_50),
.B(n_78),
.C(n_81),
.Y(n_115)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_51),
.Y(n_186)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_57),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_110),
.C(n_116),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_74),
.A2(n_75),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_94),
.C(n_96),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_76),
.B(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_86),
.C(n_90),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_77),
.B(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_99),
.C(n_104),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_81),
.A2(n_85),
.B1(n_99),
.B2(n_100),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_82),
.B(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_86),
.B(n_90),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.C(n_89),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_87),
.B(n_88),
.CI(n_89),
.CON(n_328),
.SN(n_328)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_90),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.CI(n_93),
.CON(n_90),
.SN(n_90)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_92),
.C(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_365),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_94),
.Y(n_365)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_106),
.C(n_109),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_98),
.B(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_99),
.A2(n_100),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_99),
.B(n_306),
.C(n_307),
.Y(n_327)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_104),
.B(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_338),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_109),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_109),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_109),
.B(n_334),
.C(n_337),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_110),
.B(n_116),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_115),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_111),
.A2(n_112),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_114),
.B(n_115),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_366),
.C(n_367),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_354),
.C(n_355),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_342),
.C(n_343),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_318),
.C(n_319),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_286),
.C(n_287),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_252),
.C(n_253),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_221),
.C(n_222),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_196),
.C(n_197),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_157),
.C(n_168),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_141),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_129),
.B(n_136),
.C(n_141),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_131),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_137),
.B(n_139),
.C(n_140),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_142),
.B(n_150),
.C(n_151),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_156),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_167),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_162),
.B1(n_167),
.B2(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_192),
.C(n_193),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.C(n_182),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_175),
.C(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_183)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.C(n_187),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_191),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_210),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_211),
.C(n_220),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_206),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_205),
.C(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_204),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_206),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.CI(n_209),
.CON(n_206),
.SN(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_208),
.C(n_209),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_220),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_218),
.B2(n_219),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_217),
.C(n_219),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_237),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_226),
.C(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_228),
.Y(n_371)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.CI(n_231),
.CON(n_228),
.SN(n_228)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_230),
.C(n_231),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_245),
.C(n_250),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_245),
.B1(n_250),
.B2(n_251),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_243),
.B(n_244),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_243),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_244),
.B(n_277),
.C(n_278),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_273),
.B2(n_285),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_274),
.C(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_258),
.C(n_266),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_262),
.C(n_265),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_264),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_270),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_314),
.C(n_315),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.CI(n_284),
.CON(n_279),
.SN(n_279)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_316),
.B2(n_317),
.Y(n_287)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_288),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_308),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_308),
.C(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_298),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_299),
.C(n_300),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_294),
.C(n_296),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_303),
.B1(n_304),
.B2(n_307),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_322),
.C(n_341),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_329),
.B2(n_341),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_327),
.C(n_328),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g370 ( 
.A(n_328),
.Y(n_370)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_332),
.C(n_333),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_340),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_336),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_337),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_353),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_347),
.C(n_353),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_350),
.C(n_351),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_358),
.C(n_363),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_362),
.B2(n_363),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_368),
.Y(n_369)
);


endmodule