module fake_jpeg_18886_n_216 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_32),
.B(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_48),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_29),
.B1(n_14),
.B2(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_46),
.B1(n_56),
.B2(n_30),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_29),
.B1(n_14),
.B2(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_29),
.B1(n_19),
.B2(n_17),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_41),
.B1(n_32),
.B2(n_22),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_14),
.B1(n_19),
.B2(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_72),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_15),
.B(n_22),
.C(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_67),
.B(n_81),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_76),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_42),
.A3(n_25),
.B1(n_15),
.B2(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_78),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_20),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_13),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_43),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_36),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_0),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_36),
.B1(n_30),
.B2(n_27),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_92),
.B1(n_95),
.B2(n_10),
.Y(n_122)
);

BUFx24_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_24),
.B(n_65),
.C(n_57),
.Y(n_91)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_28),
.B(n_1),
.C(n_2),
.D(n_4),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_5),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_7),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_71),
.B(n_83),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_115),
.B1(n_122),
.B2(n_125),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_110),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_98),
.B(n_73),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_9),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_10),
.B1(n_11),
.B2(n_97),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_11),
.B1(n_95),
.B2(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_83),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_102),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_147),
.B(n_108),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_96),
.B1(n_77),
.B2(n_76),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_111),
.B1(n_113),
.B2(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_70),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_119),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_121),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_79),
.Y(n_143)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_101),
.B1(n_115),
.B2(n_100),
.C(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_79),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_118),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_164),
.C(n_141),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_120),
.B(n_123),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_147),
.B(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_155),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_162),
.B(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_144),
.B1(n_136),
.B2(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_135),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_133),
.B(n_139),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_158),
.Y(n_182)
);

AOI32xp33_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_150),
.A3(n_129),
.B1(n_153),
.B2(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_171),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_170),
.B1(n_179),
.B2(n_152),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_178),
.C(n_163),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_145),
.B1(n_130),
.B2(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_139),
.C(n_103),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_133),
.B(n_134),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_176),
.C(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_186),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_161),
.C(n_160),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_178),
.C(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_174),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_179),
.B(n_156),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_194),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_168),
.B1(n_165),
.B2(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_196),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_183),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_187),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_190),
.A2(n_176),
.B(n_165),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_189),
.B(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_200),
.B(n_202),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_181),
.B(n_182),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_191),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_203),
.B1(n_185),
.B2(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_211),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_199),
.C(n_186),
.Y(n_211)
);

OAI221xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_109),
.B1(n_112),
.B2(n_111),
.C(n_124),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_212),
.C(n_98),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_109),
.Y(n_216)
);


endmodule