module fake_jpeg_14835_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_13),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_18),
.B1(n_14),
.B2(n_21),
.Y(n_38)
);

OAI22x1_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_24),
.B1(n_19),
.B2(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_16),
.B1(n_15),
.B2(n_25),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_13),
.B(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_12),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_43),
.B1(n_40),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_64),
.B1(n_52),
.B2(n_45),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_30),
.B(n_33),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_73),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_56),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_77),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_55),
.B1(n_50),
.B2(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_79),
.B1(n_80),
.B2(n_2),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_66),
.B1(n_65),
.B2(n_64),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_31),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_63),
.C(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_11),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_89),
.C(n_80),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_70),
.B(n_62),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_78),
.B(n_77),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_70),
.C(n_71),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_92),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_1),
.CI(n_2),
.CON(n_92),
.SN(n_92)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_4),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_98),
.C(n_86),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_5),
.C(n_6),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_85),
.C(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_108),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_103),
.B(n_8),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_101),
.B(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_9),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_9),
.B1(n_10),
.B2(n_111),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_113),
.Y(n_115)
);


endmodule