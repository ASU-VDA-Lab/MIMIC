module fake_jpeg_3371_n_174 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_56),
.B1(n_46),
.B2(n_54),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_77),
.B1(n_58),
.B2(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_50),
.B1(n_52),
.B2(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_76),
.B1(n_51),
.B2(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_55),
.B1(n_52),
.B2(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_56),
.B1(n_55),
.B2(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_60),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_0),
.Y(n_110)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_49),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_94),
.Y(n_105)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_97),
.B1(n_77),
.B2(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_49),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_62),
.B1(n_78),
.B2(n_58),
.Y(n_102)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_114),
.B1(n_96),
.B2(n_6),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_21),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_46),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_9),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_64),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_1),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_5),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_81),
.B(n_97),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_132),
.B(n_33),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_127),
.B1(n_101),
.B2(n_16),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_128),
.A3(n_135),
.B1(n_15),
.B2(n_16),
.C1(n_17),
.C2(n_19),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_5),
.B(n_6),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_29),
.B(n_30),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_44),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_8),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_8),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_108),
.B1(n_112),
.B2(n_106),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_14),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_14),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_15),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_112),
.B1(n_104),
.B2(n_101),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_129),
.C(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_156),
.C(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_154),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_161),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_138),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_162),
.A2(n_163),
.B1(n_123),
.B2(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_140),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_160),
.A2(n_142),
.B(n_153),
.C(n_130),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_145),
.C(n_151),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_166),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_168),
.B(n_159),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_164),
.B(n_119),
.Y(n_171)
);

AOI221xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_147),
.B1(n_158),
.B2(n_120),
.C(n_118),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_34),
.A3(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_42),
.Y(n_174)
);


endmodule