module fake_aes_1326_n_681 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_681);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_681;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_21), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_43), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_64), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_76), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_47), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_28), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_57), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_19), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_5), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_66), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_67), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_48), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_56), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_2), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_13), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_63), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_40), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_52), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_41), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_58), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_59), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_68), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_35), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_37), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_7), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_54), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_39), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_23), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_27), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_15), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_74), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_55), .Y(n_112) );
CKINVDCx14_ASAP7_75t_R g113 ( .A(n_24), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_4), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_72), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_42), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_6), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_3), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_29), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_98), .B(n_0), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_122), .B(n_0), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_84), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_107), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_93), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_113), .Y(n_130) );
AND2x6_ASAP7_75t_L g131 ( .A(n_88), .B(n_30), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_101), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_135) );
NAND2xp33_ASAP7_75t_L g136 ( .A(n_88), .B(n_32), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_89), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_89), .B(n_5), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_122), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_80), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_102), .B(n_6), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_101), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_77), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_78), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_119), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_79), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g151 ( .A(n_114), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_120), .B(n_8), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_81), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g154 ( .A1(n_121), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_82), .B(n_10), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_80), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_96), .B(n_11), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_99), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_104), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_106), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_108), .B(n_13), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_94), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_105), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
NOR2xp33_ASAP7_75t_SL g167 ( .A(n_142), .B(n_109), .Y(n_167) );
INVx6_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_142), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_160), .B(n_87), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_138), .B(n_123), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_165), .B(n_118), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
INVx1_ASAP7_75t_SL g179 ( .A(n_139), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_140), .B(n_112), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_139), .A2(n_109), .B1(n_83), .B2(n_116), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_124), .B(n_118), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_124), .B(n_117), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_156), .B(n_116), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_137), .A2(n_103), .B1(n_115), .B2(n_100), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_150), .B(n_115), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_131), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_126), .B(n_97), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_135), .A2(n_100), .B1(n_97), .B2(n_85), .Y(n_195) );
NOR2x1p5_ASAP7_75t_L g196 ( .A(n_130), .B(n_85), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_147), .B(n_83), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_130), .B(n_14), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_126), .B(n_38), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_133), .B(n_14), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_125), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_134), .B(n_146), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_141), .B(n_149), .Y(n_205) );
INVx5_ASAP7_75t_L g206 ( .A(n_131), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_144), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_151), .B(n_15), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_147), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_163), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_150), .B(n_16), .Y(n_212) );
INVxp67_ASAP7_75t_SL g213 ( .A(n_157), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_147), .B(n_45), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_129), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_153), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_153), .B(n_44), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_157), .B(n_16), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_129), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_132), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_159), .B(n_75), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_159), .B(n_18), .Y(n_222) );
OR2x6_ASAP7_75t_L g223 ( .A(n_154), .B(n_20), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_161), .B(n_22), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_153), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_206), .B(n_153), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_177), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_193), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_206), .B(n_193), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_179), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_194), .B(n_164), .Y(n_232) );
INVxp67_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_172), .B(n_145), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_185), .B(n_161), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_174), .A2(n_152), .B(n_162), .C(n_158), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_206), .B(n_153), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_192), .B(n_155), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_212), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_192), .B(n_131), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_211), .B(n_128), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_212), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_192), .B(n_131), .Y(n_244) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_214), .A2(n_136), .B(n_132), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_177), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_177), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_203), .B(n_131), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_168), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_168), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_206), .B(n_127), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_176), .B(n_131), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_205), .B(n_136), .Y(n_253) );
BUFx2_ASAP7_75t_L g254 ( .A(n_169), .Y(n_254) );
BUFx4f_ASAP7_75t_L g255 ( .A(n_200), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_167), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_200), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_190), .B(n_164), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_213), .B(n_163), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_204), .B(n_25), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_204), .A2(n_26), .B(n_31), .C(n_33), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_171), .B(n_34), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_188), .A2(n_36), .B1(n_46), .B2(n_49), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_169), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_166), .B(n_51), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_171), .B(n_53), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_200), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_171), .A2(n_60), .B(n_61), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_170), .B(n_73), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_178), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_219), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_220), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_208), .Y(n_275) );
CKINVDCx8_ASAP7_75t_R g276 ( .A(n_200), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_221), .B(n_65), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_175), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_178), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_197), .A2(n_71), .B(n_181), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_188), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_168), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_188), .A2(n_195), .B1(n_183), .B2(n_170), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_189), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_188), .B(n_191), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_175), .B(n_195), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_188), .B(n_223), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_218), .A2(n_207), .B(n_201), .C(n_223), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_191), .B(n_202), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_233), .B(n_199), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_284), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_254), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_268), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_287), .B(n_223), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_263), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_287), .A2(n_196), .B1(n_222), .B2(n_197), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_268), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_266), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_252), .A2(n_181), .B(n_217), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_234), .A2(n_224), .B1(n_186), .B2(n_180), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_240), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_235), .B(n_236), .Y(n_309) );
CKINVDCx11_ASAP7_75t_R g310 ( .A(n_287), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_248), .A2(n_217), .B(n_214), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_241), .A2(n_173), .B(n_182), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_266), .Y(n_313) );
AOI21x1_ASAP7_75t_L g314 ( .A1(n_244), .A2(n_184), .B(n_187), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_234), .A2(n_224), .B1(n_186), .B2(n_198), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_231), .B(n_198), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_231), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_260), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_278), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_283), .B(n_224), .Y(n_320) );
BUFx4f_ASAP7_75t_SL g321 ( .A(n_232), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_228), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_234), .A2(n_224), .B1(n_173), .B2(n_182), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_240), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_240), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_278), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_257), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_257), .B(n_224), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_228), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_253), .A2(n_209), .B(n_210), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_239), .A2(n_243), .B1(n_276), .B2(n_289), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_275), .B(n_209), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_242), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_288), .A2(n_210), .B(n_216), .C(n_225), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_286), .A2(n_178), .B1(n_216), .B2(n_225), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_269), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_255), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_269), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_307), .A2(n_255), .B1(n_285), .B2(n_238), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_318), .B(n_258), .Y(n_340) );
OA21x2_ASAP7_75t_L g341 ( .A1(n_334), .A2(n_262), .B(n_311), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_333), .A2(n_256), .B1(n_255), .B2(n_250), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_314), .A2(n_270), .B(n_277), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_296), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_302), .A2(n_277), .B(n_267), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_294), .B(n_250), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_321), .B(n_250), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_326), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_331), .A2(n_267), .B(n_280), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_309), .A2(n_262), .B(n_261), .Y(n_351) );
OAI21x1_ASAP7_75t_SL g352 ( .A1(n_307), .A2(n_265), .B(n_264), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_292), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_335), .A2(n_271), .B(n_237), .Y(n_354) );
NAND3xp33_ASAP7_75t_L g355 ( .A(n_320), .B(n_216), .C(n_225), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_298), .Y(n_356) );
NAND2xp33_ASAP7_75t_L g357 ( .A(n_295), .B(n_228), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_291), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_291), .B(n_249), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_322), .Y(n_361) );
OA21x2_ASAP7_75t_L g362 ( .A1(n_323), .A2(n_237), .B(n_226), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_294), .B(n_249), .Y(n_363) );
OA21x2_ASAP7_75t_L g364 ( .A1(n_305), .A2(n_226), .B(n_272), .Y(n_364) );
BUFx4_ASAP7_75t_R g365 ( .A(n_310), .Y(n_365) );
OA21x2_ASAP7_75t_L g366 ( .A1(n_312), .A2(n_315), .B(n_330), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_303), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_322), .Y(n_368) );
XOR2xp5_ASAP7_75t_L g369 ( .A(n_326), .B(n_249), .Y(n_369) );
OAI22xp33_ASAP7_75t_SL g370 ( .A1(n_358), .A2(n_293), .B1(n_313), .B2(n_301), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_344), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_344), .B(n_295), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_290), .B1(n_300), .B2(n_293), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_345), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_351), .A2(n_300), .B(n_299), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_350), .A2(n_329), .B(n_297), .Y(n_376) );
BUFx8_ASAP7_75t_L g377 ( .A(n_365), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_358), .A2(n_310), .B1(n_332), .B2(n_319), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_350), .A2(n_329), .B(n_297), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_345), .B(n_332), .Y(n_380) );
OAI221xp5_ASAP7_75t_SL g381 ( .A1(n_342), .A2(n_304), .B1(n_306), .B2(n_325), .C(n_324), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_369), .B(n_319), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_351), .A2(n_328), .B(n_251), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_349), .A2(n_308), .B1(n_297), .B2(n_338), .Y(n_386) );
OAI21xp33_ASAP7_75t_L g387 ( .A1(n_359), .A2(n_328), .B(n_336), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_353), .B(n_308), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_356), .B(n_328), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_352), .A2(n_245), .B(n_229), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_356), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_369), .B(n_338), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_367), .B(n_327), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_339), .A2(n_327), .B1(n_316), .B2(n_317), .Y(n_395) );
OAI21xp5_ASAP7_75t_L g396 ( .A1(n_339), .A2(n_251), .B(n_229), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_380), .B(n_367), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_385), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_371), .B(n_363), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_390), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_371), .B(n_368), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_380), .B(n_363), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_390), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_374), .B(n_368), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_374), .B(n_368), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_385), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_385), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_383), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_391), .A2(n_352), .B(n_355), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
INVx5_ASAP7_75t_L g413 ( .A(n_372), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_392), .B(n_362), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_392), .B(n_362), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_372), .B(n_361), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_394), .B(n_361), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_394), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_389), .B(n_364), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_384), .B(n_355), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_389), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_388), .B(n_364), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_373), .A2(n_347), .B1(n_357), .B2(n_360), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_395), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_424), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_420), .B(n_381), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_421), .B(n_362), .Y(n_434) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_397), .A2(n_370), .B(n_386), .C(n_393), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_424), .B(n_378), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_421), .B(n_362), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_421), .B(n_362), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_426), .B(n_382), .C(n_348), .D(n_387), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_423), .A2(n_347), .B1(n_396), .B2(n_225), .C(n_216), .Y(n_442) );
BUFx2_ASAP7_75t_SL g443 ( .A(n_426), .Y(n_443) );
AOI31xp33_ASAP7_75t_L g444 ( .A1(n_426), .A2(n_377), .A3(n_347), .B(n_337), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_398), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_429), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_427), .B(n_428), .C(n_430), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_413), .Y(n_449) );
NOR2xp67_ASAP7_75t_L g450 ( .A(n_413), .B(n_337), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_425), .B(n_364), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_406), .Y(n_452) );
OR2x6_ASAP7_75t_L g453 ( .A(n_431), .B(n_316), .Y(n_453) );
NAND2xp33_ASAP7_75t_SL g454 ( .A(n_431), .B(n_245), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_427), .B(n_341), .C(n_366), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_429), .B(n_336), .C(n_317), .D(n_259), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_409), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_413), .B(n_354), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_411), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_425), .B(n_364), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
OAI33xp33_ASAP7_75t_L g464 ( .A1(n_412), .A2(n_341), .A3(n_227), .B1(n_279), .B2(n_246), .B3(n_247), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_413), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_364), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_413), .A2(n_366), .B1(n_341), .B2(n_245), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_418), .B(n_341), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_397), .B(n_341), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_414), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_415), .Y(n_474) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_398), .B(n_366), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_414), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_418), .B(n_417), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_418), .B(n_366), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_415), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_428), .A2(n_316), .B1(n_366), .B2(n_350), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_456), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_433), .A2(n_429), .B1(n_423), .B2(n_413), .Y(n_483) );
OAI21x1_ASAP7_75t_L g484 ( .A1(n_475), .A2(n_419), .B(n_415), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_445), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_471), .B(n_416), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_471), .B(n_416), .Y(n_487) );
INVx4_ASAP7_75t_L g488 ( .A(n_445), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_477), .B(n_417), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_434), .B(n_430), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_434), .B(n_422), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_458), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_463), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_463), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_438), .B(n_422), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_477), .B(n_417), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g498 ( .A1(n_441), .A2(n_397), .B1(n_402), .B2(n_399), .C(n_408), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_435), .B(n_402), .C(n_399), .D(n_407), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_468), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_432), .B(n_401), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_433), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_436), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_438), .B(n_422), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_440), .B(n_422), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_473), .B(n_402), .Y(n_507) );
NAND2x1_ASAP7_75t_SL g508 ( .A(n_450), .B(n_405), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_445), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_436), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_436), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_448), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_440), .B(n_478), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_478), .B(n_422), .Y(n_514) );
OAI322xp33_ASAP7_75t_L g515 ( .A1(n_437), .A2(n_419), .A3(n_403), .B1(n_400), .B2(n_404), .C1(n_401), .C2(n_178), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_448), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_473), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_476), .B(n_401), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_460), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_476), .B(n_400), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_460), .B(n_403), .Y(n_521) );
OR2x6_ASAP7_75t_L g522 ( .A(n_453), .B(n_408), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_451), .B(n_403), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_472), .B(n_404), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_449), .B(n_405), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_449), .B(n_405), .Y(n_526) );
AOI211xp5_ASAP7_75t_L g527 ( .A1(n_457), .A2(n_408), .B(n_407), .C(n_404), .Y(n_527) );
BUFx3_ASAP7_75t_L g528 ( .A(n_446), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_439), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_451), .B(n_419), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_462), .B(n_405), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_462), .B(n_410), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_467), .B(n_447), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_467), .B(n_405), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_466), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_466), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_447), .B(n_407), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_519), .Y(n_538) );
NAND3xp33_ASAP7_75t_SL g539 ( .A(n_527), .B(n_442), .C(n_443), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_513), .B(n_475), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_488), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_513), .B(n_452), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_502), .B(n_453), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_492), .B(n_469), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_503), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_503), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_500), .B(n_453), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_519), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_492), .B(n_469), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_531), .B(n_452), .Y(n_550) );
NAND2xp33_ASAP7_75t_L g551 ( .A(n_483), .B(n_413), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_481), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_488), .B(n_444), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_496), .B(n_469), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_482), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_489), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_483), .B(n_455), .C(n_454), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_493), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_490), .B(n_453), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_497), .B(n_453), .Y(n_561) );
NOR2x1_ASAP7_75t_SL g562 ( .A(n_522), .B(n_443), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_499), .B(n_455), .C(n_480), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_496), .B(n_465), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_504), .B(n_465), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_504), .B(n_465), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_495), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_510), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_505), .B(n_469), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_479), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_491), .B(n_479), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_534), .B(n_479), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_520), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_498), .A2(n_413), .B1(n_459), .B2(n_464), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_528), .B(n_450), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_512), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_501), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_491), .B(n_474), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_533), .B(n_474), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_514), .B(n_474), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_533), .B(n_461), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_507), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_486), .B(n_470), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_514), .B(n_461), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_516), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_486), .B(n_461), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_579), .B(n_532), .Y(n_589) );
AOI33xp33_ASAP7_75t_L g590 ( .A1(n_584), .A2(n_532), .A3(n_487), .B1(n_536), .B2(n_535), .B3(n_530), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_542), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_575), .B(n_487), .Y(n_592) );
NOR3xp33_ASAP7_75t_SL g593 ( .A(n_553), .B(n_515), .C(n_518), .Y(n_593) );
XOR2x2_ASAP7_75t_L g594 ( .A(n_562), .B(n_508), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_542), .B(n_523), .Y(n_595) );
NAND3xp33_ASAP7_75t_SL g596 ( .A(n_557), .B(n_488), .C(n_537), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_577), .B(n_485), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_559), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_563), .A2(n_522), .B1(n_485), .B2(n_509), .C(n_537), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_575), .B(n_530), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_523), .Y(n_601) );
AOI32xp33_ASAP7_75t_L g602 ( .A1(n_551), .A2(n_509), .A3(n_506), .B1(n_525), .B2(n_526), .Y(n_602) );
INVxp33_ASAP7_75t_L g603 ( .A(n_562), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_559), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_541), .B(n_521), .Y(n_605) );
BUFx4f_ASAP7_75t_SL g606 ( .A(n_541), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_545), .Y(n_607) );
AO221x1_ASAP7_75t_L g608 ( .A1(n_551), .A2(n_506), .B1(n_522), .B2(n_510), .C(n_511), .Y(n_608) );
OA222x2_ASAP7_75t_L g609 ( .A1(n_560), .A2(n_522), .B1(n_506), .B2(n_524), .C1(n_511), .C2(n_529), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_SL g610 ( .A1(n_539), .A2(n_529), .B(n_452), .C(n_439), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_576), .B(n_538), .C(n_548), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_552), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_588), .B(n_439), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_561), .B(n_410), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_572), .B(n_484), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_572), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_555), .Y(n_617) );
OA21x2_ASAP7_75t_L g618 ( .A1(n_558), .A2(n_484), .B(n_354), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_556), .Y(n_619) );
OAI311xp33_ASAP7_75t_L g620 ( .A1(n_547), .A2(n_410), .A3(n_354), .B1(n_346), .C1(n_343), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_580), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_545), .A2(n_410), .B(n_343), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_550), .B(n_346), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_566), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_591), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_591), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_599), .B(n_543), .C(n_585), .D(n_540), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g628 ( .A1(n_596), .A2(n_573), .B1(n_580), .B2(n_568), .C1(n_586), .C2(n_582), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_590), .B(n_586), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_589), .B(n_582), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_611), .B(n_587), .C(n_578), .Y(n_631) );
XOR2x2_ASAP7_75t_L g632 ( .A(n_594), .B(n_567), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g633 ( .A(n_595), .B(n_550), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_606), .A2(n_549), .B1(n_544), .B2(n_570), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_SL g635 ( .A1(n_603), .A2(n_583), .B(n_581), .C(n_574), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_601), .B(n_549), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_596), .B(n_587), .C(n_578), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_621), .B(n_574), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_598), .Y(n_639) );
AOI32xp33_ASAP7_75t_L g640 ( .A1(n_609), .A2(n_544), .A3(n_570), .B1(n_567), .B2(n_565), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_614), .A2(n_565), .B1(n_554), .B2(n_564), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_597), .A2(n_583), .B(n_581), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_592), .B(n_571), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_604), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_616), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_606), .A2(n_564), .B1(n_554), .B2(n_571), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_636), .B(n_608), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_625), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g649 ( .A1(n_640), .A2(n_602), .B1(n_593), .B2(n_610), .C(n_605), .Y(n_649) );
NOR2xp67_ASAP7_75t_L g650 ( .A(n_646), .B(n_615), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_639), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_635), .A2(n_620), .B(n_624), .C(n_619), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_629), .B(n_617), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_638), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_628), .A2(n_593), .B1(n_612), .B2(n_600), .C(n_623), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_631), .A2(n_607), .B1(n_613), .B2(n_622), .C(n_569), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_646), .A2(n_618), .B1(n_569), .B2(n_546), .Y(n_657) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_637), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_626), .A2(n_618), .B(n_546), .Y(n_659) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_648), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_651), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_658), .A2(n_627), .B1(n_642), .B2(n_644), .C(n_641), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_647), .B(n_632), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_648), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_654), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_658), .A2(n_645), .B1(n_634), .B2(n_630), .C(n_643), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_649), .A2(n_634), .B(n_633), .Y(n_667) );
NOR2x1p5_ASAP7_75t_L g668 ( .A(n_663), .B(n_655), .Y(n_668) );
NAND3x1_ASAP7_75t_L g669 ( .A(n_662), .B(n_653), .C(n_656), .Y(n_669) );
NAND4xp25_ASAP7_75t_L g670 ( .A(n_667), .B(n_652), .C(n_650), .D(n_659), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_666), .B(n_657), .C(n_622), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_668), .Y(n_672) );
NAND4xp25_ASAP7_75t_L g673 ( .A(n_670), .B(n_665), .C(n_661), .D(n_660), .Y(n_673) );
NOR3x1_ASAP7_75t_L g674 ( .A(n_669), .B(n_660), .C(n_664), .Y(n_674) );
AND3x1_ASAP7_75t_L g675 ( .A(n_672), .B(n_671), .C(n_227), .Y(n_675) );
INVx4_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_676), .B(n_673), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_677), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_678), .A2(n_675), .B1(n_316), .B2(n_346), .Y(n_679) );
AOI31xp33_ASAP7_75t_L g680 ( .A1(n_679), .A2(n_246), .A3(n_247), .B(n_259), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_228), .B1(n_272), .B2(n_279), .C(n_343), .Y(n_681) );
endmodule