module fake_jpeg_1538_n_409 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_1),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_55),
.B(n_96),
.Y(n_141)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_60),
.Y(n_125)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_15),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_10),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_66),
.B(n_67),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_10),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_71),
.B(n_77),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_12),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_73),
.B(n_80),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_12),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_81),
.B(n_94),
.Y(n_158)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_91),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_1),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_97),
.Y(n_172)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_157)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_104),
.B(n_105),
.Y(n_150)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_106),
.B(n_57),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_110),
.Y(n_153)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_47),
.B1(n_25),
.B2(n_20),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_112),
.A2(n_117),
.B1(n_122),
.B2(n_141),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_47),
.B1(n_25),
.B2(n_34),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_113),
.A2(n_142),
.B1(n_144),
.B2(n_167),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_25),
.B1(n_34),
.B2(n_33),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_48),
.B1(n_37),
.B2(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_120),
.B(n_128),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_66),
.A2(n_101),
.B1(n_45),
.B2(n_42),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_124),
.A2(n_128),
.B1(n_133),
.B2(n_140),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_61),
.A2(n_31),
.B1(n_42),
.B2(n_37),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_85),
.B(n_31),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_129),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_33),
.B1(n_30),
.B2(n_26),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_30),
.B(n_26),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_134),
.B(n_118),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_23),
.B1(n_46),
.B2(n_28),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_63),
.A2(n_51),
.B1(n_46),
.B2(n_28),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_95),
.A2(n_21),
.B1(n_51),
.B2(n_17),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_96),
.A2(n_21),
.B1(n_17),
.B2(n_48),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_73),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_99),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_60),
.B(n_6),
.C(n_7),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_175),
.C(n_158),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_74),
.A2(n_9),
.B1(n_90),
.B2(n_97),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_76),
.A2(n_9),
.B1(n_91),
.B2(n_88),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_152),
.B1(n_161),
.B2(n_170),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_78),
.A2(n_100),
.B1(n_102),
.B2(n_107),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_58),
.B(n_72),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_176),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_109),
.A2(n_41),
.B1(n_43),
.B2(n_39),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_81),
.A2(n_55),
.B(n_80),
.C(n_73),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_120),
.B(n_128),
.Y(n_201)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_179),
.B(n_180),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_135),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_181),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_182),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_187),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_186),
.A2(n_208),
.B1(n_183),
.B2(n_178),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_111),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_SL g238 ( 
.A(n_189),
.B(n_201),
.C(n_224),
.Y(n_238)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_118),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_192),
.B(n_196),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_129),
.B(n_144),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_194),
.A2(n_163),
.B(n_165),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_138),
.B(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_197),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_147),
.B(n_136),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_198),
.B(n_204),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_111),
.B(n_115),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_202),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_129),
.B(n_128),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g246 ( 
.A1(n_200),
.A2(n_225),
.B(n_232),
.C(n_163),
.D(n_165),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_154),
.B(n_160),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_205),
.B(n_210),
.Y(n_261)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_207),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_154),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_173),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_211),
.B(n_214),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_157),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_168),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_216),
.Y(n_244)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_137),
.B(n_173),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_215),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_130),
.B(n_126),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_130),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_218),
.Y(n_273)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_220),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_159),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_164),
.B(n_159),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_170),
.B(n_161),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_139),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_227),
.B1(n_230),
.B2(n_132),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_229),
.A2(n_224),
.B1(n_230),
.B2(n_195),
.Y(n_269)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_214),
.B1(n_206),
.B2(n_227),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_116),
.B(n_163),
.Y(n_232)
);

AO22x2_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_165),
.B1(n_163),
.B2(n_116),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_237),
.B(n_274),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_217),
.B(n_194),
.C(n_208),
.Y(n_240)
);

AO22x1_ASAP7_75t_L g297 ( 
.A1(n_240),
.A2(n_238),
.B1(n_253),
.B2(n_237),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_248),
.B(n_250),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_209),
.A2(n_212),
.B1(n_213),
.B2(n_177),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_165),
.B(n_162),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_223),
.A2(n_184),
.B1(n_218),
.B2(n_228),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_184),
.A2(n_152),
.B1(n_131),
.B2(n_162),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_203),
.A2(n_219),
.B1(n_216),
.B2(n_225),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_179),
.A2(n_123),
.A3(n_131),
.B1(n_189),
.B2(n_203),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_257),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_183),
.A2(n_123),
.B(n_232),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_254),
.B1(n_252),
.B2(n_247),
.Y(n_289)
);

AOI32xp33_ASAP7_75t_L g268 ( 
.A1(n_183),
.A2(n_231),
.A3(n_221),
.B1(n_211),
.B2(n_190),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_250),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_195),
.B1(n_226),
.B2(n_181),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_192),
.A2(n_191),
.B(n_197),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_270),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_295),
.B1(n_237),
.B2(n_260),
.Y(n_308)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_207),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_283),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_234),
.A2(n_182),
.B1(n_244),
.B2(n_240),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_280),
.A2(n_288),
.B1(n_269),
.B2(n_260),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_249),
.B(n_267),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_281),
.B(n_282),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_241),
.B(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_273),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_235),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_266),
.C(n_272),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_256),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_286),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_251),
.B(n_245),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_248),
.A2(n_240),
.B1(n_257),
.B2(n_237),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_289),
.A2(n_274),
.B1(n_265),
.B2(n_258),
.Y(n_320)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g316 ( 
.A(n_290),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_246),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_298),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_233),
.B(n_262),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_296),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_294),
.A2(n_297),
.B(n_279),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_237),
.A2(n_245),
.B1(n_262),
.B2(n_261),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_238),
.B(n_255),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_242),
.B(n_263),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_271),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_301),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_243),
.B(n_263),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_239),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_259),
.B(n_274),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_242),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_259),
.Y(n_313)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_298),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_282),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_323),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_305),
.C(n_278),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_236),
.C(n_272),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_322),
.C(n_280),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_318),
.A2(n_329),
.B(n_330),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_239),
.B1(n_274),
.B2(n_236),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_319),
.A2(n_290),
.B1(n_287),
.B2(n_302),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_320),
.B(n_324),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_292),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_289),
.A2(n_275),
.B1(n_306),
.B2(n_292),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_275),
.A2(n_306),
.B1(n_292),
.B2(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_279),
.A2(n_294),
.B(n_288),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_307),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_339),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_333),
.B(n_322),
.Y(n_361)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_334),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_293),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_337),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_308),
.B1(n_319),
.B2(n_311),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_345),
.B1(n_297),
.B2(n_323),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_307),
.B(n_285),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_317),
.C(n_314),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_313),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_299),
.Y(n_340)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_311),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_341),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_329),
.A2(n_330),
.B(n_300),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_342),
.A2(n_347),
.B1(n_349),
.B2(n_309),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_324),
.A2(n_304),
.B(n_296),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_356),
.C(n_361),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_351),
.A2(n_354),
.B1(n_359),
.B2(n_345),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_325),
.A3(n_328),
.B1(n_321),
.B2(n_291),
.C1(n_312),
.C2(n_286),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_353),
.B(n_337),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_347),
.A2(n_325),
.B1(n_312),
.B2(n_321),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_338),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_336),
.A2(n_320),
.B1(n_316),
.B2(n_328),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_362),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_333),
.B(n_322),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_364),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_314),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_371),
.Y(n_381)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_357),
.Y(n_366)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_366),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_367),
.A2(n_370),
.B1(n_373),
.B2(n_339),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_359),
.A2(n_332),
.B1(n_341),
.B2(n_346),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_335),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_357),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_372),
.A2(n_374),
.B1(n_348),
.B2(n_349),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_332),
.B1(n_346),
.B2(n_344),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_317),
.C(n_343),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_363),
.C(n_361),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_369),
.A2(n_362),
.B(n_344),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_378),
.A2(n_379),
.B(n_354),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_366),
.A2(n_358),
.B(n_355),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_376),
.B(n_350),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_383),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_316),
.Y(n_384)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_384),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_348),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_334),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_391),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_389),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_382),
.A2(n_367),
.B1(n_370),
.B2(n_373),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_392),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_380),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_393),
.B(n_368),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_387),
.B1(n_390),
.B2(n_364),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_368),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_395),
.A2(n_398),
.B(n_375),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_384),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_401),
.C(n_402),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_400),
.B(n_383),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_397),
.A2(n_384),
.B1(n_316),
.B2(n_391),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_403),
.A2(n_405),
.B(n_315),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_396),
.C(n_398),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_376),
.C(n_342),
.Y(n_406)
);

OAI21x1_ASAP7_75t_SL g408 ( 
.A1(n_406),
.A2(n_407),
.B(n_327),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_310),
.Y(n_409)
);


endmodule