module fake_jpeg_22892_n_171 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_1),
.B(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_0),
.C(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_24),
.B1(n_21),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_57),
.B1(n_66),
.B2(n_27),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_24),
.B1(n_30),
.B2(n_26),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_16),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_40),
.B(n_39),
.C(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_43),
.B(n_41),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_66),
.B1(n_28),
.B2(n_23),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_76),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_87),
.Y(n_102)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_18),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_91)
);

OAI22x1_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_59),
.B1(n_95),
.B2(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_56),
.B(n_33),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_33),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_19),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_80),
.B(n_78),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_51),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_118),
.B1(n_48),
.B2(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_58),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_39),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_48),
.B1(n_55),
.B2(n_46),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_83),
.C(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_132),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_120),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_123),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_2),
.Y(n_125)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_83),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_78),
.B(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_88),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_86),
.C(n_79),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_134),
.Y(n_149)
);

NOR4xp25_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_20),
.C(n_17),
.D(n_82),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_135),
.B(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_70),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_126),
.A2(n_117),
.B1(n_118),
.B2(n_108),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_108),
.A3(n_102),
.B1(n_103),
.B2(n_109),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_148),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_128),
.B1(n_123),
.B2(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_105),
.B1(n_103),
.B2(n_70),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_127),
.A2(n_105),
.B1(n_102),
.B2(n_109),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_69),
.B(n_3),
.Y(n_146)
);

AOI21x1_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_133),
.B(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_2),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_121),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_157),
.B(n_146),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_156),
.B1(n_155),
.B2(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_144),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_137),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_153),
.B(n_145),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_162),
.B1(n_165),
.B2(n_163),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_10),
.B(n_5),
.Y(n_168)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_6),
.B(n_8),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_149),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_170),
.Y(n_171)
);


endmodule