module fake_jpeg_6654_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_33),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_1),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_51),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_25),
.B(n_29),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_56),
.B(n_59),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_52),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_25),
.B1(n_23),
.B2(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_57),
.B1(n_22),
.B2(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_53),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_27),
.B1(n_28),
.B2(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_21),
.B1(n_28),
.B2(n_26),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_24),
.B(n_26),
.C(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_29),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_71),
.B1(n_44),
.B2(n_19),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_76),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_82),
.B1(n_86),
.B2(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_44),
.C(n_58),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_19),
.C(n_55),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_46),
.B1(n_54),
.B2(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_46),
.B1(n_54),
.B2(n_47),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_54),
.B1(n_36),
.B2(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_48),
.B1(n_41),
.B2(n_34),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_68),
.B1(n_75),
.B2(n_29),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_64),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_72),
.B(n_70),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_98),
.B(n_95),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_96),
.B(n_86),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_49),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_14),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_105),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_49),
.C(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_106),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_96),
.A2(n_69),
.B1(n_61),
.B2(n_66),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_109),
.B1(n_115),
.B2(n_83),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_55),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_107),
.C(n_4),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_112),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_94),
.B1(n_80),
.B2(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_95),
.B1(n_68),
.B2(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_18),
.B1(n_15),
.B2(n_43),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_132),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_106),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_83),
.B1(n_85),
.B2(n_79),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_125),
.B(n_128),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_79),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_113),
.B1(n_102),
.B2(n_111),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_130),
.C(n_131),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_2),
.B(n_3),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_107),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_2),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_5),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_100),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_128),
.C(n_130),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_146),
.B(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_100),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_144),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_99),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_5),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_5),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_135),
.B(n_129),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_131),
.C(n_127),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_125),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_161),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_120),
.B(n_118),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_6),
.B(n_9),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_158),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_119),
.B(n_126),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_13),
.C(n_8),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_6),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_141),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_10),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_148),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_162),
.Y(n_177)
);

NAND2x1p5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_142),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_172),
.B(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_10),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_172),
.B(n_174),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_150),
.C(n_163),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_155),
.B1(n_161),
.B2(n_12),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_165),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_188),
.B(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_174),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_11),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_181),
.C(n_169),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_193),
.C(n_195),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_175),
.B1(n_176),
.B2(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_184),
.B(n_164),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_185),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_197),
.B(n_13),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_11),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_200),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_13),
.B(n_196),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_201),
.Y(n_202)
);


endmodule