module fake_jpeg_16328_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_26),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_15),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_21),
.B(n_22),
.C(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_47),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_59),
.Y(n_99)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_17),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_29),
.C(n_27),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_39),
.B1(n_15),
.B2(n_20),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_75),
.Y(n_105)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_28),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_20),
.B1(n_15),
.B2(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_76),
.B1(n_79),
.B2(n_31),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_26),
.Y(n_103)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_20),
.B1(n_28),
.B2(n_19),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_80),
.Y(n_93)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_19),
.B1(n_30),
.B2(n_31),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_41),
.Y(n_80)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_84),
.B(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_47),
.B1(n_41),
.B2(n_45),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_100),
.B1(n_56),
.B2(n_52),
.Y(n_127)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_65),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_110),
.C(n_17),
.Y(n_118)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_101),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_53),
.B1(n_34),
.B2(n_42),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_24),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_59),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_29),
.B1(n_27),
.B2(n_50),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_36),
.B(n_38),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_37),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_66),
.A3(n_27),
.B1(n_28),
.B2(n_21),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_118),
.Y(n_142)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_119),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_66),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_116),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_0),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_128),
.B(n_85),
.Y(n_163)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_60),
.A3(n_78),
.B1(n_50),
.B2(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_129),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_126),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_92),
.B1(n_123),
.B2(n_125),
.Y(n_161)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_14),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_134),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_14),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_117),
.Y(n_152)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_110),
.C(n_111),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_137),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_96),
.B1(n_92),
.B2(n_89),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_161),
.B1(n_163),
.B2(n_169),
.Y(n_178)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_159),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_148),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_105),
.B1(n_84),
.B2(n_100),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_153),
.A2(n_167),
.B1(n_168),
.B2(n_135),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_155),
.B(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_86),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_17),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_127),
.A2(n_102),
.B1(n_108),
.B2(n_89),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_108),
.B1(n_34),
.B2(n_36),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_0),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_0),
.B(n_1),
.Y(n_189)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_180),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_38),
.C(n_36),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_124),
.Y(n_179)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_181),
.A2(n_189),
.B(n_195),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_152),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_194),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_164),
.B(n_120),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_193),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_13),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_11),
.C(n_13),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_77),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_0),
.Y(n_195)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_1),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_201),
.B(n_2),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_145),
.A2(n_170),
.B(n_158),
.C(n_150),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_22),
.B(n_18),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_142),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_218),
.C(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_185),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_170),
.B(n_147),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_219),
.B(n_223),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_153),
.B1(n_139),
.B2(n_142),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_212),
.B1(n_220),
.B2(n_225),
.Y(n_231)
);

AOI22x1_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_168),
.B1(n_167),
.B2(n_169),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_199),
.B1(n_181),
.B2(n_175),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_154),
.B1(n_64),
.B2(n_61),
.Y(n_212)
);

AO32x1_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_8),
.A3(n_12),
.B1(n_11),
.B2(n_6),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_1),
.B(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_22),
.B1(n_25),
.B2(n_18),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_202),
.B1(n_200),
.B2(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_195),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_237),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_202),
.B1(n_184),
.B2(n_199),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_236),
.B1(n_196),
.B2(n_205),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_239),
.C(n_240),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_226),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_234),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_225),
.B1(n_211),
.B2(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_189),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_172),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_201),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_176),
.C(n_192),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_243),
.C(n_247),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_214),
.C(n_221),
.Y(n_243)
);

XOR2x1_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_213),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_207),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_205),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_176),
.C(n_37),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_37),
.C(n_38),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_247),
.C(n_240),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_223),
.B(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_9),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_256),
.C(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_203),
.C(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_241),
.C(n_229),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_190),
.B(n_173),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_2),
.B(n_3),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_231),
.C(n_236),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_25),
.C(n_18),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_220),
.B1(n_248),
.B2(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_263),
.B(n_10),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_180),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_270),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_271),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_171),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_190),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_25),
.B1(n_18),
.B2(n_9),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_274),
.B(n_12),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_280),
.C(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_279),
.B(n_12),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_257),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_272),
.A2(n_261),
.B1(n_254),
.B2(n_275),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_287),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_288),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_277),
.A2(n_252),
.B(n_256),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_266),
.B(n_280),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_254),
.B(n_255),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_25),
.C(n_3),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_2),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_268),
.B1(n_270),
.B2(n_267),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_290),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_285),
.C(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_293),
.B(n_7),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_301),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_24),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_302),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_24),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_309),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_303),
.B(n_292),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_288),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_310),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_282),
.C(n_290),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_311),
.A2(n_294),
.B(n_295),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_313),
.C(n_308),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_3),
.A3(n_4),
.B1(n_24),
.B2(n_296),
.C1(n_307),
.C2(n_306),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_4),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_24),
.Y(n_320)
);


endmodule