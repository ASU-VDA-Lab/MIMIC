module fake_jpeg_18164_n_199 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_32),
.B(n_34),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_20),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_27),
.B1(n_18),
.B2(n_14),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_53),
.B1(n_38),
.B2(n_21),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_27),
.B1(n_18),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_51),
.B1(n_64),
.B2(n_20),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_14),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_24),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_19),
.B1(n_30),
.B2(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_78),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_13),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_43),
.A3(n_31),
.B1(n_41),
.B2(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_13),
.Y(n_76)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_28),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_84),
.B1(n_72),
.B2(n_78),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_61),
.C(n_60),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_28),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_21),
.B1(n_19),
.B2(n_30),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_90),
.B1(n_16),
.B2(n_15),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_45),
.B1(n_62),
.B2(n_60),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_29),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_24),
.B(n_6),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_7),
.B(n_8),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_29),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_56),
.B1(n_15),
.B2(n_25),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_25),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_52),
.B(n_23),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_50),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_49),
.B(n_23),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_103),
.B1(n_109),
.B2(n_83),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_28),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_104),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_5),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_123),
.Y(n_140)
);

XNOR2x1_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_7),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_82),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_9),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_66),
.B1(n_69),
.B2(n_88),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_10),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_68),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_137),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_12),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_122),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_118),
.C(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_150),
.B(n_160),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_102),
.B(n_103),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_135),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_127),
.A2(n_124),
.B(n_126),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_137),
.B1(n_143),
.B2(n_104),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_134),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_168),
.B(n_169),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_143),
.B1(n_111),
.B2(n_117),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_171),
.B1(n_172),
.B2(n_131),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_138),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_160),
.B(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_116),
.C(n_153),
.Y(n_179)
);

AOI321xp33_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_101),
.A3(n_153),
.B1(n_113),
.B2(n_176),
.C(n_175),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_133),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_163),
.C(n_133),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_178),
.B(n_130),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_186),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_155),
.B(n_162),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_141),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_180),
.B1(n_140),
.B2(n_107),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_182),
.A3(n_174),
.B1(n_126),
.B2(n_125),
.C1(n_123),
.C2(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_114),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_68),
.C(n_125),
.Y(n_194)
);

NOR4xp25_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_191),
.C(n_119),
.D(n_123),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_66),
.B(n_69),
.Y(n_197)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_195),
.B(n_96),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_96),
.B(n_77),
.Y(n_199)
);


endmodule