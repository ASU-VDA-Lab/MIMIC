module fake_jpeg_25179_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_29),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_20),
.B(n_18),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_9),
.C(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_46),
.B(n_70),
.Y(n_82)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_59),
.B1(n_63),
.B2(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_20),
.B1(n_32),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_27),
.B1(n_32),
.B2(n_22),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_20),
.B1(n_27),
.B2(n_22),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_16),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_34),
.B(n_43),
.C(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_35),
.A2(n_26),
.B1(n_32),
.B2(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_36),
.B1(n_24),
.B2(n_19),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_55),
.B1(n_56),
.B2(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_39),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_48),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_26),
.B1(n_36),
.B2(n_21),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_81),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_65),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_93),
.B(n_34),
.Y(n_113)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_39),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_43),
.B1(n_21),
.B2(n_26),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_96),
.B1(n_34),
.B2(n_33),
.Y(n_122)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_115),
.B1(n_117),
.B2(n_120),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_107),
.Y(n_134)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_112),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_0),
.B(n_1),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_113),
.B(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_76),
.Y(n_128)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_55),
.B1(n_54),
.B2(n_49),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_119),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_68),
.B1(n_61),
.B2(n_65),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_28),
.B1(n_23),
.B2(n_24),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_19),
.B1(n_24),
.B2(n_16),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_86),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_96),
.B1(n_73),
.B2(n_84),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_124),
.A2(n_138),
.B1(n_89),
.B2(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_125),
.B(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_75),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_131),
.B(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_86),
.B1(n_84),
.B2(n_82),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_147),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_77),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_97),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_142),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_93),
.B(n_77),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_90),
.B(n_79),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_85),
.B1(n_82),
.B2(n_87),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_130),
.B1(n_144),
.B2(n_125),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_104),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_155),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_98),
.B(n_113),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_159),
.A2(n_162),
.B1(n_172),
.B2(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_105),
.B1(n_121),
.B2(n_110),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_161),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_102),
.B1(n_120),
.B2(n_93),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_99),
.B(n_93),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_89),
.C(n_80),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_171),
.C(n_132),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_177),
.B1(n_144),
.B2(n_137),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_140),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_74),
.B1(n_79),
.B2(n_90),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_67),
.C(n_58),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_28),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_34),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_127),
.A2(n_85),
.B1(n_90),
.B2(n_79),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_202),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_164),
.C(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_181),
.C(n_188),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_129),
.C(n_145),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_197),
.B1(n_201),
.B2(n_33),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_143),
.C(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_166),
.B1(n_154),
.B2(n_124),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_196),
.B1(n_205),
.B2(n_163),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_143),
.B1(n_150),
.B2(n_131),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_159),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_143),
.B1(n_149),
.B2(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_146),
.B1(n_123),
.B2(n_107),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_74),
.B1(n_146),
.B2(n_123),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_19),
.B1(n_24),
.B2(n_31),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_19),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_171),
.A2(n_58),
.B1(n_16),
.B2(n_31),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_221),
.C(n_228),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_153),
.B(n_170),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_209),
.B(n_211),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_213),
.B1(n_199),
.B2(n_205),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_162),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_155),
.B(n_152),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_174),
.B1(n_173),
.B2(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_220),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_200),
.B1(n_183),
.B2(n_194),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_224),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_151),
.B1(n_16),
.B2(n_31),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_219),
.A2(n_33),
.B1(n_30),
.B2(n_3),
.Y(n_249)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_23),
.C(n_31),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_28),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_227),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_8),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_187),
.C(n_181),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_23),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_230),
.C(n_30),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_23),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_204),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_253),
.B1(n_212),
.B2(n_221),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_248),
.A2(n_207),
.B1(n_230),
.B2(n_10),
.Y(n_270)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_218),
.Y(n_254)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_259),
.C(n_261),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_216),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_262),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_243),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_258),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_228),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_216),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_247),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_206),
.C(n_224),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_271),
.C(n_14),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_234),
.B(n_229),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_267),
.B(n_272),
.Y(n_281)
);

BUFx4f_ASAP7_75t_SL g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_30),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_14),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_236),
.B(n_253),
.Y(n_273)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_252),
.B1(n_245),
.B2(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_284),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_246),
.B(n_250),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_282),
.B(n_283),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_250),
.B(n_244),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_237),
.B(n_233),
.C(n_248),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_251),
.B(n_249),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_288),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_0),
.B(n_2),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_256),
.C(n_261),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_296),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_285),
.A2(n_263),
.B1(n_270),
.B2(n_268),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_271),
.B1(n_259),
.B2(n_4),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_301),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_282),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_275),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_308),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_281),
.B(n_275),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_304),
.A2(n_303),
.B(n_309),
.Y(n_312)
);

AOI21x1_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_297),
.B(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_295),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_13),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_288),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_299),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_313),
.C(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_294),
.C(n_298),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_11),
.C(n_12),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_4),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_5),
.B(n_6),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_309),
.B(n_6),
.C(n_7),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g325 ( 
.A1(n_322),
.A2(n_323),
.B(n_5),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_326),
.C(n_321),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_315),
.C(n_6),
.Y(n_326)
);

AOI21x1_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_324),
.B(n_6),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_7),
.B(n_308),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_7),
.Y(n_330)
);


endmodule