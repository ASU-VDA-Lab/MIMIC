module fake_jpeg_31780_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_17),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_27),
.C(n_39),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_80),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_46),
.B1(n_63),
.B2(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_0),
.Y(n_113)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_53),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_49),
.B1(n_65),
.B2(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_91),
.A2(n_58),
.B1(n_54),
.B2(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_65),
.B1(n_64),
.B2(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_100),
.B1(n_105),
.B2(n_106),
.Y(n_137)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_48),
.CI(n_70),
.CON(n_102),
.SN(n_102)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_103),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_66),
.C(n_1),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_62),
.C(n_67),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_9),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_64),
.B1(n_57),
.B2(n_61),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_111),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_47),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_29),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_8),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_2),
.B(n_3),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_126),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_98),
.Y(n_124)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_130),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_5),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_13),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_40),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_11),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_18),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_20),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_120),
.C(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_154),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_38),
.B(n_23),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_155),
.A2(n_139),
.B(n_119),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_148),
.C(n_128),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

AO32x1_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_147),
.A3(n_154),
.B1(n_151),
.B2(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_149),
.B1(n_155),
.B2(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_159),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_164),
.B1(n_168),
.B2(n_165),
.Y(n_171)
);

OAI221xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.C(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_122),
.Y(n_173)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_144),
.B(n_25),
.C(n_30),
.D(n_31),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_22),
.C(n_32),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_175),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_33),
.Y(n_177)
);


endmodule