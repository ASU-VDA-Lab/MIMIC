module fake_jpeg_28119_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2x1_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_32),
.B(n_39),
.C(n_23),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_50),
.Y(n_84)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_65),
.Y(n_81)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_33),
.B1(n_28),
.B2(n_18),
.Y(n_62)
);

AO21x1_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_32),
.B(n_16),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_40),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_28),
.B1(n_30),
.B2(n_18),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_55),
.B1(n_60),
.B2(n_63),
.Y(n_90)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

HB1xp67_ASAP7_75t_SL g111 ( 
.A(n_75),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_54),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_40),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_69),
.B1(n_71),
.B2(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_55),
.B1(n_58),
.B2(n_61),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_106),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_39),
.B1(n_28),
.B2(n_33),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_61),
.B1(n_58),
.B2(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_81),
.B1(n_82),
.B2(n_79),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_112),
.B(n_113),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_40),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_40),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_1),
.B(n_2),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_18),
.B(n_20),
.C(n_30),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

AOI22x1_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_102),
.B1(n_101),
.B2(n_112),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_23),
.B1(n_25),
.B2(n_20),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_24),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_98),
.B(n_97),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_82),
.B1(n_69),
.B2(n_47),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_129),
.B1(n_131),
.B2(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_68),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_47),
.B1(n_54),
.B2(n_51),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_68),
.B1(n_28),
.B2(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_32),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_16),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_23),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_104),
.B(n_2),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_166),
.B(n_26),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_104),
.B1(n_108),
.B2(n_91),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_159),
.B1(n_29),
.B2(n_24),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_155),
.B(n_21),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_98),
.B1(n_91),
.B2(n_104),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_148),
.B1(n_119),
.B2(n_128),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_103),
.B1(n_19),
.B2(n_22),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_37),
.C(n_36),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_153),
.C(n_37),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_37),
.C(n_36),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_19),
.B(n_22),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_167),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_1),
.B(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_127),
.B1(n_125),
.B2(n_117),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_170),
.B1(n_172),
.B2(n_191),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_120),
.B1(n_131),
.B2(n_119),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_SL g204 ( 
.A(n_171),
.B(n_176),
.C(n_183),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_129),
.B1(n_137),
.B2(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_179),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_25),
.B1(n_30),
.B2(n_26),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_178),
.B1(n_185),
.B2(n_149),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_25),
.B1(n_21),
.B2(n_26),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_24),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_153),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_21),
.B1(n_29),
.B2(n_35),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_145),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_189),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_146),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_157),
.C(n_150),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_211),
.C(n_193),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_164),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_203),
.B(n_208),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_164),
.B(n_144),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_141),
.B(n_166),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_140),
.B1(n_163),
.B2(n_29),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_170),
.B1(n_169),
.B2(n_175),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_24),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_189),
.B(n_10),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_213),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_10),
.B1(n_15),
.B2(n_3),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_212),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_181),
.C(n_182),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.C(n_225),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_182),
.C(n_179),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_174),
.B1(n_169),
.B2(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_174),
.C(n_187),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_178),
.B1(n_177),
.B2(n_34),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_231),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_1),
.B(n_2),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_196),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_35),
.C(n_34),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_207),
.C(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_234),
.B1(n_198),
.B2(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_195),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_238),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_249),
.C(n_229),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_196),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_228),
.CI(n_231),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_209),
.C(n_201),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_204),
.C(n_4),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_204),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_220),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_3),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_262),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_227),
.B1(n_216),
.B2(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_238),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_260),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_5),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_3),
.B(n_4),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_218),
.B(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_230),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_269),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_272),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_245),
.B(n_244),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_257),
.B(n_258),
.Y(n_277)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_245),
.C(n_236),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_271),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_280),
.Y(n_288)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_277),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_261),
.B(n_6),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_15),
.B(n_7),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_272),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_261),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_282),
.B(n_276),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_284),
.B(n_287),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_281),
.A2(n_263),
.B(n_266),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_278),
.B1(n_8),
.B2(n_10),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_5),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_286),
.C(n_12),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_7),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_7),
.C(n_11),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_289),
.B(n_293),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_11),
.B(n_12),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_296),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_15),
.Y(n_298)
);


endmodule