module fake_netlist_5_714_n_1893 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1893);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1893;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g194 ( 
.A(n_109),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_59),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_4),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_24),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_155),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_157),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_24),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_85),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_119),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_19),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_94),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_43),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_96),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_91),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_2),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_142),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_92),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_139),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_40),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_11),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_93),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_78),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_42),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_69),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_63),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_5),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_158),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_146),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_72),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_189),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_145),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_103),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_106),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_114),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_3),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_30),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_21),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_15),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_28),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_41),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_177),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_33),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_29),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_47),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_105),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_32),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_143),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_43),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_163),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_97),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_67),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_132),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_70),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_74),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_159),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_137),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_147),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_20),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_37),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_54),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_141),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_130),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_56),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_166),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_124),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_41),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_82),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_185),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_9),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_13),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_84),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_33),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_44),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_50),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_21),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_188),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_6),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_192),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_151),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_144),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_62),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_184),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_65),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_120),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_9),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_0),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_125),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_71),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_13),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_17),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_176),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_3),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_18),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_75),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_61),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_164),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_100),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_89),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_190),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_56),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_167),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_77),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_38),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_116),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_108),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_149),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_111),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_134),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_37),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_191),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_32),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_60),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_81),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_25),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_135),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_27),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_107),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_110),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_123),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_58),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_48),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_50),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_54),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_122),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_127),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_170),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_58),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_136),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_115),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_113),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_193),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_0),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_31),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_140),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_6),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_98),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_14),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_39),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_46),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_15),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_121),
.Y(n_361)
);

BUFx8_ASAP7_75t_SL g362 ( 
.A(n_60),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_30),
.Y(n_363)
);

INVx4_ASAP7_75t_R g364 ( 
.A(n_25),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_79),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_173),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_49),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_2),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_126),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_118),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_47),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_64),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_44),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_29),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_187),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_12),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_51),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_182),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_1),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_16),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_80),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_73),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_45),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_8),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_61),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_178),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_57),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_10),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_186),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_117),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_14),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_133),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_213),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_198),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_241),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_362),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_218),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_236),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_299),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_218),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_349),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_218),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_235),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_218),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_218),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_255),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_238),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_332),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_255),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_356),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_198),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_255),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_248),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_310),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_255),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_255),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_240),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_208),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_286),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_248),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_286),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_222),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_286),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_286),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_242),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_286),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_314),
.Y(n_427)
);

BUFx6f_ASAP7_75t_SL g428 ( 
.A(n_300),
.Y(n_428)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_227),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_378),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_261),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_245),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_353),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_274),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_246),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_274),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_249),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_390),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_353),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_237),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_319),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_237),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_256),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_274),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_250),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_250),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_262),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_251),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_251),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_265),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_282),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_269),
.Y(n_457)
);

BUFx2_ASAP7_75t_SL g458 ( 
.A(n_314),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_282),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_270),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_197),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_271),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_199),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_200),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_381),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_204),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_272),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_203),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_222),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_221),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_300),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_233),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_234),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_278),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_259),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_294),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_277),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_278),
.Y(n_479)
);

INVxp33_ASAP7_75t_L g480 ( 
.A(n_295),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_283),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_287),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_292),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_291),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_302),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_195),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_307),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_313),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_306),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_333),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_309),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_300),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_403),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_404),
.A2(n_220),
.B(n_211),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_404),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

BUFx8_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_393),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_402),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_407),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_405),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_406),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_409),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_458),
.B(n_211),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_412),
.A2(n_329),
.B(n_220),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_415),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_416),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_470),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_329),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_419),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_413),
.B(n_341),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_429),
.A2(n_355),
.B1(n_336),
.B2(n_388),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_419),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_484),
.A2(n_352),
.B1(n_223),
.B2(n_388),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_421),
.B(n_423),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_398),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_423),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_424),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_417),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_413),
.B(n_342),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_426),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_426),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_433),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_433),
.B(n_366),
.Y(n_538)
);

NAND2x1_ASAP7_75t_L g539 ( 
.A(n_434),
.B(n_364),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_434),
.B(n_196),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_436),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_425),
.B(n_194),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_443),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_420),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_427),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_432),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_444),
.B(n_366),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_414),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_488),
.A2(n_293),
.B1(n_223),
.B2(n_387),
.Y(n_553)
);

NOR3xp33_ASAP7_75t_L g554 ( 
.A(n_418),
.B(n_308),
.C(n_340),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_437),
.B(n_239),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_453),
.A2(n_389),
.B(n_210),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_441),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_427),
.B(n_359),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_452),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_456),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_445),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_461),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_399),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_463),
.B(n_201),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_401),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_447),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_428),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_447),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_542),
.B(n_455),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_513),
.B(n_458),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_567),
.B(n_540),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_497),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_493),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_497),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_495),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_513),
.B(n_389),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_495),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_498),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_503),
.Y(n_588)
);

OAI21xp33_ASAP7_75t_SL g589 ( 
.A1(n_513),
.A2(n_469),
.B(n_408),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_498),
.Y(n_590)
);

AOI21x1_ASAP7_75t_L g591 ( 
.A1(n_514),
.A2(n_212),
.B(n_202),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

AND2x2_ASAP7_75t_SL g593 ( 
.A(n_514),
.B(n_215),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_500),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_501),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_501),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_506),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_547),
.B(n_214),
.Y(n_599)
);

INVxp33_ASAP7_75t_L g600 ( 
.A(n_517),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_572),
.B(n_457),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_547),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_507),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_504),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_504),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_507),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_507),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_509),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_513),
.B(n_217),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_509),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_510),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_511),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_529),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_547),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_555),
.B(n_460),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_512),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_511),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_511),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_527),
.A2(n_293),
.B1(n_347),
.B2(n_232),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_512),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_522),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_527),
.A2(n_347),
.B1(n_352),
.B2(n_232),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_515),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_522),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_515),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_516),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_516),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_526),
.Y(n_630)
);

INVxp33_ASAP7_75t_L g631 ( 
.A(n_552),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_518),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_518),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_518),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_526),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_553),
.A2(n_360),
.B1(n_363),
.B2(n_357),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_553),
.B(n_431),
.Y(n_638)
);

INVx8_ASAP7_75t_L g639 ( 
.A(n_513),
.Y(n_639)
);

AND2x6_ASAP7_75t_L g640 ( 
.A(n_521),
.B(n_215),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_531),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_556),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_519),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_543),
.B(n_481),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_531),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_549),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_535),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_508),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_556),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_520),
.A2(n_253),
.B1(n_254),
.B2(n_252),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_508),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_521),
.B(n_482),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_525),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_519),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_530),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_535),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_549),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_523),
.B(n_463),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_536),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_530),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_567),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_525),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_514),
.A2(n_225),
.B(n_224),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_521),
.B(n_483),
.Y(n_667)
);

AND3x2_ASAP7_75t_L g668 ( 
.A(n_554),
.B(n_439),
.C(n_435),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_556),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_536),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_530),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_570),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_570),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_537),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_543),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_565),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_570),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_539),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_539),
.B(n_226),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_494),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_572),
.B(n_485),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_537),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_525),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_546),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_546),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_554),
.A2(n_357),
.B1(n_360),
.B2(n_363),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_570),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_525),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_570),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_548),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_525),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_505),
.B(n_489),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_520),
.B(n_475),
.C(n_449),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_525),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_548),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_541),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_570),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_532),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_532),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_532),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_541),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_532),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_540),
.B(n_491),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_545),
.Y(n_704)
);

CKINVDCx6p67_ASAP7_75t_R g705 ( 
.A(n_566),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_524),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_538),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_545),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_538),
.Y(n_710)
);

AND2x6_ASAP7_75t_L g711 ( 
.A(n_538),
.B(n_215),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_538),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_551),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_551),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_545),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_551),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_533),
.B(n_394),
.Y(n_717)
);

INVxp33_ASAP7_75t_SL g718 ( 
.A(n_550),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_551),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_545),
.B(n_466),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_664),
.B(n_574),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_664),
.B(n_557),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_577),
.B(n_560),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_616),
.B(n_499),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_577),
.B(n_534),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_589),
.B(n_411),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_710),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_710),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_703),
.B(n_534),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_655),
.B(n_558),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

INVx5_ASAP7_75t_L g732 ( 
.A(n_642),
.Y(n_732)
);

BUFx8_ASAP7_75t_L g733 ( 
.A(n_675),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_667),
.B(n_558),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_578),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_710),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_708),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_708),
.B(n_448),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_593),
.A2(n_514),
.B1(n_391),
.B2(n_496),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_589),
.B(n_675),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_580),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_639),
.B(n_502),
.Y(n_742)
);

AO221x1_ASAP7_75t_L g743 ( 
.A1(n_652),
.A2(n_215),
.B1(n_369),
.B2(n_479),
.C(n_361),
.Y(n_743)
);

INVx8_ASAP7_75t_L g744 ( 
.A(n_639),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_580),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_712),
.B(n_462),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_713),
.B(n_468),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_586),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_661),
.B(n_706),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_706),
.B(n_472),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_586),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_615),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_645),
.B(n_478),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_676),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_717),
.B(n_692),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_678),
.B(n_602),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_713),
.B(n_541),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_602),
.B(n_422),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_600),
.B(n_410),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_593),
.A2(n_528),
.B(n_496),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_678),
.B(n_499),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_588),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_714),
.B(n_541),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_714),
.A2(n_496),
.B(n_320),
.C(n_276),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_588),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_647),
.B(n_492),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_716),
.B(n_541),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_680),
.B(n_631),
.Y(n_768)
);

INVx8_ASAP7_75t_L g769 ( 
.A(n_639),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_639),
.B(n_312),
.Y(n_770)
);

INVx8_ASAP7_75t_L g771 ( 
.A(n_639),
.Y(n_771)
);

OA21x2_ASAP7_75t_L g772 ( 
.A1(n_591),
.A2(n_528),
.B(n_230),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_719),
.B(n_541),
.Y(n_773)
);

BUFx6f_ASAP7_75t_SL g774 ( 
.A(n_680),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_647),
.B(n_499),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_720),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_680),
.B(n_492),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_660),
.B(n_499),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_660),
.B(n_466),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_576),
.A2(n_564),
.B(n_569),
.C(n_473),
.Y(n_780)
);

OAI221xp5_ASAP7_75t_L g781 ( 
.A1(n_621),
.A2(n_564),
.B1(n_569),
.B2(n_382),
.C(n_316),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_L g782 ( 
.A(n_638),
.B(n_624),
.C(n_621),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_592),
.Y(n_783)
);

INVx8_ASAP7_75t_L g784 ( 
.A(n_575),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_576),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_615),
.B(n_480),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_579),
.B(n_544),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_615),
.B(n_201),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_582),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_582),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_593),
.A2(n_215),
.B1(n_369),
.B2(n_372),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_599),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_585),
.B(n_544),
.Y(n_793)
);

AO22x2_ASAP7_75t_L g794 ( 
.A1(n_707),
.A2(n_260),
.B1(n_247),
.B2(n_244),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_585),
.B(n_544),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_643),
.B(n_464),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_642),
.A2(n_571),
.B(n_563),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_587),
.B(n_544),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_592),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_643),
.B(n_205),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_693),
.B(n_502),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_643),
.B(n_205),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_587),
.B(n_206),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_590),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_599),
.B(n_206),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_590),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_718),
.A2(n_442),
.B1(n_430),
.B2(n_568),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_642),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_599),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_595),
.B(n_544),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_595),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_597),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_597),
.B(n_544),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_604),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_604),
.B(n_559),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_605),
.B(n_207),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_605),
.B(n_559),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_599),
.B(n_464),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_611),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_611),
.B(n_207),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_617),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_617),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_618),
.B(n_559),
.Y(n_823)
);

NOR2xp67_ASAP7_75t_SL g824 ( 
.A(n_642),
.B(n_369),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_618),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_596),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_680),
.B(n_209),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_622),
.B(n_209),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_642),
.A2(n_571),
.B(n_563),
.Y(n_829)
);

AND2x2_ASAP7_75t_SL g830 ( 
.A(n_624),
.B(n_369),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_623),
.B(n_559),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_575),
.A2(n_344),
.B1(n_346),
.B2(n_339),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_623),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_626),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_626),
.B(n_630),
.Y(n_835)
);

INVxp33_ASAP7_75t_L g836 ( 
.A(n_686),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_630),
.B(n_636),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_686),
.B(n_396),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_636),
.B(n_216),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_641),
.B(n_228),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_641),
.B(n_216),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_646),
.B(n_243),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_646),
.B(n_219),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_648),
.B(n_219),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_648),
.B(n_264),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_659),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_659),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_651),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_662),
.B(n_229),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_L g850 ( 
.A(n_601),
.B(n_438),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_662),
.B(n_266),
.Y(n_851)
);

AO22x2_ASAP7_75t_L g852 ( 
.A1(n_637),
.A2(n_674),
.B1(n_682),
.B2(n_670),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_681),
.B(n_575),
.Y(n_853)
);

BUFx5_ASAP7_75t_L g854 ( 
.A(n_640),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_679),
.B(n_465),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_670),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_594),
.B(n_524),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_596),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_674),
.B(n_267),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_682),
.B(n_268),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_668),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_684),
.B(n_279),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_684),
.B(n_280),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_685),
.B(n_284),
.Y(n_864)
);

BUFx2_ASAP7_75t_SL g865 ( 
.A(n_640),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_685),
.B(n_297),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_637),
.B(n_575),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_690),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_690),
.B(n_229),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_695),
.B(n_305),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_695),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_698),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_594),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_598),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_640),
.B(n_327),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_613),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_698),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_598),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_640),
.B(n_345),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_640),
.B(n_350),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_651),
.B(n_231),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_784),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_774),
.Y(n_883)
);

NOR3xp33_ASAP7_75t_L g884 ( 
.A(n_753),
.B(n_613),
.C(n_440),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_740),
.A2(n_575),
.B1(n_583),
.B2(n_609),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_737),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_830),
.A2(n_583),
.B1(n_609),
.B2(n_640),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_SL g888 ( 
.A(n_781),
.B(n_371),
.C(n_367),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_754),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_732),
.B(n_651),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_723),
.B(n_705),
.Y(n_891)
);

BUFx4f_ASAP7_75t_SL g892 ( 
.A(n_733),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_836),
.A2(n_583),
.B1(n_609),
.B2(n_679),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_808),
.B(n_699),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_808),
.B(n_699),
.Y(n_895)
);

AND2x4_ASAP7_75t_SL g896 ( 
.A(n_768),
.B(n_705),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_749),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_L g898 ( 
.A(n_791),
.B(n_640),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_733),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_740),
.B(n_700),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_833),
.B(n_700),
.Y(n_901)
);

INVx5_ASAP7_75t_L g902 ( 
.A(n_742),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_722),
.B(n_651),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_873),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_786),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_785),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_786),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_729),
.B(n_583),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_732),
.B(n_669),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_789),
.Y(n_910)
);

OAI21xp33_ASAP7_75t_SL g911 ( 
.A1(n_791),
.A2(n_583),
.B(n_609),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_722),
.B(n_669),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_723),
.B(n_669),
.Y(n_913)
);

OR2x2_ASAP7_75t_SL g914 ( 
.A(n_838),
.B(n_428),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_872),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_833),
.B(n_679),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_848),
.B(n_702),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_790),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_848),
.B(n_702),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_750),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_830),
.A2(n_609),
.B1(n_679),
.B2(n_669),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_758),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_804),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_806),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_725),
.B(n_679),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_876),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_731),
.B(n_465),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_752),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_776),
.B(n_732),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_721),
.B(n_669),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_776),
.B(n_704),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_777),
.B(n_278),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_811),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_732),
.B(n_296),
.Y(n_934)
);

AND2x6_ASAP7_75t_L g935 ( 
.A(n_867),
.B(n_704),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_726),
.B(n_374),
.C(n_373),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_877),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_812),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_726),
.A2(n_376),
.B(n_374),
.Y(n_939)
);

BUFx8_ASAP7_75t_L g940 ( 
.A(n_774),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_796),
.B(n_818),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_814),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_796),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_857),
.A2(n_376),
.B1(n_377),
.B2(n_379),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_809),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_835),
.B(n_709),
.Y(n_946)
);

OR2x6_ASAP7_75t_L g947 ( 
.A(n_784),
.B(n_467),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_782),
.A2(n_715),
.B1(n_709),
.B2(n_711),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_730),
.B(n_715),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_819),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_743),
.A2(n_711),
.B1(n_354),
.B2(n_392),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_784),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_818),
.B(n_467),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_734),
.B(n_581),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_792),
.A2(n_673),
.B1(n_672),
.B2(n_697),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_744),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_738),
.B(n_746),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_755),
.B(n_296),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_855),
.B(n_471),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_868),
.B(n_581),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_744),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_821),
.B(n_581),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_807),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_747),
.B(n_298),
.Y(n_964)
);

CKINVDCx14_ASAP7_75t_R g965 ( 
.A(n_759),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_727),
.Y(n_966)
);

NOR2xp67_ASAP7_75t_L g967 ( 
.A(n_832),
.B(n_677),
.Y(n_967)
);

NOR2x1p5_ASAP7_75t_L g968 ( 
.A(n_801),
.B(n_377),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_792),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_855),
.B(n_298),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_728),
.A2(n_711),
.B1(n_365),
.B2(n_375),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_766),
.B(n_301),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_861),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_853),
.B(n_348),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_822),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_736),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_742),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_825),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_794),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_852),
.A2(n_711),
.B1(n_687),
.B2(n_697),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_852),
.A2(n_687),
.B1(n_689),
.B2(n_711),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_834),
.B(n_471),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_846),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_769),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_847),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_794),
.Y(n_986)
);

OAI22xp33_ASAP7_75t_L g987 ( 
.A1(n_856),
.A2(n_348),
.B1(n_370),
.B2(n_386),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_779),
.B(n_351),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_SL g989 ( 
.A(n_827),
.B(n_380),
.C(n_379),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_871),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_769),
.B(n_473),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_788),
.B(n_370),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_852),
.A2(n_711),
.B1(n_701),
.B2(n_696),
.Y(n_993)
);

NOR2x2_ASAP7_75t_L g994 ( 
.A(n_794),
.B(n_368),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_840),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_757),
.A2(n_649),
.B(n_614),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_739),
.A2(n_837),
.B1(n_845),
.B2(n_842),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_803),
.B(n_584),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_815),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_816),
.B(n_584),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_828),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_724),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_816),
.B(n_386),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_820),
.B(n_315),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_R g1005 ( 
.A(n_770),
.B(n_591),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_820),
.B(n_839),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_850),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_756),
.B(n_474),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_769),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_735),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_817),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_823),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_839),
.B(n_317),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_788),
.B(n_257),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_831),
.Y(n_1015)
);

AND2x6_ASAP7_75t_L g1016 ( 
.A(n_762),
.B(n_603),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_761),
.B(n_474),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_765),
.Y(n_1018)
);

AND2x6_ASAP7_75t_L g1019 ( 
.A(n_783),
.B(n_603),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_851),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_775),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_844),
.B(n_476),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_881),
.A2(n_863),
.B1(n_859),
.B2(n_860),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_824),
.B(n_771),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_800),
.B(n_258),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_862),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_800),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_739),
.B(n_606),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_841),
.B(n_368),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_841),
.B(n_322),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_763),
.A2(n_649),
.B(n_614),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_799),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_864),
.B(n_606),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_778),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_866),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_802),
.A2(n_701),
.B1(n_696),
.B2(n_653),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_826),
.B(n_607),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_870),
.B(n_607),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_858),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_741),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_745),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_771),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_760),
.B(n_608),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_843),
.B(n_324),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_780),
.B(n_476),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_843),
.B(n_584),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_748),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_874),
.B(n_614),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_878),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_849),
.B(n_584),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_751),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_787),
.Y(n_1052)
);

INVxp33_ASAP7_75t_L g1053 ( 
.A(n_802),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_849),
.A2(n_696),
.B1(n_653),
.B2(n_665),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_869),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_898),
.A2(n_760),
.B(n_767),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_886),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_961),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_911),
.A2(n_805),
.B(n_764),
.C(n_773),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_915),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_984),
.B(n_614),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_937),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_SL g1063 ( 
.A1(n_1029),
.A2(n_865),
.B1(n_368),
.B2(n_380),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_905),
.B(n_907),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_900),
.B(n_793),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_1014),
.A2(n_797),
.B(n_829),
.C(n_798),
.Y(n_1066)
);

INVx3_ASAP7_75t_SL g1067 ( 
.A(n_883),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_900),
.B(n_795),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_1006),
.A2(n_880),
.B(n_879),
.C(n_875),
.Y(n_1069)
);

AO21x1_ASAP7_75t_L g1070 ( 
.A1(n_913),
.A2(n_813),
.B(n_810),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_894),
.A2(n_829),
.B(n_797),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_921),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_1072)
);

OAI22x1_ASAP7_75t_L g1073 ( 
.A1(n_891),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_961),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_965),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_904),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_957),
.B(n_772),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1032),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1025),
.A2(n_325),
.B1(n_326),
.B2(n_334),
.Y(n_1079)
);

OAI22x1_ASAP7_75t_L g1080 ( 
.A1(n_1034),
.A2(n_387),
.B1(n_331),
.B2(n_330),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1032),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1053),
.B(n_922),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_928),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_940),
.Y(n_1084)
);

OR2x6_ASAP7_75t_SL g1085 ( 
.A(n_963),
.B(n_263),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_1027),
.B(n_897),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_897),
.B(n_854),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_904),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1052),
.B(n_772),
.Y(n_1089)
);

INVx6_ASAP7_75t_L g1090 ( 
.A(n_882),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_964),
.B(n_273),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_895),
.A2(n_656),
.B(n_649),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_941),
.B(n_854),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_926),
.Y(n_1094)
);

CKINVDCx14_ASAP7_75t_R g1095 ( 
.A(n_899),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_895),
.A2(n_656),
.B(n_688),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_940),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1003),
.A2(n_490),
.B(n_477),
.C(n_487),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1010),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_992),
.A2(n_337),
.B1(n_338),
.B2(n_854),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_974),
.A2(n_653),
.B(n_701),
.C(n_683),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_R g1102 ( 
.A(n_1021),
.B(n_854),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_892),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_890),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_R g1105 ( 
.A(n_1002),
.B(n_854),
.Y(n_1105)
);

INVx5_ASAP7_75t_L g1106 ( 
.A(n_961),
.Y(n_1106)
);

NOR2x1p5_ASAP7_75t_SL g1107 ( 
.A(n_999),
.B(n_854),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_889),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_973),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1055),
.B(n_275),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_972),
.A2(n_490),
.B(n_477),
.C(n_487),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_890),
.A2(n_909),
.B(n_1028),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_920),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_931),
.B(n_610),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1055),
.B(n_281),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1040),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1042),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_908),
.A2(n_653),
.B(n_665),
.C(n_683),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_932),
.B(n_927),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_887),
.A2(n_285),
.B1(n_288),
.B2(n_289),
.Y(n_1120)
);

BUFx10_ASAP7_75t_L g1121 ( 
.A(n_896),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_906),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_979),
.A2(n_665),
.B1(n_683),
.B2(n_650),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_909),
.A2(n_694),
.B(n_688),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1017),
.A2(n_290),
.B1(n_303),
.B2(n_304),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_927),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1028),
.A2(n_694),
.B(n_688),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_959),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1004),
.A2(n_657),
.B(n_663),
.C(n_671),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_903),
.A2(n_912),
.B(n_1043),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_977),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_995),
.B(n_612),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1020),
.B(n_1026),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_928),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_910),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_914),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1035),
.B(n_612),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1043),
.A2(n_694),
.B(n_688),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_918),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_936),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_969),
.B(n_619),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_885),
.A2(n_311),
.B1(n_318),
.B2(n_321),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_986),
.A2(n_980),
.B1(n_948),
.B2(n_924),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_978),
.B(n_983),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_SL g1145 ( 
.A(n_956),
.B(n_323),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_954),
.A2(n_694),
.B(n_656),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1041),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1013),
.A2(n_625),
.B(n_658),
.C(n_650),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_943),
.B(n_683),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_949),
.A2(n_691),
.B(n_654),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_923),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1030),
.A2(n_1044),
.B(n_939),
.C(n_988),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_933),
.B(n_620),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_938),
.Y(n_1154)
);

AO22x1_ASAP7_75t_L g1155 ( 
.A1(n_884),
.A2(n_328),
.B1(n_335),
.B2(n_343),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_942),
.B(n_620),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_946),
.A2(n_691),
.B(n_654),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_946),
.A2(n_691),
.B(n_654),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_950),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_953),
.B(n_450),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_975),
.B(n_625),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_930),
.A2(n_691),
.B(n_654),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_985),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_990),
.A2(n_993),
.B1(n_888),
.B2(n_981),
.Y(n_1164)
);

BUFx8_ASAP7_75t_L g1165 ( 
.A(n_882),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_982),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_882),
.B(n_450),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1047),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_902),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_1042),
.B(n_666),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1001),
.B(n_7),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_996),
.A2(n_691),
.B(n_654),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_959),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_982),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_901),
.B(n_627),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_901),
.B(n_627),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1018),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_916),
.A2(n_644),
.B1(n_635),
.B2(n_634),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_902),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_997),
.A2(n_451),
.B1(n_454),
.B2(n_459),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_953),
.B(n_451),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_997),
.A2(n_925),
.B1(n_893),
.B2(n_1023),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_R g1183 ( 
.A(n_1042),
.B(n_66),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1051),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1008),
.B(n_454),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_945),
.B(n_561),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1031),
.A2(n_644),
.B(n_633),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_952),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1033),
.A2(n_633),
.B(n_632),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_958),
.A2(n_989),
.B(n_987),
.C(n_1022),
.Y(n_1190)
);

OAI21xp33_ASAP7_75t_L g1191 ( 
.A1(n_1017),
.A2(n_459),
.B(n_561),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_970),
.B(n_7),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1033),
.A2(n_632),
.B(n_629),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_947),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_SL g1195 ( 
.A1(n_934),
.A2(n_562),
.B(n_10),
.C(n_12),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_929),
.A2(n_629),
.B1(n_628),
.B2(n_562),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_968),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_902),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1007),
.B(n_8),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_SL g1200 ( 
.A(n_1005),
.B(n_573),
.C(n_571),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_SL g1201 ( 
.A1(n_944),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_935),
.A2(n_628),
.B1(n_573),
.B2(n_563),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_947),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_952),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1059),
.A2(n_956),
.B(n_1024),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1057),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1071),
.A2(n_917),
.B(n_919),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1119),
.B(n_1008),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1091),
.A2(n_1192),
.B1(n_1164),
.B2(n_1182),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1088),
.B(n_945),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1187),
.A2(n_917),
.B(n_919),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1182),
.A2(n_1000),
.A3(n_998),
.B(n_1050),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1076),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1064),
.B(n_1011),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1185),
.B(n_1012),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1164),
.A2(n_1152),
.B(n_1143),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1082),
.B(n_1015),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1127),
.A2(n_962),
.B(n_1048),
.Y(n_1218)
);

AOI221x1_ASAP7_75t_L g1219 ( 
.A1(n_1066),
.A2(n_1130),
.B1(n_1073),
.B2(n_1056),
.C(n_1112),
.Y(n_1219)
);

AO22x2_ASAP7_75t_L g1220 ( 
.A1(n_1142),
.A2(n_994),
.B1(n_976),
.B2(n_966),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1122),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1160),
.B(n_947),
.Y(n_1222)
);

NOR3xp33_ASAP7_75t_SL g1223 ( 
.A(n_1140),
.B(n_1049),
.C(n_1039),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_SL g1224 ( 
.A1(n_1125),
.A2(n_951),
.B(n_929),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1118),
.A2(n_1046),
.A3(n_1038),
.B(n_960),
.Y(n_1225)
);

INVx1_ASAP7_75t_SL g1226 ( 
.A(n_1088),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1065),
.B(n_935),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1065),
.B(n_935),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1077),
.A2(n_967),
.B(n_1038),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1190),
.A2(n_966),
.B(n_1036),
.C(n_1054),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1171),
.A2(n_935),
.B1(n_1045),
.B2(n_991),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1068),
.A2(n_1045),
.B(n_991),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1143),
.A2(n_1024),
.B1(n_984),
.B2(n_1009),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1101),
.A2(n_955),
.B(n_971),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1174),
.B(n_1009),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1189),
.A2(n_1037),
.B(n_1019),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1092),
.A2(n_984),
.B(n_1019),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_L g1238 ( 
.A1(n_1070),
.A2(n_573),
.B(n_1019),
.C(n_1016),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1087),
.A2(n_1037),
.B(n_1019),
.C(n_1016),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1126),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1181),
.B(n_22),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1188),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1063),
.A2(n_1037),
.B(n_1016),
.C(n_26),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1193),
.A2(n_1037),
.B(n_1016),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1079),
.B(n_1115),
.C(n_1110),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1096),
.A2(n_95),
.B(n_181),
.Y(n_1246)
);

NAND2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1058),
.B(n_90),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1172),
.A2(n_88),
.B(n_180),
.Y(n_1248)
);

AOI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1072),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.C(n_31),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1069),
.A2(n_101),
.B(n_179),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1089),
.A2(n_99),
.B(n_171),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1144),
.B(n_1086),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1146),
.A2(n_87),
.B(n_168),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1094),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1124),
.A2(n_86),
.B(n_161),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_L g1256 ( 
.A1(n_1180),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1135),
.B(n_34),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1188),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1108),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1139),
.B(n_35),
.Y(n_1260)
);

AO32x2_ASAP7_75t_L g1261 ( 
.A1(n_1180),
.A2(n_36),
.A3(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1162),
.A2(n_104),
.B(n_153),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1133),
.B(n_45),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1199),
.B(n_1120),
.C(n_1155),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1179),
.B(n_112),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1100),
.A2(n_102),
.B(n_150),
.Y(n_1266)
);

INVxp67_ASAP7_75t_SL g1267 ( 
.A(n_1132),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1157),
.A2(n_76),
.B(n_148),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1151),
.B(n_1154),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1159),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_SL g1271 ( 
.A1(n_1093),
.A2(n_46),
.B(n_49),
.C(n_51),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1114),
.A2(n_1175),
.B(n_1176),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1128),
.B(n_52),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1163),
.B(n_52),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1177),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1198),
.B(n_53),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1196),
.A2(n_55),
.A3(n_1158),
.B(n_1150),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1201),
.A2(n_1128),
.B1(n_1120),
.B2(n_1191),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1137),
.A2(n_1195),
.B(n_1178),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1060),
.B(n_1062),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1196),
.A2(n_1129),
.B(n_1148),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_SL g1282 ( 
.A(n_1058),
.B(n_1106),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1173),
.B(n_1113),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1188),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1200),
.A2(n_1104),
.B(n_1061),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1169),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1202),
.A2(n_1153),
.B(n_1161),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1131),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_R g1289 ( 
.A(n_1105),
.B(n_1102),
.Y(n_1289)
);

CKINVDCx6p67_ASAP7_75t_R g1290 ( 
.A(n_1067),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1061),
.A2(n_1141),
.B(n_1156),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1083),
.A2(n_1134),
.B(n_1149),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1099),
.B(n_1116),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1074),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1075),
.B(n_1109),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_SL g1296 ( 
.A1(n_1186),
.A2(n_1134),
.B(n_1184),
.C(n_1147),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1168),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1167),
.B(n_1194),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1058),
.B(n_1106),
.Y(n_1299)
);

NOR2xp67_ASAP7_75t_L g1300 ( 
.A(n_1058),
.B(n_1106),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1204),
.B(n_1145),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1078),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1080),
.A2(n_1072),
.A3(n_1081),
.B(n_1107),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1123),
.A2(n_1111),
.B(n_1098),
.Y(n_1304)
);

OAI22x1_ASAP7_75t_L g1305 ( 
.A1(n_1203),
.A2(n_1197),
.B1(n_1167),
.B2(n_1084),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1106),
.A2(n_1170),
.B(n_1117),
.Y(n_1306)
);

NOR4xp25_ASAP7_75t_L g1307 ( 
.A(n_1136),
.B(n_1085),
.C(n_1183),
.D(n_1165),
.Y(n_1307)
);

O2A1O1Ixp5_ASAP7_75t_L g1308 ( 
.A1(n_1090),
.A2(n_1165),
.B(n_1117),
.C(n_1074),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1090),
.A2(n_1121),
.B1(n_1095),
.B2(n_1097),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1090),
.A2(n_1182),
.A3(n_1118),
.B(n_1059),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1103),
.B(n_1121),
.C(n_1091),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1066),
.A2(n_732),
.B(n_808),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1058),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1119),
.B(n_897),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1094),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1091),
.A2(n_830),
.B1(n_782),
.B2(n_1006),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1182),
.A2(n_1118),
.A3(n_1059),
.B(n_1070),
.Y(n_1317)
);

NAND3x1_ASAP7_75t_L g1318 ( 
.A(n_1192),
.B(n_782),
.C(n_624),
.Y(n_1318)
);

O2A1O1Ixp5_ASAP7_75t_L g1319 ( 
.A1(n_1091),
.A2(n_1006),
.B(n_992),
.C(n_1014),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1091),
.B(n_957),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1088),
.Y(n_1321)
);

AOI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1056),
.A2(n_824),
.B(n_1043),
.Y(n_1322)
);

BUFx10_ASAP7_75t_L g1323 ( 
.A(n_1082),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1071),
.A2(n_1187),
.B(n_1138),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1091),
.A2(n_830),
.B1(n_1006),
.B2(n_723),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1091),
.B(n_957),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_R g1327 ( 
.A(n_1105),
.B(n_594),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1071),
.A2(n_1187),
.B(n_1138),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1182),
.A2(n_1118),
.A3(n_1059),
.B(n_1070),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1119),
.B(n_1166),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_L g1331 ( 
.A(n_1091),
.B(n_1025),
.C(n_1014),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1091),
.A2(n_911),
.B(n_1190),
.C(n_1025),
.Y(n_1332)
);

INVx5_ASAP7_75t_L g1333 ( 
.A(n_1074),
.Y(n_1333)
);

AO32x2_ASAP7_75t_L g1334 ( 
.A1(n_1182),
.A2(n_1164),
.A3(n_979),
.B1(n_1143),
.B2(n_1180),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1066),
.A2(n_732),
.B(n_808),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1119),
.B(n_1166),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1119),
.B(n_897),
.Y(n_1337)
);

AO21x1_ASAP7_75t_L g1338 ( 
.A1(n_1182),
.A2(n_1006),
.B(n_1164),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1075),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1066),
.A2(n_732),
.B(n_808),
.Y(n_1340)
);

AOI221x1_ASAP7_75t_L g1341 ( 
.A1(n_1182),
.A2(n_1164),
.B1(n_1091),
.B2(n_992),
.C(n_1014),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1091),
.A2(n_1006),
.B(n_911),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1091),
.A2(n_830),
.B1(n_1006),
.B2(n_723),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1071),
.A2(n_1187),
.B(n_1138),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1091),
.B(n_957),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1103),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1071),
.A2(n_1187),
.B(n_1138),
.Y(n_1347)
);

AOI211x1_ASAP7_75t_L g1348 ( 
.A1(n_1143),
.A2(n_1164),
.B(n_781),
.C(n_1006),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1182),
.A2(n_1164),
.B1(n_1091),
.B2(n_992),
.C(n_1014),
.Y(n_1349)
);

AOI221xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1142),
.A2(n_781),
.B1(n_939),
.B2(n_986),
.C(n_907),
.Y(n_1350)
);

AOI221xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1164),
.A2(n_986),
.B1(n_781),
.B2(n_1143),
.C(n_1006),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1091),
.B(n_957),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1056),
.A2(n_824),
.B(n_1043),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1182),
.A2(n_1118),
.A3(n_1059),
.B(n_1070),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1339),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1269),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1219),
.A2(n_1347),
.B(n_1344),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1221),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1254),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1290),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1331),
.A2(n_1345),
.B(n_1326),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1330),
.B(n_1336),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1352),
.B(n_1217),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1250),
.A2(n_1332),
.B(n_1229),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1236),
.A2(n_1244),
.B(n_1322),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1206),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1316),
.A2(n_1209),
.B1(n_1245),
.B2(n_1325),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1316),
.A2(n_1209),
.B1(n_1245),
.B2(n_1343),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1353),
.A2(n_1335),
.B(n_1312),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1342),
.A2(n_1216),
.B(n_1264),
.C(n_1214),
.Y(n_1370)
);

O2A1O1Ixp5_ASAP7_75t_L g1371 ( 
.A1(n_1266),
.A2(n_1251),
.B(n_1279),
.C(n_1238),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1249),
.A2(n_1264),
.B1(n_1263),
.B2(n_1220),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_SL g1373 ( 
.A1(n_1243),
.A2(n_1230),
.B(n_1228),
.C(n_1227),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1220),
.A2(n_1278),
.B1(n_1215),
.B2(n_1318),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1346),
.Y(n_1375)
);

AOI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1348),
.A2(n_1351),
.B1(n_1350),
.B2(n_1307),
.C(n_1278),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1333),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1256),
.A2(n_1340),
.A3(n_1272),
.B(n_1291),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1310),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1237),
.A2(n_1285),
.A3(n_1233),
.B(n_1246),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1232),
.A2(n_1281),
.B(n_1205),
.Y(n_1381)
);

INVx3_ASAP7_75t_SL g1382 ( 
.A(n_1315),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1253),
.A2(n_1255),
.B(n_1248),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1262),
.A2(n_1268),
.B(n_1292),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1314),
.B(n_1337),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1304),
.A2(n_1287),
.B(n_1234),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1333),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1333),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1270),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1234),
.A2(n_1306),
.B(n_1231),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1257),
.A2(n_1260),
.B1(n_1274),
.B2(n_1241),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1289),
.A2(n_1327),
.B1(n_1252),
.B2(n_1231),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1321),
.B(n_1208),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_SL g1394 ( 
.A(n_1224),
.B(n_1223),
.C(n_1307),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1235),
.A2(n_1308),
.B(n_1247),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1239),
.A2(n_1267),
.B(n_1224),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1310),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1323),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1323),
.B(n_1240),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1275),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1296),
.A2(n_1300),
.B(n_1299),
.Y(n_1401)
);

AOI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1348),
.A2(n_1351),
.B1(n_1271),
.B2(n_1305),
.C(n_1311),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1280),
.B(n_1210),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1297),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1283),
.B(n_1222),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1311),
.A2(n_1301),
.B1(n_1273),
.B2(n_1276),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_SL g1407 ( 
.A1(n_1282),
.A2(n_1293),
.B(n_1313),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1302),
.Y(n_1408)
);

OA21x2_ASAP7_75t_L g1409 ( 
.A1(n_1277),
.A2(n_1354),
.B(n_1329),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1242),
.A2(n_1258),
.B(n_1225),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1242),
.A2(n_1258),
.B(n_1225),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1259),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1288),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1225),
.A2(n_1310),
.B(n_1329),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1295),
.A2(n_1265),
.B(n_1313),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1284),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1265),
.A2(n_1309),
.B(n_1276),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1284),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1286),
.B(n_1212),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1277),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1309),
.A2(n_1334),
.B1(n_1261),
.B2(n_1294),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1334),
.A2(n_1261),
.B1(n_1294),
.B2(n_1212),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1317),
.A2(n_1329),
.B(n_1354),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1303),
.B(n_1334),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1317),
.A2(n_1354),
.B(n_1277),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1317),
.A2(n_1331),
.B1(n_1320),
.B2(n_1326),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1261),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1207),
.A2(n_1211),
.B(n_1218),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1217),
.B(n_1226),
.Y(n_1429)
);

AOI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1320),
.A2(n_1352),
.B1(n_1345),
.B2(n_1326),
.C(n_1343),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1331),
.B(n_1209),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1219),
.A2(n_1328),
.B(n_1324),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1310),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1332),
.A2(n_808),
.B(n_1331),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1331),
.A2(n_1319),
.B(n_1320),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1346),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1331),
.A2(n_830),
.B1(n_1209),
.B2(n_1320),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1316),
.A2(n_911),
.B(n_1326),
.C(n_1320),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1226),
.Y(n_1441)
);

CKINVDCx12_ASAP7_75t_R g1442 ( 
.A(n_1298),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1443)
);

O2A1O1Ixp33_ASAP7_75t_SL g1444 ( 
.A1(n_1332),
.A2(n_1331),
.B(n_1343),
.C(n_1325),
.Y(n_1444)
);

INVxp67_ASAP7_75t_SL g1445 ( 
.A(n_1338),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1269),
.Y(n_1446)
);

INVx8_ASAP7_75t_L g1447 ( 
.A(n_1333),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1331),
.A2(n_1319),
.B(n_1320),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1221),
.Y(n_1449)
);

BUFx8_ASAP7_75t_L g1450 ( 
.A(n_1213),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1219),
.A2(n_1328),
.B(n_1324),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1331),
.A2(n_830),
.B1(n_1209),
.B2(n_1320),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1269),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1219),
.A2(n_1328),
.B(n_1324),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1269),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1213),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1331),
.A2(n_1319),
.B(n_1320),
.Y(n_1457)
);

AOI21xp33_ASAP7_75t_L g1458 ( 
.A1(n_1331),
.A2(n_1326),
.B(n_1320),
.Y(n_1458)
);

AO22x2_ASAP7_75t_L g1459 ( 
.A1(n_1341),
.A2(n_1349),
.B1(n_1325),
.B2(n_1343),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1207),
.A2(n_1211),
.B(n_1218),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1331),
.B(n_1320),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1269),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1333),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1219),
.A2(n_1328),
.B(n_1324),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1221),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1219),
.A2(n_1328),
.B(n_1324),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1269),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1269),
.Y(n_1468)
);

NAND2x1_ASAP7_75t_L g1469 ( 
.A(n_1205),
.B(n_1313),
.Y(n_1469)
);

OR2x6_ASAP7_75t_L g1470 ( 
.A(n_1205),
.B(n_1348),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1316),
.A2(n_911),
.B(n_1326),
.C(n_1320),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1221),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1314),
.B(n_1337),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1314),
.B(n_1337),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1207),
.A2(n_1211),
.B(n_1218),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1207),
.A2(n_1211),
.B(n_1218),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1221),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1331),
.A2(n_1319),
.B(n_1320),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1331),
.A2(n_830),
.B1(n_1209),
.B2(n_1320),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1331),
.A2(n_1245),
.B1(n_753),
.B2(n_1091),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1331),
.A2(n_1319),
.B(n_1320),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1333),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1331),
.B(n_1326),
.C(n_1320),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1331),
.A2(n_1245),
.B1(n_753),
.B2(n_1091),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1254),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1444),
.A2(n_1431),
.B(n_1367),
.C(n_1368),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1473),
.B(n_1474),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1366),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1399),
.B(n_1429),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1419),
.B(n_1431),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1440),
.A2(n_1471),
.B(n_1480),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1485),
.A2(n_1372),
.B1(n_1479),
.B2(n_1438),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1386),
.A2(n_1371),
.B(n_1369),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1374),
.B(n_1393),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1372),
.A2(n_1438),
.B1(n_1452),
.B2(n_1479),
.Y(n_1496)
);

AOI31xp33_ASAP7_75t_L g1497 ( 
.A1(n_1452),
.A2(n_1376),
.A3(n_1374),
.B(n_1402),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1444),
.A2(n_1434),
.B(n_1364),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1379),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1371),
.A2(n_1425),
.B(n_1420),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1355),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1406),
.A2(n_1391),
.B1(n_1443),
.B2(n_1439),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1377),
.Y(n_1503)
);

O2A1O1Ixp5_ASAP7_75t_L g1504 ( 
.A1(n_1445),
.A2(n_1478),
.B(n_1435),
.C(n_1481),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1430),
.B(n_1461),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1434),
.A2(n_1364),
.B(n_1440),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1405),
.B(n_1412),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1412),
.B(n_1403),
.Y(n_1508)
);

OAI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1461),
.A2(n_1391),
.B1(n_1361),
.B2(n_1448),
.C(n_1457),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1417),
.B(n_1356),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1446),
.B(n_1453),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1430),
.B(n_1363),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1455),
.B(n_1462),
.Y(n_1513)
);

AOI21x1_ASAP7_75t_SL g1514 ( 
.A1(n_1397),
.A2(n_1433),
.B(n_1424),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1471),
.A2(n_1370),
.B(n_1484),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1406),
.A2(n_1437),
.B1(n_1482),
.B2(n_1376),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1355),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1389),
.B(n_1400),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1458),
.A2(n_1426),
.B(n_1394),
.C(n_1392),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1467),
.B(n_1468),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1377),
.A2(n_1387),
.B(n_1463),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1445),
.A2(n_1402),
.B(n_1396),
.C(n_1422),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1459),
.A2(n_1399),
.B1(n_1470),
.B2(n_1392),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1410),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1441),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1414),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1449),
.B(n_1465),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1472),
.B(n_1477),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1358),
.B(n_1456),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1404),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1411),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1469),
.A2(n_1396),
.B(n_1470),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1373),
.A2(n_1421),
.B1(n_1422),
.B2(n_1408),
.C(n_1427),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1395),
.B(n_1416),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1409),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1382),
.A2(n_1407),
.B(n_1359),
.C(n_1486),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1390),
.A2(n_1423),
.B(n_1401),
.C(n_1447),
.Y(n_1537)
);

O2A1O1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1382),
.A2(n_1413),
.B(n_1401),
.C(n_1381),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1450),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1409),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1409),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1450),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1398),
.Y(n_1543)
);

NOR2xp67_ASAP7_75t_L g1544 ( 
.A(n_1436),
.B(n_1418),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1428),
.A2(n_1460),
.B(n_1476),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1360),
.A2(n_1388),
.B1(n_1483),
.B2(n_1463),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1387),
.B(n_1483),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1387),
.A2(n_1463),
.B(n_1483),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1360),
.A2(n_1388),
.B1(n_1483),
.B2(n_1387),
.Y(n_1549)
);

AND2x4_ASAP7_75t_SL g1550 ( 
.A(n_1375),
.B(n_1442),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1447),
.A2(n_1381),
.B(n_1357),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1398),
.B(n_1388),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1375),
.A2(n_1466),
.B(n_1432),
.C(n_1464),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1451),
.A2(n_1454),
.B(n_1464),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1555)
);

OA22x2_ASAP7_75t_L g1556 ( 
.A1(n_1384),
.A2(n_1365),
.B1(n_1383),
.B2(n_1475),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1380),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1380),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1444),
.A2(n_1332),
.B(n_1326),
.C(n_1320),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1386),
.A2(n_1371),
.B(n_1369),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1385),
.B(n_1419),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1415),
.B(n_1362),
.Y(n_1562)
);

BUFx12f_ASAP7_75t_L g1563 ( 
.A(n_1436),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1444),
.A2(n_1332),
.B(n_1326),
.C(n_1320),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_SL g1565 ( 
.A1(n_1440),
.A2(n_1332),
.B(n_1341),
.Y(n_1565)
);

O2A1O1Ixp5_ASAP7_75t_L g1566 ( 
.A1(n_1371),
.A2(n_1331),
.B(n_1368),
.C(n_1367),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1386),
.A2(n_1371),
.B(n_1369),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1480),
.A2(n_1485),
.B1(n_1331),
.B2(n_1326),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1385),
.B(n_1419),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1385),
.B(n_1419),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1385),
.B(n_1419),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1444),
.A2(n_1332),
.B(n_1326),
.C(n_1320),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1450),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1430),
.B(n_1461),
.Y(n_1574)
);

NAND2xp33_ASAP7_75t_L g1575 ( 
.A(n_1480),
.B(n_1331),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1430),
.B(n_1461),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1379),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1415),
.B(n_1362),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1480),
.A2(n_1485),
.B1(n_1331),
.B2(n_1326),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1555),
.B(n_1535),
.Y(n_1580)
);

AO21x2_ASAP7_75t_L g1581 ( 
.A1(n_1498),
.A2(n_1506),
.B(n_1554),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1499),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1524),
.B(n_1531),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1532),
.B(n_1565),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1540),
.B(n_1541),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1505),
.A2(n_1576),
.B1(n_1574),
.B2(n_1497),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1489),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1534),
.Y(n_1588)
);

AO21x2_ASAP7_75t_L g1589 ( 
.A1(n_1537),
.A2(n_1522),
.B(n_1551),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1566),
.A2(n_1504),
.B(n_1522),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1500),
.B(n_1558),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1557),
.B(n_1526),
.Y(n_1592)
);

OR2x6_ASAP7_75t_L g1593 ( 
.A(n_1492),
.B(n_1515),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1526),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1545),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1533),
.A2(n_1523),
.B(n_1530),
.Y(n_1596)
);

AOI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1493),
.A2(n_1496),
.B1(n_1487),
.B2(n_1579),
.C(n_1568),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1545),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1494),
.B(n_1560),
.Y(n_1599)
);

AOI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1556),
.A2(n_1512),
.B(n_1516),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1494),
.B(n_1560),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1518),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1560),
.B(n_1567),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1553),
.B(n_1538),
.Y(n_1604)
);

AO21x2_ASAP7_75t_L g1605 ( 
.A1(n_1575),
.A2(n_1519),
.B(n_1509),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1491),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1530),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1561),
.B(n_1569),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1567),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1508),
.B(n_1507),
.Y(n_1610)
);

OAI211xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1559),
.A2(n_1564),
.B(n_1572),
.C(n_1502),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1527),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1510),
.B(n_1520),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1562),
.B(n_1578),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1567),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1528),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1511),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1488),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_1608),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1608),
.B(n_1513),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1594),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1593),
.A2(n_1586),
.B1(n_1605),
.B2(n_1590),
.Y(n_1624)
);

NAND2x1_ASAP7_75t_L g1625 ( 
.A(n_1593),
.B(n_1584),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1588),
.B(n_1583),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1587),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1606),
.B(n_1529),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1536),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1585),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1587),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1597),
.B(n_1490),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_SL g1633 ( 
.A1(n_1593),
.A2(n_1495),
.B1(n_1550),
.B2(n_1539),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1593),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1595),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1606),
.B(n_1525),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1586),
.A2(n_1517),
.B1(n_1549),
.B2(n_1546),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1582),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1593),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1591),
.B(n_1514),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1591),
.B(n_1581),
.Y(n_1641)
);

OAI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1632),
.A2(n_1597),
.B1(n_1584),
.B2(n_1604),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1627),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1627),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1622),
.B(n_1613),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1620),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1631),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1626),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1631),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1632),
.A2(n_1584),
.B1(n_1604),
.B2(n_1590),
.Y(n_1650)
);

OAI31xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1624),
.A2(n_1611),
.A3(n_1605),
.B(n_1615),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1624),
.A2(n_1605),
.B(n_1611),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1639),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1641),
.A2(n_1605),
.B1(n_1613),
.B2(n_1614),
.C(n_1602),
.Y(n_1654)
);

AND2x2_ASAP7_75t_SL g1655 ( 
.A(n_1639),
.B(n_1590),
.Y(n_1655)
);

CKINVDCx16_ASAP7_75t_R g1656 ( 
.A(n_1621),
.Y(n_1656)
);

OAI211xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1633),
.A2(n_1602),
.B(n_1552),
.C(n_1614),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1630),
.B(n_1628),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_L g1659 ( 
.A(n_1633),
.B(n_1600),
.C(n_1634),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1636),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1637),
.A2(n_1584),
.B1(n_1604),
.B2(n_1590),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1637),
.B(n_1590),
.C(n_1604),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1639),
.A2(n_1584),
.B1(n_1589),
.B2(n_1604),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1625),
.B(n_1604),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1641),
.A2(n_1612),
.B1(n_1617),
.B2(n_1607),
.C(n_1618),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1622),
.B(n_1610),
.Y(n_1666)
);

INVx5_ASAP7_75t_SL g1667 ( 
.A(n_1629),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1641),
.A2(n_1612),
.B1(n_1617),
.B2(n_1607),
.C(n_1618),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1626),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1639),
.A2(n_1589),
.B1(n_1615),
.B2(n_1596),
.Y(n_1670)
);

OA21x2_ASAP7_75t_L g1671 ( 
.A1(n_1635),
.A2(n_1609),
.B(n_1601),
.Y(n_1671)
);

OAI21xp33_ASAP7_75t_L g1672 ( 
.A1(n_1640),
.A2(n_1600),
.B(n_1592),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1634),
.B(n_1501),
.C(n_1503),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1635),
.A2(n_1609),
.B(n_1603),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1625),
.B(n_1629),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1639),
.A2(n_1550),
.B(n_1542),
.C(n_1539),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1640),
.A2(n_1603),
.B(n_1601),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1638),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1623),
.Y(n_1679)
);

OAI31xp33_ASAP7_75t_L g1680 ( 
.A1(n_1640),
.A2(n_1543),
.A3(n_1592),
.B(n_1615),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1656),
.B(n_1542),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1645),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1643),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1643),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1644),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1671),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1662),
.A2(n_1629),
.B(n_1589),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1676),
.B(n_1573),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1678),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1652),
.A2(n_1601),
.B(n_1599),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1675),
.Y(n_1691)
);

INVx4_ASAP7_75t_SL g1692 ( 
.A(n_1653),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1664),
.B(n_1629),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1661),
.A2(n_1629),
.B(n_1581),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1678),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1674),
.Y(n_1696)
);

INVx4_ASAP7_75t_SL g1697 ( 
.A(n_1653),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1677),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1677),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1646),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

OA21x2_ASAP7_75t_L g1702 ( 
.A1(n_1672),
.A2(n_1616),
.B(n_1598),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1647),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1679),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1653),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1649),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1649),
.Y(n_1707)
);

NOR2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1648),
.B(n_1573),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1658),
.B(n_1636),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1683),
.Y(n_1710)
);

NAND2x1_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1679),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1686),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1687),
.A2(n_1651),
.B(n_1654),
.C(n_1663),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1709),
.B(n_1658),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1694),
.A2(n_1642),
.B(n_1650),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1708),
.B(n_1692),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1688),
.B(n_1563),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1701),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1682),
.B(n_1660),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1684),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1684),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1700),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1704),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1708),
.B(n_1669),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1691),
.B(n_1669),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1691),
.B(n_1669),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1692),
.B(n_1655),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1685),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1692),
.B(n_1655),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1692),
.B(n_1675),
.Y(n_1732)
);

NOR2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1709),
.B(n_1639),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1695),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1704),
.B(n_1666),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1695),
.B(n_1665),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1692),
.B(n_1667),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1686),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1686),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1681),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1689),
.B(n_1668),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1686),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1703),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1697),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1690),
.B(n_1636),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1693),
.A2(n_1659),
.B1(n_1673),
.B2(n_1657),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1696),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1697),
.B(n_1675),
.Y(n_1748)
);

AOI21xp33_ASAP7_75t_L g1749 ( 
.A1(n_1713),
.A2(n_1690),
.B(n_1702),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1740),
.B(n_1501),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1734),
.B(n_1628),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1740),
.B(n_1621),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_SL g1753 ( 
.A(n_1715),
.B(n_1701),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1736),
.B(n_1706),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1724),
.B(n_1706),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1721),
.B(n_1619),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1725),
.B(n_1707),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1710),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1711),
.A2(n_1694),
.B(n_1690),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1710),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1716),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1720),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1720),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1719),
.B(n_1735),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1746),
.A2(n_1664),
.B1(n_1693),
.B2(n_1670),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1737),
.B(n_1697),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1722),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1722),
.Y(n_1768)
);

OR2x6_ASAP7_75t_L g1769 ( 
.A(n_1744),
.B(n_1711),
.Y(n_1769)
);

NOR2x1_ASAP7_75t_L g1770 ( 
.A(n_1744),
.B(n_1701),
.Y(n_1770)
);

AOI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1741),
.A2(n_1702),
.B(n_1701),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1737),
.B(n_1697),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1727),
.Y(n_1773)
);

OAI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1745),
.A2(n_1629),
.B1(n_1664),
.B2(n_1693),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1723),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1716),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1718),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1716),
.B(n_1697),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1723),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1730),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1735),
.B(n_1714),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1717),
.B(n_1705),
.Y(n_1782)
);

INVxp67_ASAP7_75t_SL g1783 ( 
.A(n_1718),
.Y(n_1783)
);

OA21x2_ASAP7_75t_L g1784 ( 
.A1(n_1712),
.A2(n_1699),
.B(n_1698),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1730),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1769),
.B(n_1729),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1766),
.B(n_1729),
.Y(n_1787)
);

BUFx2_ASAP7_75t_L g1788 ( 
.A(n_1770),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1758),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1772),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1784),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1760),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1769),
.B(n_1731),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1784),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1778),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1769),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1762),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1753),
.A2(n_1749),
.B(n_1759),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1761),
.B(n_1731),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1781),
.B(n_1714),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1763),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1777),
.Y(n_1802)
);

NAND2xp33_ASAP7_75t_L g1803 ( 
.A(n_1764),
.B(n_1733),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1773),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1751),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1776),
.B(n_1732),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1767),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1783),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1768),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1750),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1757),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1757),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1804),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1790),
.B(n_1752),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1790),
.B(n_1754),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1804),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_SL g1817 ( 
.A(n_1786),
.B(n_1753),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1809),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1809),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1796),
.B(n_1754),
.Y(n_1820)
);

AOI221x1_ASAP7_75t_L g1821 ( 
.A1(n_1798),
.A2(n_1749),
.B1(n_1771),
.B2(n_1718),
.C(n_1782),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1800),
.B(n_1756),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1798),
.A2(n_1771),
.B(n_1765),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1808),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1788),
.A2(n_1680),
.B(n_1748),
.C(n_1732),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1810),
.A2(n_1755),
.B(n_1774),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1787),
.B(n_1726),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1810),
.A2(n_1755),
.B1(n_1745),
.B2(n_1785),
.C(n_1779),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1809),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1788),
.A2(n_1693),
.B1(n_1732),
.B2(n_1748),
.Y(n_1830)
);

XOR2xp5_ASAP7_75t_L g1831 ( 
.A(n_1787),
.B(n_1748),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1796),
.B(n_1775),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1809),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1824),
.B(n_1808),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1827),
.B(n_1799),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1813),
.B(n_1795),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1824),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1816),
.B(n_1795),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1818),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1817),
.A2(n_1803),
.B1(n_1799),
.B2(n_1806),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1827),
.B(n_1806),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1814),
.B(n_1811),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1819),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1831),
.B(n_1806),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1826),
.B(n_1811),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1845),
.A2(n_1823),
.B(n_1821),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1834),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1842),
.B(n_1820),
.Y(n_1848)
);

NOR2x1_ASAP7_75t_L g1849 ( 
.A(n_1834),
.B(n_1829),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1835),
.B(n_1832),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1837),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1841),
.B(n_1815),
.Y(n_1852)
);

NAND3xp33_ASAP7_75t_L g1853 ( 
.A(n_1840),
.B(n_1825),
.C(n_1828),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1844),
.B(n_1812),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1836),
.B(n_1812),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1838),
.A2(n_1825),
.B(n_1830),
.Y(n_1856)
);

O2A1O1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1846),
.A2(n_1839),
.B(n_1843),
.C(n_1833),
.Y(n_1857)
);

AOI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1853),
.A2(n_1793),
.B(n_1786),
.Y(n_1858)
);

AOI221x1_ASAP7_75t_L g1859 ( 
.A1(n_1851),
.A2(n_1802),
.B1(n_1807),
.B2(n_1789),
.C(n_1792),
.Y(n_1859)
);

AOI322xp5_ASAP7_75t_L g1860 ( 
.A1(n_1848),
.A2(n_1786),
.A3(n_1793),
.B1(n_1791),
.B2(n_1794),
.C1(n_1806),
.C2(n_1801),
.Y(n_1860)
);

O2A1O1Ixp5_ASAP7_75t_L g1861 ( 
.A1(n_1856),
.A2(n_1854),
.B(n_1793),
.C(n_1850),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1849),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1855),
.A2(n_1852),
.B1(n_1847),
.B2(n_1805),
.C(n_1822),
.Y(n_1863)
);

AOI211xp5_ASAP7_75t_L g1864 ( 
.A1(n_1846),
.A2(n_1807),
.B(n_1801),
.C(n_1789),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1862),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1860),
.B(n_1792),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1858),
.B(n_1805),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1859),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1861),
.Y(n_1869)
);

BUFx12f_ASAP7_75t_L g1870 ( 
.A(n_1863),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1864),
.B(n_1805),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1868),
.B(n_1857),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_R g1873 ( 
.A1(n_1865),
.A2(n_1802),
.B1(n_1794),
.B2(n_1791),
.Y(n_1873)
);

AOI211xp5_ASAP7_75t_L g1874 ( 
.A1(n_1866),
.A2(n_1797),
.B(n_1802),
.C(n_1544),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1867),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_SL g1876 ( 
.A(n_1870),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1873),
.Y(n_1877)
);

INVxp33_ASAP7_75t_L g1878 ( 
.A(n_1872),
.Y(n_1878)
);

OAI22xp33_ASAP7_75t_SL g1879 ( 
.A1(n_1875),
.A2(n_1866),
.B1(n_1871),
.B2(n_1869),
.Y(n_1879)
);

AND3x2_ASAP7_75t_L g1880 ( 
.A(n_1877),
.B(n_1874),
.C(n_1876),
.Y(n_1880)
);

AOI322xp5_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1879),
.A3(n_1878),
.B1(n_1791),
.B2(n_1794),
.C1(n_1797),
.C2(n_1742),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1881),
.B(n_1800),
.Y(n_1882)
);

XNOR2xp5_ASAP7_75t_L g1883 ( 
.A(n_1881),
.B(n_1780),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1883),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1882),
.B(n_1727),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1885),
.A2(n_1738),
.B1(n_1739),
.B2(n_1747),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1884),
.A2(n_1738),
.B1(n_1742),
.B2(n_1747),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1887),
.Y(n_1888)
);

OAI22x1_ASAP7_75t_SL g1889 ( 
.A1(n_1888),
.A2(n_1886),
.B1(n_1712),
.B2(n_1739),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_SL g1890 ( 
.A1(n_1889),
.A2(n_1705),
.B1(n_1728),
.B2(n_1726),
.Y(n_1890)
);

INVxp67_ASAP7_75t_L g1891 ( 
.A(n_1890),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1891),
.A2(n_1728),
.B1(n_1705),
.B2(n_1743),
.Y(n_1892)
);

AOI211xp5_ASAP7_75t_L g1893 ( 
.A1(n_1892),
.A2(n_1548),
.B(n_1521),
.C(n_1547),
.Y(n_1893)
);


endmodule