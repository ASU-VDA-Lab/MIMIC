module fake_netlist_5_1951_n_98 (n_16, n_0, n_12, n_9, n_25, n_18, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_98);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_98;

wire n_91;
wire n_82;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_45;
wire n_46;
wire n_94;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_29;
wire n_79;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_77;
wire n_64;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_0),
.A2(n_15),
.B1(n_11),
.B2(n_1),
.Y(n_30)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_1),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_14),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_18),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_4),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_26),
.B(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_29),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_29),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_58),
.B(n_49),
.C(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_32),
.B(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_33),
.Y(n_70)
);

NAND2x1p5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_31),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_40),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVxp67_ASAP7_75t_SL g82 ( 
.A(n_81),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_76),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

AOI211x1_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_75),
.B(n_78),
.C(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_72),
.C(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_77),
.Y(n_92)
);

AOI221xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_38),
.B1(n_89),
.B2(n_64),
.C(n_70),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_70),
.B1(n_43),
.B2(n_48),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_93),
.Y(n_97)
);

OR2x6_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_96),
.Y(n_98)
);


endmodule