module fake_jpeg_29368_n_171 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx3_ASAP7_75t_SL g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx3_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_16),
.B(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_26),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_66),
.Y(n_85)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_78),
.Y(n_80)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_48),
.B1(n_69),
.B2(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_82),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_90),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_52),
.B1(n_64),
.B2(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_50),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_69),
.B1(n_68),
.B2(n_51),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_49),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_63),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_110),
.Y(n_133)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_63),
.B1(n_45),
.B2(n_56),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_45),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_111),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_2),
.C(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_60),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_15),
.B(n_41),
.C(n_36),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_113),
.B(n_7),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_109),
.B(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_0),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_1),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_6),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_22),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_138),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_144),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_125),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_14),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_124),
.Y(n_156)
);

XOR2x2_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_153),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_114),
.C(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_161),
.C(n_152),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_152),
.A2(n_143),
.B1(n_137),
.B2(n_150),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_157),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_163),
.A2(n_164),
.B1(n_161),
.B2(n_154),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_159),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_158),
.B(n_141),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_142),
.B(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_21),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_27),
.Y(n_171)
);


endmodule