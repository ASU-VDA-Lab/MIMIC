module fake_netlist_5_1999_n_964 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_964);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_964;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_620;
wire n_367;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_368;
wire n_247;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_568;
wire n_509;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_579;
wire n_394;
wire n_250;
wire n_341;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_291;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_395;
wire n_553;
wire n_432;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_866;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_477;
wire n_571;
wire n_461;
wire n_693;
wire n_333;
wire n_338;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_891;
wire n_239;
wire n_466;
wire n_630;
wire n_420;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_647;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_857;
wire n_832;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_129),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_99),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_39),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_94),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_143),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_93),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_41),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_9),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_74),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_45),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_114),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_49),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_170),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_123),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_192),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_111),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_27),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_51),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_64),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_83),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_151),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_154),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_136),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_113),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_160),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_56),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_220),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_148),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_65),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_102),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_180),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_28),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_120),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_69),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_198),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_199),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_159),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_145),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_209),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_183),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_165),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_171),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_217),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_162),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_109),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_130),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_221),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_189),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_90),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_75),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_73),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_127),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_3),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_196),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_202),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_98),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_38),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_70),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_71),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_62),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_108),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_18),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_1),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_166),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_218),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_193),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_215),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_116),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_100),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_104),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_16),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_115),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_152),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_67),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_128),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_76),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_24),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_18),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_150),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_204),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_52),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_97),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_141),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_91),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_203),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_140),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_226),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_149),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_107),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_216),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_137),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_101),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_228),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_60),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_153),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_13),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_50),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_118),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_163),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_20),
.B(n_186),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_119),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_161),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_122),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_173),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_213),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_124),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_117),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_144),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_72),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_229),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_42),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_14),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_35),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_58),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_133),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_181),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_86),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_25),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_182),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_169),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_57),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_80),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_48),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_88),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_105),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_219),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_194),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_20),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_41),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_66),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_47),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_81),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_2),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_225),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_201),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_35),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_139),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_187),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_251),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_296),
.Y(n_386)
);

OAI22x1_ASAP7_75t_L g387 ( 
.A1(n_235),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_296),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

OAI22x1_ASAP7_75t_R g390 ( 
.A1(n_322),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_296),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_296),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_326),
.B(n_5),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_280),
.B(n_7),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_302),
.B(n_7),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_319),
.B(n_8),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_236),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_326),
.B(n_8),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_311),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_239),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_9),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_312),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_240),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_10),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_254),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_312),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_299),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_281),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_266),
.B(n_11),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_271),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_254),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_312),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_300),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_281),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_293),
.Y(n_418)
);

BUFx12f_ASAP7_75t_L g419 ( 
.A(n_292),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_306),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_348),
.B(n_12),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_358),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_234),
.B(n_15),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_304),
.B(n_16),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_237),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_295),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_238),
.Y(n_428)
);

OAI22x1_ASAP7_75t_R g429 ( 
.A1(n_364),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_292),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_310),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_374),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_337),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_310),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_382),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_368),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_232),
.Y(n_438)
);

BUFx8_ASAP7_75t_SL g439 ( 
.A(n_379),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_255),
.Y(n_440)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_337),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_255),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_383),
.B(n_22),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_337),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_324),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_327),
.B(n_23),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_284),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_290),
.B(n_23),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_255),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

BUFx8_ASAP7_75t_SL g452 ( 
.A(n_336),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_255),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_243),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_244),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_246),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_307),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_247),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_255),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_233),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_250),
.B(n_24),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_245),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_290),
.B(n_25),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_252),
.B(n_26),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_253),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_257),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_258),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_325),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_469)
);

XNOR2x1_ASAP7_75t_L g470 ( 
.A(n_357),
.B(n_359),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_366),
.B(n_29),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_259),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_264),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_265),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_248),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_267),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_372),
.B(n_30),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g479 ( 
.A1(n_273),
.A2(n_31),
.B(n_32),
.Y(n_479)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_314),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_274),
.B(n_33),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_276),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_278),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_279),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_283),
.Y(n_485)
);

BUFx12f_ASAP7_75t_L g486 ( 
.A(n_249),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_285),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_242),
.Y(n_488)
);

INVx6_ASAP7_75t_L g489 ( 
.A(n_346),
.Y(n_489)
);

BUFx12f_ASAP7_75t_L g490 ( 
.A(n_256),
.Y(n_490)
);

NAND2x1p5_ASAP7_75t_L g491 ( 
.A(n_262),
.B(n_55),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_298),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_301),
.B(n_34),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_351),
.Y(n_494)
);

AOI22x1_ASAP7_75t_SL g495 ( 
.A1(n_351),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_303),
.B(n_37),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_355),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_305),
.B(n_40),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_308),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_355),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_316),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_317),
.B(n_43),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_318),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_320),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_260),
.Y(n_506)
);

CKINVDCx8_ASAP7_75t_R g507 ( 
.A(n_261),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_452),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_388),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_426),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_428),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_476),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_486),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_388),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_394),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_418),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_490),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_R g518 ( 
.A(n_507),
.B(n_269),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_439),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_463),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_488),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_R g522 ( 
.A(n_406),
.B(n_44),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_461),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_506),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_494),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_419),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_494),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_475),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_400),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_497),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_480),
.B(n_323),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_497),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_405),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_399),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_405),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_503),
.Y(n_537)
);

BUFx10_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_503),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_448),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_385),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g542 ( 
.A(n_448),
.B(n_331),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_406),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_413),
.B(n_270),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_415),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_427),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_386),
.B(n_332),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_412),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_458),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_R g551 ( 
.A(n_430),
.B(n_263),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_489),
.A2(n_478),
.B1(n_471),
.B2(n_396),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_411),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_417),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_431),
.B(n_435),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_R g559 ( 
.A(n_434),
.B(n_268),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_385),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_437),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_501),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_472),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_473),
.Y(n_564)
);

INVxp33_ASAP7_75t_SL g565 ( 
.A(n_395),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_477),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_501),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_446),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_390),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_451),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_451),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_409),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_404),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_453),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_453),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_485),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_456),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_457),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_457),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_565),
.B(n_421),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_516),
.B(n_552),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_541),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_541),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_549),
.B(n_464),
.C(n_449),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_572),
.B(n_386),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_557),
.B(n_421),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_516),
.B(n_424),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_521),
.B(n_391),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_536),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_558),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_510),
.B(n_425),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_511),
.B(n_444),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_579),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_569),
.B(n_496),
.C(n_493),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_512),
.B(n_444),
.Y(n_595)
);

AO221x1_ASAP7_75t_L g596 ( 
.A1(n_521),
.A2(n_387),
.B1(n_340),
.B2(n_341),
.C(n_339),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_523),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_538),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_391),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_547),
.B(n_392),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_514),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_568),
.B(n_502),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_531),
.B(n_392),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_538),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_571),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_514),
.B(n_392),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_509),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_520),
.B(n_397),
.Y(n_608)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_543),
.B(n_469),
.C(n_500),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g610 ( 
.A(n_562),
.B(n_402),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_514),
.B(n_402),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_515),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_556),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_529),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_524),
.B(n_398),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_563),
.B(n_441),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_564),
.B(n_441),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_535),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_570),
.B(n_407),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

BUFx5_ASAP7_75t_L g622 ( 
.A(n_566),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_574),
.B(n_447),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_575),
.B(n_462),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_554),
.B(n_465),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_551),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_545),
.Y(n_627)
);

BUFx5_ASAP7_75t_L g628 ( 
.A(n_576),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_567),
.B(n_465),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_553),
.B(n_481),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_577),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_518),
.B(n_555),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_560),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_540),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_542),
.B(n_498),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_546),
.B(n_275),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_559),
.B(n_438),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_532),
.B(n_438),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_573),
.B(n_443),
.Y(n_639)
);

BUFx5_ASAP7_75t_L g640 ( 
.A(n_522),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_550),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_596),
.A2(n_479),
.B1(n_548),
.B2(n_345),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_640),
.B(n_513),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_640),
.B(n_517),
.Y(n_644)
);

AND2x6_ASAP7_75t_SL g645 ( 
.A(n_581),
.B(n_429),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_580),
.B(n_533),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_601),
.Y(n_647)
);

AO22x1_ASAP7_75t_L g648 ( 
.A1(n_584),
.A2(n_539),
.B1(n_347),
.B2(n_349),
.Y(n_648)
);

OR2x2_ASAP7_75t_SL g649 ( 
.A(n_609),
.B(n_495),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_582),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_611),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_583),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_639),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_611),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_623),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_589),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_605),
.B(n_631),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_621),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_587),
.A2(n_334),
.B1(n_344),
.B2(n_272),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_597),
.A2(n_527),
.B1(n_530),
.B2(n_525),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_630),
.Y(n_661)
);

OR2x6_ASAP7_75t_L g662 ( 
.A(n_598),
.B(n_604),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_591),
.B(n_561),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_599),
.B(n_350),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_640),
.A2(n_479),
.B1(n_352),
.B2(n_353),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_627),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_592),
.B(n_537),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_595),
.B(n_526),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_637),
.B(n_354),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_590),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_633),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_519),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_608),
.B(n_508),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_611),
.Y(n_674)
);

NAND2x1_ASAP7_75t_L g675 ( 
.A(n_614),
.B(n_360),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_640),
.B(n_528),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_607),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_614),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_626),
.B(n_370),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_613),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_634),
.Y(n_681)
);

AND2x2_ASAP7_75t_SL g682 ( 
.A(n_594),
.B(n_495),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_616),
.B(n_491),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_615),
.B(n_423),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_625),
.B(n_277),
.Y(n_685)
);

NOR2x1p5_ASAP7_75t_L g686 ( 
.A(n_635),
.B(n_410),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_586),
.B(n_410),
.Y(n_687)
);

AND2x6_ASAP7_75t_L g688 ( 
.A(n_620),
.B(n_408),
.Y(n_688)
);

NOR2x1p5_ASAP7_75t_L g689 ( 
.A(n_593),
.B(n_416),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_455),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_628),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_619),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_632),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_629),
.B(n_282),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_624),
.B(n_416),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_628),
.B(n_466),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_641),
.B(n_468),
.C(n_466),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_606),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_610),
.B(n_286),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_612),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_628),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_588),
.B(n_287),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_617),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_618),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_691),
.A2(n_602),
.B(n_585),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_651),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_646),
.B(n_653),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_665),
.A2(n_422),
.B1(n_432),
.B2(n_420),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_661),
.B(n_636),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_651),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_687),
.A2(n_440),
.B1(n_442),
.B2(n_414),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_SL g712 ( 
.A(n_660),
.B(n_667),
.C(n_679),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_651),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_672),
.B(n_288),
.Y(n_714)
);

OAI21x1_ASAP7_75t_L g715 ( 
.A1(n_691),
.A2(n_600),
.B(n_603),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_683),
.B(n_289),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_701),
.B(n_450),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_674),
.A2(n_460),
.B(n_454),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_657),
.B(n_420),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_659),
.A2(n_367),
.B(n_294),
.C(n_297),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_692),
.B(n_291),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_649),
.A2(n_422),
.B1(n_432),
.B2(n_436),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_647),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_693),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_668),
.B(n_309),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_669),
.B(n_313),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_650),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_662),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_652),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_677),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_686),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_673),
.Y(n_732)
);

AOI21x1_ASAP7_75t_L g733 ( 
.A1(n_690),
.A2(n_393),
.B(n_389),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_655),
.B(n_695),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_663),
.B(n_389),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_643),
.B(n_328),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_644),
.B(n_329),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_681),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_703),
.B(n_330),
.Y(n_739)
);

AOI21x1_ASAP7_75t_L g740 ( 
.A1(n_696),
.A2(n_335),
.B(n_333),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_695),
.B(n_338),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_645),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_684),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_671),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_703),
.B(n_343),
.Y(n_745)
);

INVx3_ASAP7_75t_SL g746 ( 
.A(n_682),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_684),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_689),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_704),
.B(n_356),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_697),
.B(n_459),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_704),
.B(n_361),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_664),
.A2(n_381),
.B(n_365),
.C(n_369),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_694),
.B(n_362),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_676),
.B(n_373),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_642),
.B(n_378),
.C(n_377),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_656),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_710),
.B(n_654),
.Y(n_757)
);

OAI21x1_ASAP7_75t_L g758 ( 
.A1(n_715),
.A2(n_647),
.B(n_675),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_755),
.A2(n_688),
.B(n_685),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_730),
.Y(n_760)
);

BUFx12f_ASAP7_75t_L g761 ( 
.A(n_724),
.Y(n_761)
);

BUFx2_ASAP7_75t_SL g762 ( 
.A(n_738),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_744),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_707),
.B(n_648),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_732),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_728),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_743),
.B(n_698),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_727),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_710),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_723),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_747),
.B(n_698),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_717),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_705),
.A2(n_670),
.B(n_680),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_729),
.B(n_698),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_717),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_733),
.A2(n_666),
.B(n_658),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_756),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_725),
.B(n_714),
.Y(n_778)
);

CKINVDCx16_ASAP7_75t_R g779 ( 
.A(n_719),
.Y(n_779)
);

AO21x2_ASAP7_75t_L g780 ( 
.A1(n_740),
.A2(n_699),
.B(n_702),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_719),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_748),
.Y(n_782)
);

BUFx2_ASAP7_75t_SL g783 ( 
.A(n_734),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_735),
.B(n_700),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_718),
.A2(n_700),
.B(n_678),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_746),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_709),
.A2(n_678),
.B(n_59),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_717),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_750),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_731),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_712),
.B(n_706),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_713),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_742),
.Y(n_793)
);

BUFx2_ASAP7_75t_SL g794 ( 
.A(n_722),
.Y(n_794)
);

AND2x2_ASAP7_75t_SL g795 ( 
.A(n_736),
.B(n_459),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_752),
.A2(n_146),
.B(n_61),
.Y(n_796)
);

NAND2x1p5_ASAP7_75t_L g797 ( 
.A(n_711),
.B(n_467),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_739),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_711),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_721),
.B(n_722),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_745),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_741),
.B(n_474),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_749),
.A2(n_147),
.B(n_63),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_708),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_751),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_726),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_760),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_778),
.A2(n_708),
.B1(n_716),
.B2(n_753),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_759),
.A2(n_754),
.B(n_737),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_763),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_800),
.A2(n_505),
.B1(n_482),
.B2(n_483),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_763),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_777),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_788),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_794),
.A2(n_764),
.B1(n_795),
.B2(n_804),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_795),
.A2(n_720),
.B1(n_474),
.B2(n_492),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_SL g817 ( 
.A1(n_764),
.A2(n_492),
.B1(n_505),
.B2(n_504),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_790),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_784),
.B(n_482),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_757),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_758),
.A2(n_142),
.B(n_68),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_765),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_799),
.A2(n_504),
.B1(n_499),
.B2(n_487),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_798),
.A2(n_499),
.B1(n_487),
.B2(n_484),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_766),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_768),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_805),
.A2(n_46),
.B1(n_77),
.B2(n_78),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_792),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_773),
.Y(n_829)
);

CKINVDCx11_ASAP7_75t_R g830 ( 
.A(n_761),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_766),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_805),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_774),
.B(n_85),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_767),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_770),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_779),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_781),
.Y(n_838)
);

BUFx6f_ASAP7_75t_SL g839 ( 
.A(n_793),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_771),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_762),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_765),
.Y(n_842)
);

BUFx12f_ASAP7_75t_L g843 ( 
.A(n_761),
.Y(n_843)
);

CKINVDCx16_ASAP7_75t_R g844 ( 
.A(n_786),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_SL g845 ( 
.A1(n_783),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_807),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_815),
.B(n_801),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_815),
.B(n_806),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_809),
.A2(n_791),
.B1(n_806),
.B2(n_771),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_834),
.B(n_791),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_819),
.B(n_789),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_826),
.B(n_789),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_808),
.A2(n_802),
.B(n_796),
.C(n_789),
.Y(n_853)
);

OAI21x1_ASAP7_75t_L g854 ( 
.A1(n_821),
.A2(n_787),
.B(n_776),
.Y(n_854)
);

CKINVDCx14_ASAP7_75t_R g855 ( 
.A(n_830),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_834),
.B(n_797),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_SL g857 ( 
.A(n_844),
.B(n_793),
.C(n_782),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_818),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_842),
.B(n_769),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_822),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_811),
.A2(n_788),
.B1(n_757),
.B2(n_775),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_813),
.Y(n_862)
);

BUFx2_ASAP7_75t_SL g863 ( 
.A(n_839),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_828),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_843),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_837),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_816),
.A2(n_827),
.B1(n_817),
.B2(n_838),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_R g868 ( 
.A(n_812),
.B(n_772),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_835),
.B(n_780),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_841),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_840),
.B(n_803),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_836),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_817),
.A2(n_785),
.B1(n_95),
.B2(n_96),
.Y(n_873)
);

INVx4_ASAP7_75t_SL g874 ( 
.A(n_820),
.Y(n_874)
);

CKINVDCx11_ASAP7_75t_R g875 ( 
.A(n_825),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_820),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_814),
.B(n_223),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_810),
.Y(n_878)
);

BUFx12f_ASAP7_75t_L g879 ( 
.A(n_831),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_869),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_864),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_870),
.B(n_823),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_862),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_846),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_850),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_R g886 ( 
.A(n_857),
.B(n_814),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_856),
.Y(n_887)
);

AO21x2_ASAP7_75t_L g888 ( 
.A1(n_853),
.A2(n_829),
.B(n_832),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_848),
.B(n_847),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_850),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_852),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_848),
.B(n_833),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_871),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_847),
.B(n_845),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_859),
.B(n_824),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_872),
.B(n_824),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_879),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_858),
.B(n_845),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_866),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_854),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_878),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_849),
.B(n_103),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_849),
.B(n_851),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_876),
.B(n_867),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_860),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_856),
.B(n_110),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_877),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_889),
.B(n_863),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_885),
.B(n_874),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_898),
.B(n_861),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_891),
.B(n_873),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_885),
.B(n_865),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_884),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_891),
.B(n_875),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_880),
.B(n_868),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_883),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_880),
.B(n_855),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_890),
.B(n_112),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_881),
.B(n_121),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_893),
.B(n_125),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_887),
.B(n_126),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_893),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_907),
.B(n_131),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_887),
.B(n_132),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_922),
.B(n_887),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_914),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_908),
.B(n_903),
.Y(n_927)
);

NAND4xp25_ASAP7_75t_L g928 ( 
.A(n_910),
.B(n_882),
.C(n_901),
.D(n_904),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_917),
.B(n_899),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_912),
.B(n_894),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_916),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_910),
.A2(n_892),
.B1(n_902),
.B2(n_895),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_913),
.B(n_900),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_911),
.A2(n_902),
.B1(n_896),
.B2(n_897),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_921),
.B(n_886),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_928),
.B(n_915),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_932),
.A2(n_887),
.B1(n_906),
.B2(n_924),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_932),
.A2(n_921),
.B(n_924),
.C(n_920),
.Y(n_938)
);

NOR3xp33_ASAP7_75t_L g939 ( 
.A(n_929),
.B(n_923),
.C(n_919),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_938),
.A2(n_934),
.B1(n_926),
.B2(n_927),
.Y(n_940)
);

XNOR2xp5_ASAP7_75t_L g941 ( 
.A(n_939),
.B(n_905),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_SL g942 ( 
.A1(n_937),
.A2(n_930),
.B(n_925),
.Y(n_942)
);

AOI31xp33_ASAP7_75t_L g943 ( 
.A1(n_936),
.A2(n_935),
.A3(n_909),
.B(n_918),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_SL g944 ( 
.A1(n_942),
.A2(n_943),
.B(n_941),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_940),
.B(n_931),
.Y(n_945)
);

NOR3x1_ASAP7_75t_L g946 ( 
.A(n_944),
.B(n_935),
.C(n_933),
.Y(n_946)
);

NOR2x1p5_ASAP7_75t_SL g947 ( 
.A(n_946),
.B(n_945),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_947),
.Y(n_948)
);

NOR2x1_ASAP7_75t_L g949 ( 
.A(n_948),
.B(n_888),
.Y(n_949)
);

NAND4xp75_ASAP7_75t_L g950 ( 
.A(n_949),
.B(n_134),
.C(n_135),
.D(n_138),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_950),
.Y(n_951)
);

XNOR2xp5_ASAP7_75t_L g952 ( 
.A(n_951),
.B(n_155),
.Y(n_952)
);

AOI31xp33_ASAP7_75t_L g953 ( 
.A1(n_952),
.A2(n_156),
.A3(n_157),
.B(n_158),
.Y(n_953)
);

AOI31xp33_ASAP7_75t_L g954 ( 
.A1(n_952),
.A2(n_164),
.A3(n_167),
.B(n_168),
.Y(n_954)
);

OAI22x1_ASAP7_75t_L g955 ( 
.A1(n_953),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_954),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_956),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_955),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_958),
.Y(n_959)
);

AOI31xp67_ASAP7_75t_L g960 ( 
.A1(n_957),
.A2(n_179),
.A3(n_184),
.B(n_185),
.Y(n_960)
);

OAI321xp33_ASAP7_75t_L g961 ( 
.A1(n_959),
.A2(n_188),
.A3(n_190),
.B1(n_191),
.B2(n_195),
.C(n_197),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_960),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_961),
.B(n_210),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_SL g964 ( 
.A1(n_963),
.A2(n_962),
.B1(n_211),
.B2(n_212),
.Y(n_964)
);


endmodule