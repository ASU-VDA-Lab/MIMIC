module fake_jpeg_28775_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_15),
.B(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_59),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_82),
.Y(n_83)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_55),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_90),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_46),
.B(n_57),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_93),
.B(n_94),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_25),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_46),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_70),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_56),
.B(n_45),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_56),
.B(n_49),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_48),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_30),
.C(n_43),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_28),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_106),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_47),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_114),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_117),
.B1(n_99),
.B2(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_0),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_113),
.C(n_115),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_26),
.B(n_41),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_18),
.B(n_36),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_24),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_31),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR4xp25_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_23),
.C(n_40),
.D(n_39),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_127),
.B(n_130),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_19),
.C(n_38),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_129),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_108),
.B(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_114),
.B(n_33),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_136),
.B1(n_119),
.B2(n_126),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_124),
.B1(n_122),
.B2(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_137),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_135),
.B(n_131),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_139),
.B1(n_125),
.B2(n_14),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_13),
.B(n_32),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_35),
.Y(n_146)
);


endmodule