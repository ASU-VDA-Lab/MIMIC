module fake_jpeg_17599_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_24),
.B1(n_17),
.B2(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_49),
.B1(n_52),
.B2(n_61),
.Y(n_70)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_27),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_26),
.B1(n_29),
.B2(n_18),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_16),
.B(n_25),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_38),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_27),
.B(n_1),
.Y(n_51)
);

OR2x4_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_19),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_29),
.B1(n_20),
.B2(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_59),
.B1(n_33),
.B2(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_75),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_69),
.B(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_72),
.Y(n_84)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_78),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_61),
.B(n_53),
.C(n_49),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_40),
.B1(n_19),
.B2(n_28),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_83),
.B1(n_47),
.B2(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_73),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_34),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_34),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_79),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_55),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_53),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_89),
.B1(n_95),
.B2(n_98),
.Y(n_111)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_94),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_75),
.C(n_82),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_79),
.C(n_77),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_72),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_105),
.Y(n_122)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_60),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_16),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_62),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_54),
.B1(n_56),
.B2(n_44),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_54),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_66),
.B(n_70),
.C(n_73),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_128),
.B(n_85),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_60),
.C(n_34),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_91),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_56),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_127),
.B1(n_86),
.B2(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_106),
.B1(n_47),
.B2(n_84),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_84),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_113),
.B1(n_108),
.B2(n_120),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_30),
.B(n_22),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_134),
.C(n_146),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_94),
.B1(n_93),
.B2(n_102),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_147),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_93),
.B1(n_97),
.B2(n_87),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_93),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_97),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_122),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_125),
.Y(n_152)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_103),
.B1(n_80),
.B2(n_65),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_151),
.B1(n_156),
.B2(n_165),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_114),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_164),
.B1(n_139),
.B2(n_138),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_128),
.B1(n_111),
.B2(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_158),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_116),
.B1(n_119),
.B2(n_118),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_108),
.B(n_116),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_16),
.B(n_25),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_122),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_47),
.B1(n_112),
.B2(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_139),
.B1(n_117),
.B2(n_145),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_124),
.B1(n_54),
.B2(n_112),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_131),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_145),
.B1(n_140),
.B2(n_44),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_176),
.B1(n_181),
.B2(n_161),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_159),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_38),
.A3(n_35),
.B1(n_37),
.B2(n_36),
.C1(n_47),
.C2(n_30),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_30),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_162),
.C(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_149),
.B1(n_156),
.B2(n_165),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_155),
.CI(n_158),
.CON(n_182),
.SN(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_0),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_181),
.B(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_187),
.A2(n_170),
.B1(n_176),
.B2(n_167),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_0),
.C(n_1),
.Y(n_201)
);

NAND4xp25_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_22),
.C(n_38),
.D(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_14),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_201),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_187),
.A2(n_167),
.B1(n_180),
.B2(n_14),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_200),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_191),
.B1(n_189),
.B2(n_183),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_184),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_190),
.B(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_206),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_185),
.C(n_186),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_196),
.B(n_203),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_194),
.B1(n_202),
.B2(n_7),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_186),
.B(n_6),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_4),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_214),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.C(n_207),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_197),
.C(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_6),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_218),
.B(n_219),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_221),
.B(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_208),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_9),
.C(n_10),
.Y(n_226)
);

OAI21x1_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_216),
.B(n_8),
.Y(n_224)
);

AO21x2_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_7),
.B(n_8),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_226),
.B(n_222),
.C(n_10),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_225),
.B(n_11),
.C(n_12),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_9),
.Y(n_229)
);


endmodule