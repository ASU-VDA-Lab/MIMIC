module fake_jpeg_16492_n_354 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_0),
.CON(n_44),
.SN(n_44)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_50),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_12),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_58),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_66),
.Y(n_89)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_70),
.B(n_76),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_18),
.C(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_73),
.B(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_34),
.B1(n_26),
.B2(n_21),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_83),
.A2(n_101),
.B1(n_118),
.B2(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_14),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_26),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_43),
.B(n_21),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_106),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_20),
.B1(n_32),
.B2(n_2),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_29),
.B1(n_24),
.B2(n_18),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_103),
.A2(n_96),
.B1(n_105),
.B2(n_81),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_40),
.B(n_35),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_29),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_112),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_65),
.B(n_0),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_1),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_1),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_48),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_4),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_126),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_54),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_142),
.C(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_5),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_57),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_128),
.A2(n_164),
.B(n_165),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_60),
.B1(n_52),
.B2(n_57),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_134),
.B1(n_143),
.B2(n_147),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_130),
.B(n_132),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_69),
.B1(n_7),
.B2(n_8),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_71),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_146),
.Y(n_178)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_140),
.A2(n_141),
.B(n_148),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_84),
.A2(n_117),
.B1(n_102),
.B2(n_98),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_11),
.B1(n_7),
.B2(n_10),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_161),
.B1(n_158),
.B2(n_156),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_10),
.B1(n_11),
.B2(n_93),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_79),
.A2(n_10),
.B1(n_11),
.B2(n_92),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_10),
.B1(n_101),
.B2(n_74),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_102),
.A2(n_107),
.B1(n_72),
.B2(n_104),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_151),
.A2(n_158),
.B1(n_166),
.B2(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_80),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_162),
.Y(n_185)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_73),
.B(n_77),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_132),
.Y(n_187)
);

AOI22x1_ASAP7_75t_L g158 ( 
.A1(n_82),
.A2(n_80),
.B1(n_97),
.B2(n_100),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_72),
.A2(n_104),
.B1(n_115),
.B2(n_88),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_105),
.A2(n_81),
.B1(n_97),
.B2(n_100),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_82),
.A2(n_50),
.B1(n_84),
.B2(n_83),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_131),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_128),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_191),
.C(n_168),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_194),
.B1(n_171),
.B2(n_170),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_190),
.C(n_191),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_121),
.B1(n_155),
.B2(n_153),
.Y(n_216)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_133),
.C(n_126),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_137),
.C(n_136),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_204),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_130),
.B1(n_124),
.B2(n_154),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_135),
.C(n_149),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_200),
.Y(n_209)
);

NAND2x1_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_123),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_197),
.B(n_202),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_124),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_199),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_159),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_134),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_164),
.A2(n_141),
.B1(n_122),
.B2(n_144),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_165),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_153),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_170),
.A2(n_197),
.B1(n_202),
.B2(n_172),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_211),
.B(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_229),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_230),
.Y(n_262)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_225),
.B(n_235),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_197),
.B(n_205),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_204),
.B1(n_207),
.B2(n_186),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_228),
.B1(n_241),
.B2(n_211),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_207),
.A2(n_169),
.B1(n_195),
.B2(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_187),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_238),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_173),
.B(n_187),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_190),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_225),
.B(n_238),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_180),
.A2(n_182),
.B1(n_193),
.B2(n_188),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_184),
.C(n_198),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_267),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_227),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_245),
.B(n_254),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_182),
.B1(n_193),
.B2(n_179),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_247),
.A2(n_251),
.B1(n_270),
.B2(n_233),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_234),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_261),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_226),
.B1(n_215),
.B2(n_211),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_271),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_212),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_265),
.B1(n_266),
.B2(n_250),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_210),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_269),
.B(n_266),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_213),
.B1(n_236),
.B2(n_237),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_242),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_252),
.B(n_248),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_209),
.C(n_240),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_SL g269 ( 
.A(n_209),
.B(n_241),
.C(n_230),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_231),
.A2(n_208),
.B1(n_223),
.B2(n_232),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_273),
.A2(n_277),
.B(n_279),
.Y(n_308)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_275),
.B(n_286),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_268),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_249),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_246),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_285),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_283),
.B1(n_289),
.B2(n_292),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_269),
.B1(n_253),
.B2(n_251),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_263),
.A2(n_248),
.B1(n_258),
.B2(n_253),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_262),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_244),
.A2(n_268),
.B1(n_247),
.B2(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_243),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_294),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_260),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_260),
.B1(n_264),
.B2(n_256),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_295),
.Y(n_300)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_264),
.B1(n_271),
.B2(n_257),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_307),
.B(n_312),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_245),
.B(n_255),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_306),
.B(n_282),
.Y(n_319)
);

XOR2x2_ASAP7_75t_SL g306 ( 
.A(n_275),
.B(n_267),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_270),
.B(n_292),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_278),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_311),
.C(n_291),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_276),
.C(n_288),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_281),
.A2(n_273),
.B(n_279),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_274),
.A2(n_276),
.B1(n_287),
.B2(n_272),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_313),
.A2(n_272),
.B(n_293),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_304),
.B(n_289),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_275),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_318),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_321),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_324),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_325),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_294),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_280),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_290),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_299),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_329),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_317),
.A2(n_308),
.B(n_312),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_334),
.A2(n_302),
.B(n_306),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_307),
.B(n_308),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_327),
.B(n_325),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_296),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_338),
.A2(n_334),
.B1(n_305),
.B2(n_333),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_342),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_321),
.C(n_316),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_343),
.C(n_330),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_336),
.A2(n_305),
.B1(n_314),
.B2(n_326),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_345),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_331),
.C(n_332),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_346),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_348),
.B(n_298),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_350),
.A2(n_351),
.B(n_347),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_298),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_344),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_345),
.Y(n_354)
);


endmodule