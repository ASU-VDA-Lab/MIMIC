module real_aes_9880_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1873;
wire n_1313;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1893;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_355;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1800;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1855;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_719;
wire n_465;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1691;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1889;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1277;
wire n_1049;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_1851;
wire n_780;
wire n_931;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1891;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AO221x1_ASAP7_75t_L g1603 ( .A1(n_0), .A2(n_137), .B1(n_1558), .B2(n_1604), .C(n_1606), .Y(n_1603) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_1), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g1592 ( .A1(n_2), .A2(n_124), .B1(n_1558), .B2(n_1562), .Y(n_1592) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_3), .A2(n_303), .B1(n_577), .B2(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g658 ( .A(n_3), .Y(n_658) );
INVx1_ASAP7_75t_L g1820 ( .A(n_4), .Y(n_1820) );
INVx1_ASAP7_75t_L g1249 ( .A(n_5), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1855 ( .A1(n_6), .A2(n_97), .B1(n_753), .B2(n_756), .Y(n_1855) );
INVx1_ASAP7_75t_L g1888 ( .A(n_6), .Y(n_1888) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_7), .A2(n_206), .B1(n_433), .B2(n_437), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_7), .A2(n_206), .B1(n_473), .B2(n_475), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_8), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_9), .A2(n_198), .B1(n_634), .B2(n_712), .C(n_1066), .Y(n_1183) );
OAI22xp33_ASAP7_75t_L g1188 ( .A1(n_9), .A2(n_301), .B1(n_544), .B2(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1533 ( .A(n_10), .Y(n_1533) );
INVx1_ASAP7_75t_L g1060 ( .A(n_11), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_11), .A2(n_106), .B1(n_583), .B2(n_1077), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1310 ( .A1(n_12), .A2(n_31), .B1(n_1311), .B2(n_1312), .C(n_1314), .Y(n_1310) );
INVx1_ASAP7_75t_L g1373 ( .A(n_12), .Y(n_1373) );
OAI22xp33_ASAP7_75t_L g1462 ( .A1(n_13), .A2(n_95), .B1(n_614), .B2(n_643), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g1468 ( .A1(n_13), .A2(n_95), .B1(n_588), .B2(n_697), .C(n_1469), .Y(n_1468) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_14), .A2(n_258), .B1(n_770), .B2(n_1020), .C(n_1025), .Y(n_1229) );
OAI22xp33_ASAP7_75t_L g1235 ( .A1(n_14), .A2(n_104), .B1(n_867), .B2(n_870), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_15), .A2(n_113), .B1(n_705), .B2(n_1068), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g1074 ( .A1(n_15), .A2(n_113), .B1(n_988), .B2(n_1007), .Y(n_1074) );
INVx1_ASAP7_75t_L g819 ( .A(n_16), .Y(n_819) );
OAI211xp5_ASAP7_75t_SL g849 ( .A1(n_16), .A2(n_614), .B(n_850), .C(n_860), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g1799 ( .A(n_17), .Y(n_1799) );
INVx1_ASAP7_75t_L g1607 ( .A(n_18), .Y(n_1607) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_19), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_20), .A2(n_66), .B1(n_753), .B2(n_756), .Y(n_752) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_20), .A2(n_182), .B1(n_359), .B2(n_522), .Y(n_763) );
AO22x2_ASAP7_75t_L g371 ( .A1(n_21), .A2(n_372), .B1(n_524), .B2(n_525), .Y(n_371) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_21), .Y(n_524) );
INVx1_ASAP7_75t_L g1402 ( .A(n_22), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_22), .A2(n_117), .B1(n_481), .B2(n_484), .Y(n_1436) );
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_23), .A2(n_89), .B1(n_705), .B2(n_1070), .Y(n_1069) );
INVxp67_ASAP7_75t_SL g1091 ( .A(n_23), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_24), .A2(n_340), .B1(n_487), .B2(n_788), .Y(n_1153) );
INVxp67_ASAP7_75t_SL g1174 ( .A(n_24), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_25), .A2(n_131), .B1(n_1297), .B2(n_1298), .Y(n_1296) );
INVx1_ASAP7_75t_L g1341 ( .A(n_25), .Y(n_1341) );
INVx1_ASAP7_75t_L g747 ( .A(n_26), .Y(n_747) );
OAI222xp33_ASAP7_75t_L g760 ( .A1(n_26), .A2(n_227), .B1(n_313), .B2(n_506), .C1(n_761), .C2(n_762), .Y(n_760) );
OAI222xp33_ASAP7_75t_L g940 ( .A1(n_27), .A2(n_61), .B1(n_142), .B2(n_685), .C1(n_941), .C2(n_944), .Y(n_940) );
INVx1_ASAP7_75t_L g961 ( .A(n_27), .Y(n_961) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_28), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g1302 ( .A(n_29), .Y(n_1302) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_30), .A2(n_130), .B1(n_578), .B2(n_591), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_30), .A2(n_130), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g1369 ( .A(n_31), .Y(n_1369) );
INVx1_ASAP7_75t_L g681 ( .A(n_32), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_32), .A2(n_316), .B1(n_439), .B2(n_712), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g1854 ( .A(n_33), .B(n_751), .Y(n_1854) );
INVx1_ASAP7_75t_L g1886 ( .A(n_33), .Y(n_1886) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_34), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_35), .A2(n_152), .B1(n_592), .B2(n_725), .Y(n_999) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_35), .A2(n_152), .B1(n_451), .B2(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_36), .A2(n_248), .B1(n_444), .B2(n_449), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_36), .A2(n_248), .B1(n_479), .B2(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g350 ( .A(n_37), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_38), .A2(n_112), .B1(n_750), .B2(n_751), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_38), .A2(n_112), .B1(n_707), .B2(n_716), .Y(n_774) );
INVx1_ASAP7_75t_L g1252 ( .A(n_39), .Y(n_1252) );
OAI211xp5_ASAP7_75t_SL g1273 ( .A1(n_39), .A2(n_614), .B(n_1274), .C(n_1279), .Y(n_1273) );
AOI22xp5_ASAP7_75t_L g1557 ( .A1(n_40), .A2(n_143), .B1(n_1558), .B2(n_1562), .Y(n_1557) );
INVxp67_ASAP7_75t_SL g1061 ( .A(n_41), .Y(n_1061) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_41), .A2(n_175), .B1(n_685), .B2(n_941), .Y(n_1085) );
INVx1_ASAP7_75t_L g1098 ( .A(n_42), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_42), .A2(n_215), .B1(n_712), .B2(n_771), .Y(n_1127) );
INVx1_ASAP7_75t_L g765 ( .A(n_43), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_43), .A2(n_225), .B1(n_487), .B2(n_788), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_44), .A2(n_144), .B1(n_631), .B2(n_771), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_44), .A2(n_144), .B1(n_695), .B2(n_697), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_45), .A2(n_236), .B1(n_583), .B2(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g650 ( .A(n_45), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g1413 ( .A(n_46), .Y(n_1413) );
AOI22x1_ASAP7_75t_SL g738 ( .A1(n_47), .A2(n_739), .B1(n_789), .B2(n_790), .Y(n_738) );
INVx1_ASAP7_75t_L g789 ( .A(n_47), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g1794 ( .A1(n_48), .A2(n_339), .B1(n_1432), .B2(n_1793), .Y(n_1794) );
OAI22xp33_ASAP7_75t_L g1827 ( .A1(n_48), .A2(n_318), .B1(n_643), .B2(n_665), .Y(n_1827) );
INVx1_ASAP7_75t_L g1509 ( .A(n_49), .Y(n_1509) );
INVx1_ASAP7_75t_L g1285 ( .A(n_50), .Y(n_1285) );
XNOR2xp5_ASAP7_75t_L g793 ( .A(n_51), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g1207 ( .A(n_52), .Y(n_1207) );
OAI221xp5_ASAP7_75t_L g1215 ( .A1(n_52), .A2(n_643), .B1(n_848), .B2(n_1216), .C(n_1220), .Y(n_1215) );
INVx1_ASAP7_75t_L g888 ( .A(n_53), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_53), .A2(n_614), .B1(n_909), .B2(n_917), .C(n_923), .Y(n_908) );
AO221x2_ASAP7_75t_L g1690 ( .A1(n_54), .A2(n_269), .B1(n_1604), .B2(n_1691), .C(n_1693), .Y(n_1690) );
OAI22xp33_ASAP7_75t_L g1259 ( .A1(n_55), .A2(n_235), .B1(n_537), .B2(n_544), .Y(n_1259) );
INVx1_ASAP7_75t_L g1277 ( .A(n_55), .Y(n_1277) );
INVx1_ASAP7_75t_L g1149 ( .A(n_56), .Y(n_1149) );
INVx1_ASAP7_75t_L g690 ( .A(n_57), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_57), .A2(n_179), .B1(n_705), .B2(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g968 ( .A(n_58), .Y(n_968) );
AOI22xp33_ASAP7_75t_SL g985 ( .A1(n_58), .A2(n_111), .B1(n_697), .B2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g1447 ( .A(n_59), .Y(n_1447) );
AOI221xp5_ASAP7_75t_L g1464 ( .A1(n_59), .A2(n_244), .B1(n_697), .B2(n_1465), .C(n_1467), .Y(n_1464) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_60), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g973 ( .A1(n_61), .A2(n_292), .B1(n_631), .B2(n_719), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_62), .A2(n_294), .B1(n_1558), .B2(n_1562), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_63), .A2(n_194), .B1(n_705), .B2(n_921), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_63), .A2(n_194), .B1(n_481), .B2(n_988), .Y(n_1129) );
AOI22xp5_ASAP7_75t_L g1591 ( .A1(n_64), .A2(n_321), .B1(n_1546), .B2(n_1554), .Y(n_1591) );
XOR2xp5_ASAP7_75t_L g1784 ( .A(n_64), .B(n_1785), .Y(n_1784) );
AOI22xp5_ASAP7_75t_L g1836 ( .A1(n_64), .A2(n_1837), .B1(n_1891), .B2(n_1894), .Y(n_1836) );
INVx1_ASAP7_75t_L g1818 ( .A(n_65), .Y(n_1818) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_66), .A2(n_140), .B1(n_433), .B2(n_771), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_67), .Y(n_880) );
INVxp33_ASAP7_75t_SL g1490 ( .A(n_68), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_68), .A2(n_332), .B1(n_1299), .B2(n_1522), .Y(n_1521) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_69), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_70), .A2(n_147), .B1(n_770), .B2(n_771), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_70), .A2(n_147), .B1(n_484), .B2(n_783), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g1321 ( .A(n_71), .Y(n_1321) );
OAI22xp33_ASAP7_75t_L g828 ( .A1(n_72), .A2(n_333), .B1(n_829), .B2(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g862 ( .A(n_72), .Y(n_862) );
AO22x1_ASAP7_75t_L g1568 ( .A1(n_73), .A2(n_253), .B1(n_1562), .B2(n_1569), .Y(n_1568) );
AOI22xp33_ASAP7_75t_L g1789 ( .A1(n_74), .A2(n_300), .B1(n_1311), .B2(n_1790), .Y(n_1789) );
INVx1_ASAP7_75t_L g1806 ( .A(n_74), .Y(n_1806) );
INVx1_ASAP7_75t_L g912 ( .A(n_75), .Y(n_912) );
OAI22xp33_ASAP7_75t_L g928 ( .A1(n_75), .A2(n_167), .B1(n_537), .B2(n_544), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g1303 ( .A1(n_76), .A2(n_239), .B1(n_1304), .B2(n_1307), .Y(n_1303) );
OAI221xp5_ASAP7_75t_L g1352 ( .A1(n_76), .A2(n_239), .B1(n_1353), .B2(n_1357), .C(n_1360), .Y(n_1352) );
INVx1_ASAP7_75t_L g1256 ( .A(n_77), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_77), .A2(n_224), .B1(n_836), .B2(n_837), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_78), .A2(n_334), .B1(n_584), .B2(n_588), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_78), .A2(n_643), .B1(n_645), .B2(n_657), .C(n_662), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_79), .Y(n_1419) );
AO22x1_ASAP7_75t_L g1570 ( .A1(n_80), .A2(n_252), .B1(n_1546), .B2(n_1554), .Y(n_1570) );
INVx1_ASAP7_75t_L g1099 ( .A(n_81), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_81), .A2(n_165), .B1(n_705), .B2(n_1126), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_82), .A2(n_245), .B1(n_481), .B2(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g513 ( .A(n_82), .Y(n_513) );
INVxp67_ASAP7_75t_SL g1499 ( .A(n_83), .Y(n_1499) );
AOI221xp5_ASAP7_75t_L g1527 ( .A1(n_83), .A2(n_335), .B1(n_1528), .B2(n_1529), .C(n_1530), .Y(n_1527) );
INVx1_ASAP7_75t_L g403 ( .A(n_84), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_84), .A2(n_193), .B1(n_503), .B2(n_506), .Y(n_502) );
INVx1_ASAP7_75t_L g826 ( .A(n_85), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_85), .A2(n_284), .B1(n_836), .B2(n_837), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g1142 ( .A(n_86), .Y(n_1142) );
XNOR2x2_ASAP7_75t_L g1439 ( .A(n_87), .B(n_1440), .Y(n_1439) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_88), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_88), .A2(n_250), .B1(n_988), .B2(n_1080), .Y(n_1079) );
INVxp33_ASAP7_75t_L g1090 ( .A(n_89), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g1456 ( .A(n_90), .Y(n_1456) );
BUFx2_ASAP7_75t_L g425 ( .A(n_91), .Y(n_425) );
INVx1_ASAP7_75t_L g462 ( .A(n_91), .Y(n_462) );
BUFx2_ASAP7_75t_L g490 ( .A(n_91), .Y(n_490) );
OR2x2_ASAP7_75t_L g1336 ( .A(n_91), .B(n_610), .Y(n_1336) );
AOI22xp33_ASAP7_75t_SL g773 ( .A1(n_92), .A2(n_231), .B1(n_444), .B2(n_707), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_92), .A2(n_231), .B1(n_778), .B2(n_780), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g1417 ( .A(n_93), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_94), .A2(n_328), .B1(n_695), .B2(n_697), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_94), .A2(n_328), .B1(n_712), .B2(n_719), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g1391 ( .A(n_96), .Y(n_1391) );
INVx1_ASAP7_75t_L g1850 ( .A(n_97), .Y(n_1850) );
INVx1_ASAP7_75t_L g918 ( .A(n_98), .Y(n_918) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_98), .A2(n_195), .B1(n_867), .B2(n_870), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_99), .A2(n_153), .B1(n_684), .B2(n_685), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_99), .A2(n_153), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_100), .Y(n_1445) );
INVx1_ASAP7_75t_L g550 ( .A(n_101), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_101), .A2(n_279), .B1(n_630), .B2(n_631), .C(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g891 ( .A(n_102), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_102), .A2(n_107), .B1(n_836), .B2(n_837), .Y(n_896) );
OAI221xp5_ASAP7_75t_L g1491 ( .A1(n_103), .A2(n_181), .B1(n_1353), .B2(n_1360), .C(n_1492), .Y(n_1491) );
OAI22xp5_ASAP7_75t_L g1524 ( .A1(n_103), .A2(n_181), .B1(n_1304), .B2(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1227 ( .A(n_104), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_105), .A2(n_203), .B1(n_712), .B2(n_1072), .Y(n_1071) );
INVxp67_ASAP7_75t_SL g1083 ( .A(n_105), .Y(n_1083) );
INVxp33_ASAP7_75t_L g1056 ( .A(n_106), .Y(n_1056) );
INVx1_ASAP7_75t_L g890 ( .A(n_107), .Y(n_890) );
AO221x1_ASAP7_75t_L g1024 ( .A1(n_108), .A2(n_199), .B1(n_434), .B2(n_720), .C(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1039 ( .A(n_108), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_109), .A2(n_263), .B1(n_484), .B2(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1375 ( .A(n_109), .Y(n_1375) );
INVx1_ASAP7_75t_L g956 ( .A(n_110), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_110), .A2(n_218), .B1(n_592), .B2(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g959 ( .A(n_111), .Y(n_959) );
AO221x1_ASAP7_75t_L g1575 ( .A1(n_114), .A2(n_126), .B1(n_1558), .B2(n_1562), .C(n_1576), .Y(n_1575) );
AO22x2_ASAP7_75t_L g935 ( .A1(n_115), .A2(n_936), .B1(n_937), .B2(n_991), .Y(n_935) );
INVxp67_ASAP7_75t_SL g936 ( .A(n_115), .Y(n_936) );
AO221x1_ASAP7_75t_L g1583 ( .A1(n_115), .A2(n_306), .B1(n_1558), .B2(n_1562), .C(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g1586 ( .A(n_116), .Y(n_1586) );
INVx1_ASAP7_75t_L g1407 ( .A(n_117), .Y(n_1407) );
INVx1_ASAP7_75t_L g1251 ( .A(n_118), .Y(n_1251) );
OAI221xp5_ASAP7_75t_L g1265 ( .A1(n_118), .A2(n_643), .B1(n_662), .B2(n_1266), .C(n_1269), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_119), .A2(n_273), .B1(n_695), .B2(n_1001), .Y(n_1000) );
AOI221xp5_ASAP7_75t_L g1019 ( .A1(n_119), .A2(n_273), .B1(n_770), .B2(n_1020), .C(n_1021), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_120), .A2(n_201), .B1(n_630), .B2(n_631), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_120), .A2(n_201), .B1(n_695), .B2(n_697), .Y(n_982) );
INVx1_ASAP7_75t_L g884 ( .A(n_121), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_122), .Y(n_1203) );
INVx1_ASAP7_75t_L g1580 ( .A(n_123), .Y(n_1580) );
AOI22xp5_ASAP7_75t_L g1545 ( .A1(n_125), .A2(n_148), .B1(n_1546), .B2(n_1554), .Y(n_1545) );
INVx1_ASAP7_75t_L g1180 ( .A(n_127), .Y(n_1180) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_127), .A2(n_198), .B1(n_867), .B2(n_870), .Y(n_1190) );
XNOR2xp5_ASAP7_75t_L g529 ( .A(n_128), .B(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_129), .A2(n_161), .B1(n_475), .B2(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g520 ( .A(n_129), .Y(n_520) );
INVx1_ASAP7_75t_L g1350 ( .A(n_131), .Y(n_1350) );
INVx1_ASAP7_75t_L g1158 ( .A(n_132), .Y(n_1158) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_132), .A2(n_643), .B1(n_662), .B2(n_1170), .C(n_1172), .Y(n_1169) );
INVx1_ASAP7_75t_L g1694 ( .A(n_133), .Y(n_1694) );
INVx1_ASAP7_75t_L g1114 ( .A(n_134), .Y(n_1114) );
AOI22xp33_ASAP7_75t_SL g1132 ( .A1(n_134), .A2(n_299), .B1(n_697), .B2(n_986), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_135), .A2(n_156), .B1(n_592), .B2(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g733 ( .A(n_135), .Y(n_733) );
CKINVDCx5p33_ASAP7_75t_R g1451 ( .A(n_136), .Y(n_1451) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_138), .A2(n_197), .B1(n_591), .B2(n_592), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_138), .A2(n_197), .B1(n_665), .B2(n_667), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_139), .Y(n_554) );
INVx1_ASAP7_75t_L g743 ( .A(n_140), .Y(n_743) );
CKINVDCx5p33_ASAP7_75t_R g1851 ( .A(n_141), .Y(n_1851) );
INVx1_ASAP7_75t_L g963 ( .A(n_142), .Y(n_963) );
XOR2xp5_ASAP7_75t_L g1480 ( .A(n_143), .B(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1550 ( .A(n_145), .Y(n_1550) );
OAI22xp33_ASAP7_75t_L g1212 ( .A1(n_146), .A2(n_317), .B1(n_829), .B2(n_831), .Y(n_1212) );
INVx1_ASAP7_75t_L g1231 ( .A(n_146), .Y(n_1231) );
INVx1_ASAP7_75t_L g1585 ( .A(n_149), .Y(n_1585) );
INVx1_ASAP7_75t_L g1109 ( .A(n_150), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_150), .A2(n_192), .B1(n_481), .B2(n_556), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_151), .A2(n_338), .B1(n_822), .B2(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1217 ( .A(n_151), .Y(n_1217) );
INVx1_ASAP7_75t_L g1057 ( .A(n_154), .Y(n_1057) );
INVx1_ASAP7_75t_L g1403 ( .A(n_155), .Y(n_1403) );
AOI221xp5_ASAP7_75t_L g1431 ( .A1(n_155), .A2(n_208), .B1(n_480), .B2(n_1432), .C(n_1434), .Y(n_1431) );
INVx1_ASAP7_75t_L g734 ( .A(n_156), .Y(n_734) );
INVx1_ASAP7_75t_L g1244 ( .A(n_157), .Y(n_1244) );
INVx1_ASAP7_75t_L g1551 ( .A(n_158), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_158), .B(n_1549), .Y(n_1556) );
INVx1_ASAP7_75t_L g1210 ( .A(n_159), .Y(n_1210) );
OAI211xp5_ASAP7_75t_SL g1224 ( .A1(n_159), .A2(n_614), .B(n_1225), .C(n_1230), .Y(n_1224) );
INVx1_ASAP7_75t_L g392 ( .A(n_160), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_160), .A2(n_185), .B1(n_454), .B2(n_457), .Y(n_453) );
INVx1_ASAP7_75t_L g495 ( .A(n_161), .Y(n_495) );
INVx1_ASAP7_75t_L g1393 ( .A(n_162), .Y(n_1393) );
AOI21xp33_ASAP7_75t_L g1428 ( .A1(n_162), .A2(n_1005), .B(n_1429), .Y(n_1428) );
INVx2_ASAP7_75t_L g362 ( .A(n_163), .Y(n_362) );
INVx1_ASAP7_75t_L g1394 ( .A(n_164), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_164), .A2(n_222), .B1(n_482), .B2(n_822), .Y(n_1427) );
INVx1_ASAP7_75t_L g1102 ( .A(n_165), .Y(n_1102) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_166), .A2(n_205), .B1(n_831), .B2(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1185 ( .A(n_166), .Y(n_1185) );
INVx1_ASAP7_75t_L g919 ( .A(n_167), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_168), .A2(n_260), .B1(n_716), .B2(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_168), .A2(n_260), .B1(n_577), .B2(n_592), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g1868 ( .A(n_169), .Y(n_1868) );
BUFx3_ASAP7_75t_L g382 ( .A(n_170), .Y(n_382) );
INVx1_ASAP7_75t_L g398 ( .A(n_170), .Y(n_398) );
INVx1_ASAP7_75t_L g1228 ( .A(n_171), .Y(n_1228) );
OAI22xp33_ASAP7_75t_L g1234 ( .A1(n_171), .A2(n_258), .B1(n_544), .B2(n_1189), .Y(n_1234) );
CKINVDCx5p33_ASAP7_75t_R g1860 ( .A(n_172), .Y(n_1860) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_173), .Y(n_1028) );
INVx1_ASAP7_75t_L g1815 ( .A(n_174), .Y(n_1815) );
INVx1_ASAP7_75t_L g1062 ( .A(n_175), .Y(n_1062) );
CKINVDCx5p33_ASAP7_75t_R g1852 ( .A(n_176), .Y(n_1852) );
INVxp33_ASAP7_75t_SL g1487 ( .A(n_177), .Y(n_1487) );
AOI221xp5_ASAP7_75t_L g1517 ( .A1(n_177), .A2(n_285), .B1(n_484), .B2(n_1432), .C(n_1518), .Y(n_1517) );
OAI22xp5_ASAP7_75t_L g1461 ( .A1(n_178), .A2(n_305), .B1(n_836), .B2(n_837), .Y(n_1461) );
INVx1_ASAP7_75t_L g1473 ( .A(n_178), .Y(n_1473) );
INVx1_ASAP7_75t_L g691 ( .A(n_179), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g1103 ( .A1(n_180), .A2(n_243), .B1(n_685), .B2(n_1104), .C(n_1105), .Y(n_1103) );
INVx1_ASAP7_75t_L g1112 ( .A(n_180), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_182), .A2(n_227), .B1(n_785), .B2(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g1160 ( .A(n_183), .Y(n_1160) );
OAI211xp5_ASAP7_75t_SL g1175 ( .A1(n_183), .A2(n_614), .B(n_1176), .C(n_1184), .Y(n_1175) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_184), .Y(n_1010) );
INVx1_ASAP7_75t_L g417 ( .A(n_185), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g1006 ( .A1(n_186), .A2(n_341), .B1(n_556), .B2(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1014 ( .A(n_186), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_187), .A2(n_200), .B1(n_1292), .B2(n_1293), .C(n_1294), .Y(n_1291) );
INVx1_ASAP7_75t_L g1348 ( .A(n_187), .Y(n_1348) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_188), .A2(n_342), .B1(n_439), .B2(n_634), .C(n_770), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g866 ( .A1(n_188), .A2(n_278), .B1(n_867), .B2(n_870), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1795 ( .A1(n_189), .A2(n_318), .B1(n_1163), .B2(n_1796), .Y(n_1795) );
OAI22xp33_ASAP7_75t_L g1803 ( .A1(n_189), .A2(n_339), .B1(n_614), .B2(n_667), .Y(n_1803) );
CKINVDCx5p33_ASAP7_75t_R g1801 ( .A(n_190), .Y(n_1801) );
INVx1_ASAP7_75t_L g1608 ( .A(n_191), .Y(n_1608) );
INVx1_ASAP7_75t_L g1110 ( .A(n_192), .Y(n_1110) );
INVx1_ASAP7_75t_L g409 ( .A(n_193), .Y(n_409) );
INVx1_ASAP7_75t_L g915 ( .A(n_195), .Y(n_915) );
INVx1_ASAP7_75t_L g1696 ( .A(n_196), .Y(n_1696) );
INVx1_ASAP7_75t_L g1041 ( .A(n_199), .Y(n_1041) );
INVx1_ASAP7_75t_L g1345 ( .A(n_200), .Y(n_1345) );
INVx1_ASAP7_75t_L g423 ( .A(n_202), .Y(n_423) );
INVx1_ASAP7_75t_L g541 ( .A(n_202), .Y(n_541) );
INVxp33_ASAP7_75t_L g1087 ( .A(n_203), .Y(n_1087) );
OAI22xp33_ASAP7_75t_L g1260 ( .A1(n_204), .A2(n_267), .B1(n_867), .B2(n_870), .Y(n_1260) );
AOI221xp5_ASAP7_75t_L g1278 ( .A1(n_204), .A2(n_235), .B1(n_1020), .B2(n_1025), .C(n_1223), .Y(n_1278) );
INVx1_ASAP7_75t_L g1186 ( .A(n_205), .Y(n_1186) );
CKINVDCx5p33_ASAP7_75t_R g1872 ( .A(n_207), .Y(n_1872) );
INVx1_ASAP7_75t_L g1405 ( .A(n_208), .Y(n_1405) );
INVx1_ASAP7_75t_L g1511 ( .A(n_209), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_210), .A2(n_312), .B1(n_697), .B2(n_1003), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1023 ( .A1(n_210), .A2(n_614), .B1(n_1024), .B2(n_1026), .C(n_1029), .Y(n_1023) );
INVx1_ASAP7_75t_L g818 ( .A(n_211), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g838 ( .A1(n_211), .A2(n_643), .B1(n_839), .B2(n_845), .C(n_848), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_212), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_213), .Y(n_385) );
INVx1_ASAP7_75t_L g1577 ( .A(n_214), .Y(n_1577) );
INVx1_ASAP7_75t_L g1106 ( .A(n_215), .Y(n_1106) );
INVxp67_ASAP7_75t_SL g1500 ( .A(n_216), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_216), .A2(n_287), .B1(n_785), .B2(n_788), .Y(n_1531) );
AOI22xp5_ASAP7_75t_L g1566 ( .A1(n_217), .A2(n_343), .B1(n_1546), .B2(n_1554), .Y(n_1566) );
INVx1_ASAP7_75t_L g955 ( .A(n_218), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g1460 ( .A(n_219), .Y(n_1460) );
OAI221xp5_ASAP7_75t_L g1474 ( .A1(n_219), .A2(n_562), .B1(n_571), .B2(n_596), .C(n_1475), .Y(n_1474) );
CKINVDCx5p33_ASAP7_75t_R g1411 ( .A(n_220), .Y(n_1411) );
INVx1_ASAP7_75t_L g894 ( .A(n_221), .Y(n_894) );
INVx1_ASAP7_75t_L g1389 ( .A(n_222), .Y(n_1389) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_223), .Y(n_1246) );
INVx1_ASAP7_75t_L g1254 ( .A(n_224), .Y(n_1254) );
INVx1_ASAP7_75t_L g766 ( .A(n_225), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g1821 ( .A(n_226), .Y(n_1821) );
CKINVDCx5p33_ASAP7_75t_R g1101 ( .A(n_228), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g892 ( .A1(n_229), .A2(n_311), .B1(n_829), .B2(n_831), .Y(n_892) );
INVx1_ASAP7_75t_L g926 ( .A(n_229), .Y(n_926) );
CKINVDCx16_ASAP7_75t_R g1049 ( .A(n_230), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1792 ( .A1(n_232), .A2(n_247), .B1(n_1432), .B2(n_1793), .Y(n_1792) );
INVx1_ASAP7_75t_L g1812 ( .A(n_232), .Y(n_1812) );
INVx1_ASAP7_75t_L g1198 ( .A(n_233), .Y(n_1198) );
INVx1_ASAP7_75t_L g887 ( .A(n_234), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_234), .A2(n_643), .B1(n_848), .B2(n_898), .C(n_904), .Y(n_897) );
INVx1_ASAP7_75t_L g654 ( .A(n_236), .Y(n_654) );
INVx1_ASAP7_75t_L g1242 ( .A(n_237), .Y(n_1242) );
INVx1_ASAP7_75t_L g413 ( .A(n_238), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_238), .A2(n_329), .B1(n_433), .B2(n_437), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_240), .Y(n_1453) );
OAI22xp5_ASAP7_75t_L g1843 ( .A1(n_241), .A2(n_264), .B1(n_1844), .B2(n_1846), .Y(n_1843) );
INVx1_ASAP7_75t_L g1878 ( .A(n_241), .Y(n_1878) );
INVx1_ASAP7_75t_L g1202 ( .A(n_242), .Y(n_1202) );
AOI21xp33_ASAP7_75t_L g1222 ( .A1(n_242), .A2(n_1021), .B(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1113 ( .A(n_243), .Y(n_1113) );
AOI21xp33_ASAP7_75t_L g1448 ( .A1(n_244), .A2(n_611), .B(n_1021), .Y(n_1448) );
INVx1_ASAP7_75t_L g517 ( .A(n_245), .Y(n_517) );
INVx1_ASAP7_75t_L g1332 ( .A(n_246), .Y(n_1332) );
INVx1_ASAP7_75t_L g1810 ( .A(n_247), .Y(n_1810) );
OAI211xp5_ASAP7_75t_L g1847 ( .A1(n_249), .A2(n_646), .B(n_969), .C(n_1848), .Y(n_1847) );
INVx1_ASAP7_75t_L g1875 ( .A(n_249), .Y(n_1875) );
INVx1_ASAP7_75t_L g1053 ( .A(n_250), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g1326 ( .A(n_251), .Y(n_1326) );
XNOR2xp5_ASAP7_75t_L g1195 ( .A(n_253), .B(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g878 ( .A(n_254), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g1211 ( .A1(n_255), .A2(n_280), .B1(n_804), .B2(n_1080), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_255), .A2(n_280), .B1(n_665), .B2(n_667), .Y(n_1214) );
BUFx3_ASAP7_75t_L g383 ( .A(n_256), .Y(n_383) );
INVx1_ASAP7_75t_L g420 ( .A(n_256), .Y(n_420) );
INVx1_ASAP7_75t_L g1262 ( .A(n_257), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_259), .Y(n_1009) );
AO22x2_ASAP7_75t_L g1094 ( .A1(n_261), .A2(n_1095), .B1(n_1134), .B2(n_1135), .Y(n_1094) );
INVxp67_ASAP7_75t_L g1134 ( .A(n_261), .Y(n_1134) );
XNOR2xp5_ASAP7_75t_L g1237 ( .A(n_262), .B(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1367 ( .A(n_263), .Y(n_1367) );
INVx1_ASAP7_75t_L g1877 ( .A(n_264), .Y(n_1877) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_265), .Y(n_358) );
INVx1_ASAP7_75t_L g466 ( .A(n_265), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_265), .B(n_320), .Y(n_610) );
AND2x2_ASAP7_75t_L g618 ( .A(n_265), .B(n_465), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_266), .Y(n_1027) );
INVx1_ASAP7_75t_L g1276 ( .A(n_267), .Y(n_1276) );
AOI21xp33_ASAP7_75t_L g1454 ( .A1(n_268), .A2(n_434), .B(n_1025), .Y(n_1454) );
INVx1_ASAP7_75t_L g1477 ( .A(n_268), .Y(n_1477) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_270), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g379 ( .A(n_271), .Y(n_379) );
OR2x2_ASAP7_75t_L g540 ( .A(n_271), .B(n_541), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g1329 ( .A(n_272), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_274), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_275), .Y(n_1444) );
CKINVDCx5p33_ASAP7_75t_R g1865 ( .A(n_276), .Y(n_1865) );
INVx1_ASAP7_75t_L g1506 ( .A(n_277), .Y(n_1506) );
INVx1_ASAP7_75t_L g854 ( .A(n_278), .Y(n_854) );
INVx1_ASAP7_75t_L g542 ( .A(n_279), .Y(n_542) );
INVx1_ASAP7_75t_L g858 ( .A(n_281), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g865 ( .A1(n_281), .A2(n_342), .B1(n_537), .B2(n_544), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g1450 ( .A(n_282), .Y(n_1450) );
INVx1_ASAP7_75t_L g1384 ( .A(n_283), .Y(n_1384) );
INVx1_ASAP7_75t_L g823 ( .A(n_284), .Y(n_823) );
INVxp33_ASAP7_75t_L g1489 ( .A(n_285), .Y(n_1489) );
INVx1_ASAP7_75t_L g951 ( .A(n_286), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_286), .A2(n_297), .B1(n_705), .B2(n_843), .Y(n_974) );
INVxp33_ASAP7_75t_L g1495 ( .A(n_287), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g1873 ( .A(n_288), .Y(n_1873) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_289), .A2(n_304), .B1(n_697), .B2(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g736 ( .A(n_289), .Y(n_736) );
AOI22x1_ASAP7_75t_L g993 ( .A1(n_290), .A2(n_994), .B1(n_995), .B2(n_1042), .Y(n_993) );
INVxp67_ASAP7_75t_SL g1042 ( .A(n_290), .Y(n_1042) );
XOR2xp5_ASAP7_75t_L g1838 ( .A(n_291), .B(n_1839), .Y(n_1838) );
INVx1_ASAP7_75t_L g947 ( .A(n_292), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g1161 ( .A1(n_293), .A2(n_322), .B1(n_1162), .B2(n_1163), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_293), .A2(n_322), .B1(n_836), .B2(n_837), .Y(n_1168) );
INVx1_ASAP7_75t_L g1139 ( .A(n_294), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_295), .A2(n_336), .B1(n_712), .B2(n_1066), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_295), .A2(n_336), .B1(n_402), .B2(n_695), .Y(n_1075) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_296), .Y(n_569) );
INVx1_ASAP7_75t_L g950 ( .A(n_297), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g1416 ( .A(n_298), .Y(n_1416) );
INVx1_ASAP7_75t_L g1119 ( .A(n_299), .Y(n_1119) );
INVx1_ASAP7_75t_L g1807 ( .A(n_300), .Y(n_1807) );
INVx1_ASAP7_75t_L g1182 ( .A(n_301), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g1257 ( .A1(n_302), .A2(n_327), .B1(n_829), .B2(n_831), .Y(n_1257) );
INVx1_ASAP7_75t_L g1281 ( .A(n_302), .Y(n_1281) );
INVx1_ASAP7_75t_L g660 ( .A(n_303), .Y(n_660) );
INVx1_ASAP7_75t_L g728 ( .A(n_304), .Y(n_728) );
INVx1_ASAP7_75t_L g1472 ( .A(n_305), .Y(n_1472) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_307), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_307), .B(n_350), .Y(n_1553) );
AND3x2_ASAP7_75t_L g1561 ( .A(n_307), .B(n_350), .C(n_1550), .Y(n_1561) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_308), .Y(n_833) );
INVx2_ASAP7_75t_L g363 ( .A(n_309), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_310), .Y(n_882) );
INVx1_ASAP7_75t_L g924 ( .A(n_311), .Y(n_924) );
INVx1_ASAP7_75t_L g1022 ( .A(n_312), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_313), .Y(n_746) );
XNOR2xp5_ASAP7_75t_L g872 ( .A(n_314), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g600 ( .A(n_315), .Y(n_600) );
INVx1_ASAP7_75t_L g687 ( .A(n_316), .Y(n_687) );
INVx1_ASAP7_75t_L g1232 ( .A(n_317), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1396 ( .A1(n_319), .A2(n_323), .B1(n_1353), .B2(n_1357), .C(n_1397), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g1422 ( .A1(n_319), .A2(n_323), .B1(n_1307), .B2(n_1423), .C(n_1425), .Y(n_1422) );
INVx1_ASAP7_75t_L g365 ( .A(n_320), .Y(n_365) );
INVx2_ASAP7_75t_L g465 ( .A(n_320), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g1842 ( .A(n_324), .Y(n_1842) );
INVx1_ASAP7_75t_L g1512 ( .A(n_325), .Y(n_1512) );
INVx1_ASAP7_75t_L g1824 ( .A(n_326), .Y(n_1824) );
INVx1_ASAP7_75t_L g1280 ( .A(n_327), .Y(n_1280) );
INVx1_ASAP7_75t_L g400 ( .A(n_329), .Y(n_400) );
INVx1_ASAP7_75t_L g1459 ( .A(n_330), .Y(n_1459) );
HB1xp67_ASAP7_75t_L g1475 ( .A(n_330), .Y(n_1475) );
OAI211xp5_ASAP7_75t_L g1856 ( .A1(n_331), .A2(n_748), .B(n_1857), .C(n_1858), .Y(n_1856) );
INVx1_ASAP7_75t_L g1889 ( .A(n_331), .Y(n_1889) );
INVxp33_ASAP7_75t_SL g1485 ( .A(n_332), .Y(n_1485) );
INVx1_ASAP7_75t_L g861 ( .A(n_333), .Y(n_861) );
OAI211xp5_ASAP7_75t_SL g613 ( .A1(n_334), .A2(n_614), .B(n_619), .C(n_636), .Y(n_613) );
INVxp33_ASAP7_75t_SL g1496 ( .A(n_335), .Y(n_1496) );
INVx1_ASAP7_75t_L g1148 ( .A(n_337), .Y(n_1148) );
INVx1_ASAP7_75t_L g1219 ( .A(n_338), .Y(n_1219) );
INVxp33_ASAP7_75t_SL g1173 ( .A(n_340), .Y(n_1173) );
INVx1_ASAP7_75t_L g1015 ( .A(n_341), .Y(n_1015) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_366), .B(n_1537), .Y(n_344) );
INVx3_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_353), .Y(n_347) );
AND2x4_ASAP7_75t_L g1835 ( .A(n_348), .B(n_354), .Y(n_1835) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_SL g1893 ( .A(n_349), .Y(n_1893) );
NAND2xp5_ASAP7_75t_L g1896 ( .A(n_349), .B(n_351), .Y(n_1896) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g1892 ( .A(n_351), .B(n_1893), .Y(n_1892) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_355), .B(n_359), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g523 ( .A(n_356), .B(n_490), .Y(n_523) );
OR2x6_ASAP7_75t_L g737 ( .A(n_356), .B(n_490), .Y(n_737) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g431 ( .A(n_357), .B(n_365), .Y(n_431) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_358), .B(n_512), .Y(n_1021) );
INVx8_ASAP7_75t_L g519 ( .A(n_359), .Y(n_519) );
OR2x6_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
OR2x6_ASAP7_75t_L g522 ( .A(n_360), .B(n_511), .Y(n_522) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_360), .Y(n_653) );
INVx2_ASAP7_75t_SL g907 ( .A(n_360), .Y(n_907) );
INVx1_ASAP7_75t_L g914 ( .A(n_360), .Y(n_914) );
BUFx2_ASAP7_75t_L g1272 ( .A(n_360), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_360), .B(n_1336), .Y(n_1335) );
INVx2_ASAP7_75t_SL g1401 ( .A(n_360), .Y(n_1401) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g436 ( .A(n_362), .B(n_363), .Y(n_436) );
INVx1_ASAP7_75t_L g441 ( .A(n_362), .Y(n_441) );
INVx2_ASAP7_75t_L g446 ( .A(n_362), .Y(n_446) );
AND2x4_ASAP7_75t_L g452 ( .A(n_362), .B(n_442), .Y(n_452) );
INVx1_ASAP7_75t_L g508 ( .A(n_362), .Y(n_508) );
INVx2_ASAP7_75t_L g442 ( .A(n_363), .Y(n_442) );
INVx1_ASAP7_75t_L g448 ( .A(n_363), .Y(n_448) );
INVx1_ASAP7_75t_L g505 ( .A(n_363), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_363), .B(n_446), .Y(n_623) );
INVx1_ASAP7_75t_L g649 ( .A(n_363), .Y(n_649) );
AND2x4_ASAP7_75t_L g504 ( .A(n_364), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g506 ( .A(n_365), .B(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g731 ( .A(n_365), .B(n_507), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_1381), .B2(n_1536), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
XNOR2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_1043), .Y(n_368) );
XNOR2x1_ASAP7_75t_L g369 ( .A(n_370), .B(n_674), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_526), .B1(n_672), .B2(n_673), .Y(n_370) );
INVx2_ASAP7_75t_L g672 ( .A(n_371), .Y(n_672) );
INVx1_ASAP7_75t_L g525 ( .A(n_372), .Y(n_525) );
AOI211x1_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_421), .B(n_426), .C(n_493), .Y(n_372) );
NAND4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_384), .C(n_399), .D(n_412), .Y(n_373) );
INVx5_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_375), .A2(n_681), .B(n_682), .C(n_683), .Y(n_680) );
CKINVDCx8_ASAP7_75t_R g748 ( .A(n_375), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_375), .B(n_940), .Y(n_939) );
AOI211xp5_ASAP7_75t_L g1082 ( .A1(n_375), .A2(n_1083), .B(n_1084), .C(n_1085), .Y(n_1082) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
OAI21xp33_ASAP7_75t_L g1105 ( .A1(n_376), .A2(n_477), .B(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x6_ASAP7_75t_L g418 ( .A(n_377), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g754 ( .A(n_377), .Y(n_754) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_377), .B(n_402), .Y(n_1084) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x6_ASAP7_75t_L g410 ( .A(n_378), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_379), .Y(n_388) );
INVx1_ASAP7_75t_L g395 ( .A(n_379), .Y(n_395) );
AND2x2_ASAP7_75t_L g471 ( .A(n_379), .B(n_423), .Y(n_471) );
INVx2_ASAP7_75t_L g492 ( .A(n_379), .Y(n_492) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_380), .Y(n_402) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_380), .Y(n_477) );
INVx2_ASAP7_75t_L g698 ( .A(n_380), .Y(n_698) );
INVx1_ASAP7_75t_L g799 ( .A(n_380), .Y(n_799) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_381), .Y(n_586) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx2_ASAP7_75t_L g390 ( .A(n_382), .Y(n_390) );
AND2x4_ASAP7_75t_L g419 ( .A(n_382), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g391 ( .A(n_383), .Y(n_391) );
AND2x4_ASAP7_75t_L g397 ( .A(n_383), .B(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_392), .B2(n_393), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_385), .A2(n_519), .B1(n_520), .B2(n_521), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_386), .A2(n_414), .B1(n_687), .B2(n_688), .Y(n_686) );
INVx4_ASAP7_75t_L g756 ( .A(n_386), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_386), .A2(n_414), .B1(n_947), .B2(n_948), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_386), .A2(n_1057), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_386), .A2(n_418), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1100) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
AND2x4_ASAP7_75t_L g405 ( .A(n_387), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_SL g1861 ( .A(n_387), .B(n_406), .Y(n_1861) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx6_ASAP7_75t_L g416 ( .A(n_389), .Y(n_416) );
INVx2_ASAP7_75t_L g485 ( .A(n_389), .Y(n_485) );
BUFx2_ASAP7_75t_L g583 ( .A(n_389), .Y(n_583) );
AND2x2_ASAP7_75t_L g603 ( .A(n_389), .B(n_567), .Y(n_603) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g411 ( .A(n_390), .Y(n_411) );
INVx1_ASAP7_75t_L g408 ( .A(n_391), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_393), .A2(n_418), .B1(n_690), .B2(n_691), .Y(n_689) );
INVx4_ASAP7_75t_L g751 ( .A(n_393), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_393), .A2(n_418), .B1(n_950), .B2(n_951), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_393), .A2(n_418), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_393), .A2(n_414), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AND2x6_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
AND2x4_ASAP7_75t_L g414 ( .A(n_394), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_394), .B(n_415), .Y(n_1088) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g942 ( .A(n_395), .B(n_943), .Y(n_942) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_396), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g1080 ( .A(n_396), .Y(n_1080) );
INVx2_ASAP7_75t_L g1164 ( .A(n_396), .Y(n_1164) );
BUFx6f_ASAP7_75t_L g1205 ( .A(n_396), .Y(n_1205) );
INVx1_ASAP7_75t_L g1879 ( .A(n_396), .Y(n_1879) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_397), .Y(n_482) );
INVx1_ASAP7_75t_L g538 ( .A(n_397), .Y(n_538) );
INVx2_ASAP7_75t_L g581 ( .A(n_397), .Y(n_581) );
INVx1_ASAP7_75t_L g781 ( .A(n_397), .Y(n_781) );
INVx1_ASAP7_75t_L g547 ( .A(n_398), .Y(n_547) );
AOI222xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_403), .B2(n_404), .C1(n_409), .C2(n_410), .Y(n_399) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_402), .Y(n_682) );
BUFx4f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g684 ( .A(n_405), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_405), .A2(n_410), .B1(n_746), .B2(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g943 ( .A(n_407), .Y(n_943) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g564 ( .A(n_408), .Y(n_564) );
INVx3_ASAP7_75t_L g685 ( .A(n_410), .Y(n_685) );
AOI322xp5_ASAP7_75t_L g1858 ( .A1(n_410), .A2(n_1471), .A3(n_1851), .B1(n_1852), .B2(n_1859), .C1(n_1860), .C2(n_1861), .Y(n_1858) );
BUFx3_ASAP7_75t_L g573 ( .A(n_411), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_417), .B2(n_418), .Y(n_412) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_416), .Y(n_589) );
INVx2_ASAP7_75t_L g696 ( .A(n_416), .Y(n_696) );
INVx1_ASAP7_75t_L g986 ( .A(n_416), .Y(n_986) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_416), .Y(n_1005) );
HB1xp67_ASAP7_75t_L g1466 ( .A(n_416), .Y(n_1466) );
CKINVDCx6p67_ASAP7_75t_R g750 ( .A(n_418), .Y(n_750) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_419), .Y(n_480) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_419), .Y(n_488) );
INVx2_ASAP7_75t_SL g557 ( .A(n_419), .Y(n_557) );
BUFx2_ASAP7_75t_L g577 ( .A(n_419), .Y(n_577) );
BUFx3_ASAP7_75t_L g804 ( .A(n_419), .Y(n_804) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_419), .Y(n_822) );
BUFx2_ASAP7_75t_L g988 ( .A(n_419), .Y(n_988) );
BUFx6f_ASAP7_75t_L g1471 ( .A(n_419), .Y(n_1471) );
INVx1_ASAP7_75t_L g548 ( .A(n_420), .Y(n_548) );
AO211x2_ASAP7_75t_L g678 ( .A1(n_421), .A2(n_679), .B(n_692), .C(n_726), .Y(n_678) );
BUFx6f_ASAP7_75t_L g952 ( .A(n_421), .Y(n_952) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
AND2x4_ASAP7_75t_L g757 ( .A(n_422), .B(n_424), .Y(n_757) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g491 ( .A(n_423), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g1037 ( .A(n_424), .Y(n_1037) );
BUFx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g430 ( .A(n_425), .Y(n_430) );
OR2x6_ASAP7_75t_L g1365 ( .A(n_425), .B(n_1021), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_467), .Y(n_426) );
AOI33xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_432), .A3(n_443), .B1(n_453), .B2(n_458), .B3(n_459), .Y(n_427) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_429), .B(n_715), .C(n_718), .Y(n_714) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
OR2x6_ASAP7_75t_L g469 ( .A(n_430), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g605 ( .A(n_430), .Y(n_605) );
BUFx2_ASAP7_75t_L g671 ( .A(n_430), .Y(n_671) );
OR2x2_ASAP7_75t_L g701 ( .A(n_430), .B(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g768 ( .A(n_430), .B(n_431), .Y(n_768) );
OR2x2_ASAP7_75t_L g801 ( .A(n_430), .B(n_470), .Y(n_801) );
INVx1_ASAP7_75t_L g656 ( .A(n_431), .Y(n_656) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g611 ( .A(n_435), .Y(n_611) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_435), .Y(n_1223) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_436), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g727 ( .A1(n_437), .A2(n_499), .B(n_728), .C(n_729), .Y(n_727) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g960 ( .A(n_438), .Y(n_960) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g1066 ( .A(n_439), .Y(n_1066) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g498 ( .A(n_440), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_440), .B(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_440), .Y(n_720) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_440), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1117 ( .A(n_440), .Y(n_1117) );
AND2x4_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_445), .Y(n_456) );
AND2x4_ASAP7_75t_L g510 ( .A(n_445), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g666 ( .A(n_445), .B(n_618), .Y(n_666) );
INVx1_ASAP7_75t_L g706 ( .A(n_445), .Y(n_706) );
BUFx2_ASAP7_75t_L g716 ( .A(n_445), .Y(n_716) );
BUFx6f_ASAP7_75t_L g1018 ( .A(n_445), .Y(n_1018) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g641 ( .A(n_446), .Y(n_641) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_450), .A2(n_659), .B1(n_1173), .B2(n_1174), .Y(n_1172) );
OAI221xp5_ASAP7_75t_L g1225 ( .A1(n_450), .A2(n_1226), .B1(n_1227), .B2(n_1228), .C(n_1229), .Y(n_1225) );
OAI221xp5_ASAP7_75t_L g1274 ( .A1(n_450), .A2(n_1275), .B1(n_1276), .B2(n_1277), .C(n_1278), .Y(n_1274) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_450), .A2(n_1302), .B1(n_1329), .B2(n_1371), .Y(n_1376) );
INVx4_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g457 ( .A(n_451), .Y(n_457) );
INVx2_ASAP7_75t_SL g1374 ( .A(n_451), .Y(n_1374) );
INVx2_ASAP7_75t_SL g1808 ( .A(n_451), .Y(n_1808) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g516 ( .A(n_452), .Y(n_516) );
INVx1_ASAP7_75t_L g628 ( .A(n_452), .Y(n_628) );
INVx3_ASAP7_75t_L g710 ( .A(n_452), .Y(n_710) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_456), .B(n_1344), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_456), .B(n_1344), .Y(n_1395) );
INVx1_ASAP7_75t_L g1412 ( .A(n_457), .Y(n_1412) );
AOI33xp33_ASAP7_75t_L g767 ( .A1(n_459), .A2(n_768), .A3(n_769), .B1(n_773), .B2(n_774), .B3(n_775), .Y(n_767) );
AOI33xp33_ASAP7_75t_L g1064 ( .A1(n_459), .A2(n_768), .A3(n_1065), .B1(n_1067), .B2(n_1069), .B3(n_1071), .Y(n_1064) );
INVx2_ASAP7_75t_L g1890 ( .A(n_459), .Y(n_1890) );
INVx6_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx5_ASAP7_75t_L g713 ( .A(n_460), .Y(n_713) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_461), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g539 ( .A(n_462), .B(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g1344 ( .A(n_462), .B(n_618), .Y(n_1344) );
INVx2_ASAP7_75t_L g635 ( .A(n_463), .Y(n_635) );
BUFx2_ASAP7_75t_L g1025 ( .A(n_463), .Y(n_1025) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g501 ( .A(n_464), .Y(n_501) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g512 ( .A(n_465), .Y(n_512) );
AOI33xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_472), .A3(n_478), .B1(n_483), .B2(n_486), .B3(n_489), .Y(n_467) );
AOI33xp33_ASAP7_75t_L g776 ( .A1(n_468), .A2(n_489), .A3(n_777), .B1(n_782), .B2(n_784), .B3(n_787), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g575 ( .A(n_469), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g1145 ( .A1(n_469), .A2(n_1146), .B1(n_1154), .B2(n_1156), .Y(n_1145) );
CKINVDCx5p33_ASAP7_75t_R g1788 ( .A(n_469), .Y(n_1788) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g702 ( .A(n_471), .Y(n_702) );
INVx2_ASAP7_75t_SL g1316 ( .A(n_471), .Y(n_1316) );
BUFx3_ASAP7_75t_L g1435 ( .A(n_471), .Y(n_1435) );
INVx1_ASAP7_75t_L g1530 ( .A(n_471), .Y(n_1530) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_474), .Y(n_785) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_477), .Y(n_786) );
INVx1_ASAP7_75t_L g1313 ( .A(n_477), .Y(n_1313) );
AND2x4_ASAP7_75t_L g1322 ( .A(n_477), .B(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1433 ( .A(n_477), .Y(n_1433) );
BUFx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_SL g779 ( .A(n_480), .Y(n_779) );
AND2x4_ASAP7_75t_L g1300 ( .A(n_480), .B(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1523 ( .A(n_480), .Y(n_1523) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g879 ( .A(n_482), .Y(n_879) );
INVx1_ASAP7_75t_L g1243 ( .A(n_482), .Y(n_1243) );
BUFx3_ASAP7_75t_L g1318 ( .A(n_482), .Y(n_1318) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g552 ( .A(n_485), .Y(n_552) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx4f_ASAP7_75t_L g591 ( .A(n_488), .Y(n_591) );
INVx1_ASAP7_75t_L g871 ( .A(n_488), .Y(n_871) );
INVx4_ASAP7_75t_L g827 ( .A(n_489), .Y(n_827) );
BUFx4f_ASAP7_75t_L g1155 ( .A(n_489), .Y(n_1155) );
AOI221xp5_ASAP7_75t_L g1463 ( .A1(n_489), .A2(n_575), .B1(n_1464), .B2(n_1468), .C(n_1474), .Y(n_1463) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x4_ASAP7_75t_L g593 ( .A(n_490), .B(n_491), .Y(n_593) );
AND2x4_ASAP7_75t_L g602 ( .A(n_490), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g1295 ( .A(n_491), .Y(n_1295) );
CKINVDCx5p33_ASAP7_75t_R g1429 ( .A(n_491), .Y(n_1429) );
INVx2_ASAP7_75t_SL g1520 ( .A(n_491), .Y(n_1520) );
AND2x4_ASAP7_75t_L g567 ( .A(n_492), .B(n_568), .Y(n_567) );
AOI31xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_509), .A3(n_518), .B(n_523), .Y(n_493) );
AOI211xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_499), .C(n_502), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g630 ( .A(n_497), .Y(n_630) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g615 ( .A(n_498), .B(n_616), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g759 ( .A(n_499), .B(n_760), .C(n_763), .Y(n_759) );
CKINVDCx11_ASAP7_75t_R g969 ( .A(n_499), .Y(n_969) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_L g966 ( .A(n_501), .Y(n_966) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g730 ( .A(n_504), .Y(n_730) );
INVx2_ASAP7_75t_L g761 ( .A(n_504), .Y(n_761) );
AOI222xp33_ASAP7_75t_L g1111 ( .A1(n_504), .A2(n_964), .B1(n_1112), .B2(n_1113), .C1(n_1114), .C2(n_1115), .Y(n_1111) );
AOI322xp5_ASAP7_75t_L g1848 ( .A1(n_504), .A2(n_964), .A3(n_1845), .B1(n_1849), .B2(n_1850), .C1(n_1851), .C2(n_1852), .Y(n_1848) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_505), .Y(n_638) );
INVx1_ASAP7_75t_L g1034 ( .A(n_505), .Y(n_1034) );
AOI22xp5_ASAP7_75t_L g1458 ( .A1(n_505), .A2(n_1359), .B1(n_1459), .B2(n_1460), .Y(n_1458) );
INVx1_ASAP7_75t_L g965 ( .A(n_507), .Y(n_965) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g648 ( .A(n_508), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_508), .B(n_649), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_513), .B1(n_514), .B2(n_517), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_510), .A2(n_514), .B1(n_733), .B2(n_734), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_510), .A2(n_514), .B1(n_765), .B2(n_766), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_510), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_510), .A2(n_957), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_510), .A2(n_957), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
AND2x4_ASAP7_75t_L g514 ( .A(n_511), .B(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g957 ( .A(n_511), .B(n_515), .Y(n_957) );
INVx1_ASAP7_75t_L g1845 ( .A(n_511), .Y(n_1845) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx5_ASAP7_75t_SL g1846 ( .A(n_514), .Y(n_1846) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_516), .Y(n_661) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_519), .A2(n_521), .B1(n_688), .B2(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_519), .A2(n_521), .B1(n_948), .B2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_519), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_519), .A2(n_1058), .B1(n_1101), .B2(n_1119), .Y(n_1118) );
AOI211xp5_ASAP7_75t_L g1841 ( .A1(n_519), .A2(n_1842), .B(n_1843), .C(n_1847), .Y(n_1841) );
INVx5_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx4_ASAP7_75t_L g1058 ( .A(n_522), .Y(n_1058) );
OAI211xp5_ASAP7_75t_L g1840 ( .A1(n_523), .A2(n_1841), .B(n_1853), .C(n_1862), .Y(n_1840) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g673 ( .A(n_529), .Y(n_673) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_599), .C(n_612), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_558), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_549), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_542), .B2(n_543), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_535), .A2(n_554), .B1(n_620), .B2(n_624), .C(n_629), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g1038 ( .A1(n_536), .A2(n_551), .B1(n_602), .B2(n_1027), .C1(n_1030), .C2(n_1039), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_536), .A2(n_543), .B1(n_1451), .B2(n_1453), .Y(n_1478) );
AOI222xp33_ASAP7_75t_L g1828 ( .A1(n_536), .A2(n_551), .B1(n_602), .B2(n_1818), .C1(n_1821), .C2(n_1824), .Y(n_1828) );
CKINVDCx6p67_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_538), .A2(n_803), .B1(n_890), .B2(n_891), .Y(n_889) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_538), .B(n_539), .Y(n_1189) );
INVx2_ASAP7_75t_L g1791 ( .A(n_538), .Y(n_1791) );
OR2x6_ASAP7_75t_L g544 ( .A(n_539), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g553 ( .A(n_539), .Y(n_553) );
OR2x2_ASAP7_75t_L g867 ( .A(n_539), .B(n_868), .Y(n_867) );
OR2x2_ASAP7_75t_L g870 ( .A(n_539), .B(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g1301 ( .A(n_540), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_540), .B(n_755), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_540), .B(n_581), .Y(n_1331) );
INVx1_ASAP7_75t_L g568 ( .A(n_541), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_543), .A2(n_555), .B1(n_1028), .B2(n_1041), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1829 ( .A1(n_543), .A2(n_555), .B1(n_1815), .B2(n_1820), .Y(n_1829) );
CKINVDCx6p67_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g815 ( .A1(n_545), .A2(n_816), .B1(n_818), .B2(n_819), .Y(n_815) );
BUFx3_ASAP7_75t_L g883 ( .A(n_545), .Y(n_883) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g813 ( .A(n_546), .Y(n_813) );
BUFx4f_ASAP7_75t_L g1152 ( .A(n_546), .Y(n_1152) );
INVx1_ASAP7_75t_L g1209 ( .A(n_546), .Y(n_1209) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
OR2x2_ASAP7_75t_L g755 ( .A(n_547), .B(n_548), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B1(n_554), .B2(n_555), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g1476 ( .A1(n_551), .A2(n_555), .B1(n_602), .B2(n_1450), .C1(n_1456), .C2(n_1477), .Y(n_1476) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
BUFx2_ASAP7_75t_L g1793 ( .A(n_552), .Y(n_1793) );
AND2x2_ASAP7_75t_L g555 ( .A(n_553), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g725 ( .A(n_557), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g1876 ( .A1(n_557), .A2(n_1877), .B1(n_1878), .B2(n_1879), .Y(n_1876) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_574), .C(n_594), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_569), .B2(n_570), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_560), .A2(n_569), .B1(n_637), .B2(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g1166 ( .A(n_561), .Y(n_1166) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g830 ( .A(n_562), .Y(n_830) );
INVx1_ASAP7_75t_L g1800 ( .A(n_562), .Y(n_1800) );
NAND2x1p5_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g1306 ( .A(n_564), .Y(n_1306) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OR2x6_ASAP7_75t_L g571 ( .A(n_566), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g598 ( .A(n_566), .Y(n_598) );
OR2x2_ASAP7_75t_L g831 ( .A(n_566), .B(n_572), .Y(n_831) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_567), .B(n_1306), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_567), .B(n_573), .Y(n_1308) );
INVx1_ASAP7_75t_L g1324 ( .A(n_567), .Y(n_1324) );
AND2x4_ASAP7_75t_L g1424 ( .A(n_567), .B(n_1306), .Y(n_1424) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_570), .A2(n_797), .B1(n_830), .B2(n_1009), .C(n_1010), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1798 ( .A1(n_570), .A2(n_797), .B1(n_1799), .B2(n_1800), .C(n_1801), .Y(n_1798) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g1525 ( .A(n_572), .B(n_1324), .Y(n_1525) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI33xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .A3(n_582), .B1(n_587), .B2(n_590), .B3(n_593), .Y(n_574) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g592 ( .A(n_579), .Y(n_592) );
INVx2_ASAP7_75t_SL g807 ( .A(n_579), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_579), .A2(n_1470), .B1(n_1472), .B2(n_1473), .Y(n_1469) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g1299 ( .A(n_580), .Y(n_1299) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g1870 ( .A(n_581), .Y(n_1870) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g744 ( .A(n_585), .Y(n_744) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_586), .Y(n_597) );
BUFx3_ASAP7_75t_L g783 ( .A(n_586), .Y(n_783) );
BUFx4f_ASAP7_75t_L g1001 ( .A(n_586), .Y(n_1001) );
INVx1_ASAP7_75t_L g1078 ( .A(n_586), .Y(n_1078) );
AND2x4_ASAP7_75t_L g1320 ( .A(n_586), .B(n_1301), .Y(n_1320) );
INVx4_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g723 ( .A(n_589), .Y(n_723) );
INVx1_ASAP7_75t_L g1293 ( .A(n_589), .Y(n_1293) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_593), .B(n_722), .C(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g990 ( .A(n_593), .Y(n_990) );
AOI33xp33_ASAP7_75t_L g997 ( .A1(n_593), .A2(n_998), .A3(n_999), .B1(n_1000), .B2(n_1002), .B3(n_1006), .Y(n_997) );
AOI33xp33_ASAP7_75t_L g1073 ( .A1(n_593), .A2(n_998), .A3(n_1074), .B1(n_1075), .B2(n_1076), .B3(n_1079), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g1131 ( .A(n_593), .B(n_1132), .C(n_1133), .Y(n_1131) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
BUFx2_ASAP7_75t_SL g1529 ( .A(n_597), .Y(n_1529) );
AND2x2_ASAP7_75t_L g797 ( .A(n_598), .B(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_601), .B(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_601), .B(n_894), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_601), .B(n_1142), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_601), .B(n_1198), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_601), .B(n_1262), .Y(n_1261) );
OR2x6_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx2_ASAP7_75t_L g1337 ( .A(n_602), .Y(n_1337) );
NOR2xp67_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx2_ASAP7_75t_L g863 ( .A(n_605), .Y(n_863) );
INVx1_ASAP7_75t_L g1823 ( .A(n_606), .Y(n_1823) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .Y(n_606) );
AND2x2_ASAP7_75t_L g637 ( .A(n_607), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g925 ( .A(n_607), .B(n_638), .Y(n_925) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x6_ASAP7_75t_L g640 ( .A(n_608), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g662 ( .A(n_608), .B(n_663), .Y(n_662) );
OR2x6_ASAP7_75t_L g848 ( .A(n_608), .B(n_663), .Y(n_848) );
INVx1_ASAP7_75t_L g1035 ( .A(n_608), .Y(n_1035) );
AOI21xp33_ASAP7_75t_L g1825 ( .A1(n_608), .A2(n_905), .B(n_1826), .Y(n_1825) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g712 ( .A(n_611), .Y(n_712) );
OAI31xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_642), .A3(n_664), .B(n_669), .Y(n_612) );
INVx8_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g668 ( .A(n_616), .B(n_627), .Y(n_668) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g644 ( .A(n_618), .B(n_633), .Y(n_644) );
BUFx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g659 ( .A(n_622), .Y(n_659) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_622), .Y(n_841) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g853 ( .A(n_623), .Y(n_853) );
INVx1_ASAP7_75t_L g901 ( .A(n_623), .Y(n_901) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g717 ( .A(n_626), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g1884 ( .A1(n_626), .A2(n_851), .B1(n_1865), .B2(n_1868), .Y(n_1884) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g1029 ( .A1(n_631), .A2(n_1030), .B(n_1031), .C(n_1035), .Y(n_1029) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g1849 ( .A(n_632), .Y(n_1849) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_633), .Y(n_770) );
INVx1_ASAP7_75t_L g916 ( .A(n_634), .Y(n_916) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_637), .A2(n_639), .B1(n_861), .B2(n_862), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g1184 ( .A1(n_637), .A2(n_639), .B1(n_1185), .B2(n_1186), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_637), .A2(n_639), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_639), .A2(n_924), .B1(n_925), .B2(n_926), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_639), .A2(n_925), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
CKINVDCx11_ASAP7_75t_R g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g1359 ( .A(n_641), .Y(n_1359) );
CKINVDCx6p67_ASAP7_75t_R g643 ( .A(n_644), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_644), .A2(n_1017), .B1(n_1019), .B2(n_1022), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B1(n_651), .B2(n_654), .C(n_655), .Y(n_645) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_646), .A2(n_1400), .B1(n_1402), .B2(n_1403), .Y(n_1399) );
OAI22xp33_ASAP7_75t_L g1414 ( .A1(n_646), .A2(n_1415), .B1(n_1416), .B2(n_1417), .Y(n_1414) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g1171 ( .A(n_647), .Y(n_1171) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g663 ( .A(n_648), .Y(n_663) );
INVx2_ASAP7_75t_L g762 ( .A(n_648), .Y(n_762) );
INVx3_ASAP7_75t_L g905 ( .A(n_648), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g1170 ( .A1(n_651), .A2(n_655), .B1(n_1148), .B2(n_1149), .C(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g845 ( .A1(n_653), .A2(n_655), .B1(n_811), .B2(n_814), .C(n_846), .Y(n_845) );
BUFx2_ASAP7_75t_L g1415 ( .A(n_653), .Y(n_1415) );
OAI22xp33_ASAP7_75t_L g1881 ( .A1(n_653), .A2(n_1872), .B1(n_1873), .B2(n_1882), .Y(n_1881) );
OAI22xp33_ASAP7_75t_L g1887 ( .A1(n_653), .A2(n_910), .B1(n_1888), .B2(n_1889), .Y(n_1887) );
OAI221xp5_ASAP7_75t_L g904 ( .A1(n_655), .A2(n_882), .B1(n_884), .B2(n_905), .C(n_906), .Y(n_904) );
OAI221xp5_ASAP7_75t_L g1269 ( .A1(n_655), .A2(n_905), .B1(n_1246), .B2(n_1249), .C(n_1270), .Y(n_1269) );
OAI221xp5_ASAP7_75t_L g1809 ( .A1(n_655), .A2(n_762), .B1(n_1810), .B2(n_1811), .C(n_1812), .Y(n_1809) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_659), .A2(n_708), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_659), .A2(n_922), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
OAI22xp5_ASAP7_75t_L g1449 ( .A1(n_659), .A2(n_708), .B1(n_1450), .B2(n_1451), .Y(n_1449) );
INVx1_ASAP7_75t_L g903 ( .A(n_661), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_663), .B(n_1458), .Y(n_1457) );
HB1xp67_ASAP7_75t_L g1497 ( .A(n_663), .Y(n_1497) );
INVx1_ASAP7_75t_L g1883 ( .A(n_663), .Y(n_1883) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx3_ASAP7_75t_L g836 ( .A(n_666), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_666), .A2(n_668), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx3_ASAP7_75t_L g837 ( .A(n_668), .Y(n_837) );
OAI31xp33_ASAP7_75t_L g895 ( .A1(n_669), .A2(n_896), .A3(n_897), .B(n_908), .Y(n_895) );
OAI31xp33_ASAP7_75t_L g1263 ( .A1(n_669), .A2(n_1264), .A3(n_1265), .B(n_1273), .Y(n_1263) );
AOI31xp33_ASAP7_75t_L g1420 ( .A1(n_669), .A2(n_1421), .A3(n_1430), .B(n_1437), .Y(n_1420) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
CKINVDCx8_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
XNOR2x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_931), .Y(n_674) );
XNOR2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_791), .Y(n_675) );
XNOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_738), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_686), .C(n_689), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g692 ( .A(n_693), .B(n_703), .C(n_714), .D(n_721), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_699), .C(n_700), .Y(n_693) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g981 ( .A(n_700), .B(n_982), .C(n_983), .Y(n_981) );
NAND3xp33_ASAP7_75t_L g1128 ( .A(n_700), .B(n_1129), .C(n_1130), .Y(n_1128) );
INVx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_711), .C(n_713), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g1068 ( .A(n_708), .Y(n_1068) );
INVx1_ASAP7_75t_L g1268 ( .A(n_708), .Y(n_1268) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g844 ( .A(n_709), .Y(n_844) );
INVx2_ASAP7_75t_L g922 ( .A(n_709), .Y(n_922) );
INVx1_ASAP7_75t_L g1503 ( .A(n_709), .Y(n_1503) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_710), .Y(n_857) );
INVx3_ASAP7_75t_L g979 ( .A(n_710), .Y(n_979) );
NAND3xp33_ASAP7_75t_L g972 ( .A(n_713), .B(n_973), .C(n_974), .Y(n_972) );
NAND3xp33_ASAP7_75t_L g1124 ( .A(n_713), .B(n_1125), .C(n_1127), .Y(n_1124) );
CKINVDCx8_ASAP7_75t_R g1379 ( .A(n_713), .Y(n_1379) );
INVx1_ASAP7_75t_L g1181 ( .A(n_717), .Y(n_1181) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_SL g772 ( .A(n_720), .Y(n_772) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_720), .Y(n_1072) );
AOI31xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_732), .A3(n_735), .B(n_737), .Y(n_726) );
INVx1_ASAP7_75t_L g962 ( .A(n_730), .Y(n_962) );
AO21x1_ASAP7_75t_SL g758 ( .A1(n_737), .A2(n_759), .B(n_764), .Y(n_758) );
CKINVDCx16_ASAP7_75t_R g970 ( .A(n_737), .Y(n_970) );
AND4x1_ASAP7_75t_L g739 ( .A(n_740), .B(n_758), .C(n_767), .D(n_776), .Y(n_739) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_740), .B(n_758), .C(n_767), .D(n_776), .Y(n_790) );
OAI31xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_749), .A3(n_752), .B(n_757), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_745), .C(n_748), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g1859 ( .A(n_754), .Y(n_1859) );
BUFx2_ASAP7_75t_L g810 ( .A(n_755), .Y(n_810) );
INVx1_ASAP7_75t_L g817 ( .A(n_755), .Y(n_817) );
INVx2_ASAP7_75t_L g869 ( .A(n_755), .Y(n_869) );
INVx1_ASAP7_75t_SL g1092 ( .A(n_757), .Y(n_1092) );
OAI31xp33_ASAP7_75t_SL g1853 ( .A1(n_757), .A2(n_1854), .A3(n_1855), .B(n_1856), .Y(n_1853) );
OAI21xp33_ASAP7_75t_L g1452 ( .A1(n_762), .A2(n_1453), .B(n_1454), .Y(n_1452) );
NAND3xp33_ASAP7_75t_L g975 ( .A(n_768), .B(n_976), .C(n_980), .Y(n_975) );
NAND3xp33_ASAP7_75t_L g1121 ( .A(n_768), .B(n_1122), .C(n_1123), .Y(n_1121) );
A2O1A1Ixp33_ASAP7_75t_L g1455 ( .A1(n_770), .A2(n_1035), .B(n_1456), .C(n_1457), .Y(n_1455) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g1253 ( .A1(n_779), .A2(n_1254), .B1(n_1255), .B2(n_1256), .Y(n_1253) );
INVx1_ASAP7_75t_L g1297 ( .A(n_779), .Y(n_1297) );
OAI22xp5_ASAP7_75t_L g1467 ( .A1(n_779), .A2(n_781), .B1(n_1444), .B2(n_1445), .Y(n_1467) );
INVx1_ASAP7_75t_L g1528 ( .A(n_779), .Y(n_1528) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g788 ( .A(n_781), .Y(n_788) );
INVx1_ASAP7_75t_L g825 ( .A(n_781), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_872), .B2(n_930), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND4x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_832), .C(n_834), .D(n_864), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_800), .C(n_828), .Y(n_795) );
NOR3xp33_ASAP7_75t_SL g874 ( .A(n_796), .B(n_875), .C(n_892), .Y(n_874) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_797), .Y(n_1144) );
NOR3xp33_ASAP7_75t_SL g1199 ( .A(n_797), .B(n_1200), .C(n_1212), .Y(n_1199) );
NOR3xp33_ASAP7_75t_SL g1239 ( .A(n_797), .B(n_1240), .C(n_1257), .Y(n_1239) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1292 ( .A(n_799), .Y(n_1292) );
OAI33xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .A3(n_809), .B1(n_815), .B2(n_820), .B3(n_827), .Y(n_800) );
OAI33xp33_ASAP7_75t_L g875 ( .A1(n_801), .A2(n_827), .A3(n_876), .B1(n_881), .B2(n_885), .B3(n_889), .Y(n_875) );
INVx1_ASAP7_75t_SL g998 ( .A(n_801), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_801), .A2(n_1154), .B1(n_1201), .B2(n_1206), .Y(n_1200) );
OAI33xp33_ASAP7_75t_L g1240 ( .A1(n_801), .A2(n_827), .A3(n_1241), .B1(n_1245), .B2(n_1250), .B3(n_1253), .Y(n_1240) );
OAI33xp33_ASAP7_75t_L g1863 ( .A1(n_801), .A2(n_827), .A3(n_1864), .B1(n_1871), .B2(n_1874), .B3(n_1876), .Y(n_1863) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_805), .B1(n_806), .B2(n_808), .Y(n_802) );
INVx2_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
BUFx3_ASAP7_75t_L g1162 ( .A(n_804), .Y(n_1162) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_805), .A2(n_808), .B1(n_840), .B2(n_842), .Y(n_839) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_814), .Y(n_809) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_810), .A2(n_882), .B1(n_883), .B2(n_884), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_810), .A2(n_1159), .B1(n_1202), .B2(n_1203), .C(n_1204), .Y(n_1201) );
OAI221xp5_ASAP7_75t_L g1206 ( .A1(n_810), .A2(n_1207), .B1(n_1208), .B2(n_1210), .C(n_1211), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g945 ( .A(n_813), .Y(n_945) );
BUFx2_ASAP7_75t_L g1147 ( .A(n_816), .Y(n_1147) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B1(n_824), .B2(n_826), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g877 ( .A(n_822), .Y(n_877) );
BUFx2_ASAP7_75t_L g1311 ( .A(n_822), .Y(n_1311) );
BUFx3_ASAP7_75t_L g1796 ( .A(n_822), .Y(n_1796) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g1797 ( .A(n_827), .Y(n_1797) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI31xp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_838), .A3(n_849), .B(n_863), .Y(n_834) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g911 ( .A(n_846), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_846), .B(n_1032), .Y(n_1031) );
BUFx3_ASAP7_75t_L g1221 ( .A(n_846), .Y(n_1221) );
OAI221xp5_ASAP7_75t_L g1819 ( .A1(n_846), .A2(n_913), .B1(n_916), .B2(n_1820), .C(n_1821), .Y(n_1819) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_854), .B1(n_855), .B2(n_858), .C(n_859), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
BUFx2_ASAP7_75t_L g1505 ( .A(n_853), .Y(n_1505) );
OR2x2_ASAP7_75t_L g1844 ( .A(n_853), .B(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g1126 ( .A(n_857), .Y(n_1126) );
INVx2_ASAP7_75t_SL g1409 ( .A(n_857), .Y(n_1409) );
INVx2_ASAP7_75t_L g1508 ( .A(n_857), .Y(n_1508) );
INVx2_ASAP7_75t_L g1817 ( .A(n_857), .Y(n_1817) );
OAI31xp33_ASAP7_75t_L g1167 ( .A1(n_863), .A2(n_1168), .A3(n_1169), .B(n_1175), .Y(n_1167) );
OAI31xp33_ASAP7_75t_L g1441 ( .A1(n_863), .A2(n_1442), .A3(n_1461), .B(n_1462), .Y(n_1441) );
INVx1_ASAP7_75t_L g1514 ( .A(n_863), .Y(n_1514) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g886 ( .A(n_869), .Y(n_886) );
INVx2_ASAP7_75t_L g1157 ( .A(n_869), .Y(n_1157) );
INVx1_ASAP7_75t_L g930 ( .A(n_872), .Y(n_930) );
AND4x1_ASAP7_75t_L g873 ( .A(n_874), .B(n_893), .C(n_895), .D(n_927), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_876) );
OAI22xp33_ASAP7_75t_L g1241 ( .A1(n_877), .A2(n_1242), .B1(n_1243), .B2(n_1244), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_878), .A2(n_880), .B1(n_899), .B2(n_902), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_883), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g1874 ( .A1(n_883), .A2(n_886), .B1(n_1842), .B2(n_1875), .Y(n_1874) );
OAI22xp33_ASAP7_75t_L g1245 ( .A1(n_886), .A2(n_1246), .B1(n_1247), .B2(n_1249), .Y(n_1245) );
OAI22xp33_ASAP7_75t_L g1250 ( .A1(n_886), .A2(n_1159), .B1(n_1251), .B2(n_1252), .Y(n_1250) );
OAI22xp33_ASAP7_75t_SL g1871 ( .A1(n_886), .A2(n_1208), .B1(n_1872), .B2(n_1873), .Y(n_1871) );
OAI22xp5_ASAP7_75t_SL g917 ( .A1(n_899), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_899), .A2(n_1217), .B1(n_1218), .B2(n_1219), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_899), .A2(n_1242), .B1(n_1244), .B2(n_1267), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1805 ( .A1(n_899), .A2(n_1806), .B1(n_1807), .B2(n_1808), .Y(n_1805) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx2_ASAP7_75t_L g1226 ( .A(n_900), .Y(n_1226) );
INVx2_ASAP7_75t_L g1275 ( .A(n_900), .Y(n_1275) );
INVx2_ASAP7_75t_SL g1814 ( .A(n_900), .Y(n_1814) );
BUFx3_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g1179 ( .A(n_901), .Y(n_1179) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g1446 ( .A1(n_905), .A2(n_1447), .B(n_1448), .Y(n_1446) );
BUFx2_ASAP7_75t_L g1378 ( .A(n_906), .Y(n_1378) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_912), .B1(n_913), .B2(n_915), .C(n_916), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g1510 ( .A1(n_910), .A2(n_1378), .B1(n_1511), .B2(n_1512), .Y(n_1510) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g1368 ( .A(n_911), .Y(n_1368) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_913), .A2(n_1367), .B1(n_1368), .B2(n_1369), .Y(n_1366) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_922), .Y(n_921) );
INVx2_ASAP7_75t_L g1070 ( .A(n_922), .Y(n_1070) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
OAI22x1_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_935), .B1(n_992), .B2(n_993), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g991 ( .A(n_937), .Y(n_991) );
AOI221x1_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_952), .B1(n_953), .B2(n_970), .C(n_971), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_946), .C(n_949), .Y(n_938) );
INVx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g1104 ( .A(n_942), .Y(n_1104) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
AOI221x1_ASAP7_75t_L g1095 ( .A1(n_952), .A2(n_970), .B1(n_1096), .B2(n_1107), .C(n_1120), .Y(n_1095) );
NAND4xp25_ASAP7_75t_SL g953 ( .A(n_954), .B(n_958), .C(n_967), .D(n_969), .Y(n_953) );
AOI222xp33_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_960), .B1(n_961), .B2(n_962), .C1(n_963), .C2(n_964), .Y(n_958) );
AOI222xp33_ASAP7_75t_L g1059 ( .A1(n_960), .A2(n_962), .B1(n_964), .B2(n_1060), .C1(n_1061), .C2(n_1062), .Y(n_1059) );
AND2x4_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g1032 ( .A1(n_965), .A2(n_1009), .B1(n_1010), .B2(n_1033), .Y(n_1032) );
NAND4xp25_ASAP7_75t_SL g1051 ( .A(n_969), .B(n_1052), .C(n_1055), .D(n_1059), .Y(n_1051) );
NAND4xp25_ASAP7_75t_SL g1107 ( .A(n_969), .B(n_1108), .C(n_1111), .D(n_1118), .Y(n_1107) );
AOI211xp5_ASAP7_75t_L g1050 ( .A1(n_970), .A2(n_1051), .B(n_1063), .C(n_1081), .Y(n_1050) );
NAND4xp25_ASAP7_75t_L g971 ( .A(n_972), .B(n_975), .C(n_981), .D(n_984), .Y(n_971) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
AND2x4_ASAP7_75t_L g1343 ( .A(n_979), .B(n_1344), .Y(n_1343) );
NAND3xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_987), .C(n_989), .Y(n_984) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx2_ASAP7_75t_SL g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
NAND4xp75_ASAP7_75t_L g995 ( .A(n_996), .B(n_1011), .C(n_1038), .D(n_1040), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_997), .B(n_1008), .Y(n_996) );
INVx2_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
OAI21xp5_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1023), .B(n_1036), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1016), .Y(n_1012) );
AND2x6_ASAP7_75t_L g1346 ( .A(n_1020), .B(n_1344), .Y(n_1346) );
NAND2x1p5_ASAP7_75t_L g1361 ( .A(n_1020), .B(n_1356), .Y(n_1361) );
NAND2x1_ASAP7_75t_SL g1355 ( .A(n_1033), .B(n_1356), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1826 ( .A1(n_1033), .A2(n_1359), .B1(n_1799), .B2(n_1801), .Y(n_1826) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
OAI31xp33_ASAP7_75t_L g1213 ( .A1(n_1036), .A2(n_1214), .A3(n_1215), .B(n_1224), .Y(n_1213) );
BUFx8_ASAP7_75t_SL g1036 ( .A(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1037), .Y(n_1288) );
OAI31xp33_ASAP7_75t_L g1802 ( .A1(n_1037), .A2(n_1803), .A3(n_1804), .B(n_1827), .Y(n_1802) );
XNOR2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1192), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1046), .B1(n_1137), .B2(n_1191), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
HB1xp67_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
OA22x2_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1093), .B1(n_1094), .B2(n_1136), .Y(n_1047) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1048), .Y(n_1136) );
XNOR2xp5_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1050), .Y(n_1048) );
NAND2xp5_ASAP7_75t_SL g1063 ( .A(n_1064), .B(n_1073), .Y(n_1063) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
AOI31xp33_ASAP7_75t_SL g1081 ( .A1(n_1082), .A2(n_1086), .A3(n_1089), .B(n_1092), .Y(n_1081) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1084), .Y(n_1857) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1095), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1100), .Y(n_1096) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
NAND4xp25_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1124), .C(n_1128), .D(n_1131), .Y(n_1120) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1126), .Y(n_1218) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1137), .Y(n_1191) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
XNOR2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1140), .Y(n_1138) );
AND4x1_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1143), .C(n_1167), .D(n_1187), .Y(n_1140) );
NOR3xp33_ASAP7_75t_SL g1143 ( .A(n_1144), .B(n_1145), .C(n_1165), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1148), .B1(n_1149), .B2(n_1150), .C(n_1153), .Y(n_1146) );
BUFx2_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1152), .Y(n_1159) );
INVx2_ASAP7_75t_SL g1426 ( .A(n_1152), .Y(n_1426) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_1155), .Y(n_1154) );
OAI221xp5_ASAP7_75t_L g1156 ( .A1(n_1157), .A2(n_1158), .B1(n_1159), .B2(n_1160), .C(n_1161), .Y(n_1156) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
OAI221xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1180), .B1(n_1181), .B2(n_1182), .C(n_1183), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
INVx2_ASAP7_75t_L g1406 ( .A(n_1178), .Y(n_1406) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1190), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1194), .B1(n_1283), .B2(n_1380), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
AO22x2_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1236), .B1(n_1237), .B2(n_1282), .Y(n_1194) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1195), .Y(n_1282) );
AND4x1_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1199), .C(n_1213), .D(n_1233), .Y(n_1196) );
OAI21xp33_ASAP7_75t_L g1220 ( .A1(n_1203), .A2(n_1221), .B(n_1222), .Y(n_1220) );
INVx2_ASAP7_75t_SL g1255 ( .A(n_1205), .Y(n_1255) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1209), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g1377 ( .A1(n_1221), .A2(n_1321), .B1(n_1326), .B2(n_1378), .Y(n_1377) );
AND2x4_ASAP7_75t_L g1349 ( .A(n_1223), .B(n_1344), .Y(n_1349) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1226), .Y(n_1372) );
NOR2xp33_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1235), .Y(n_1233) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
AND4x1_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1258), .C(n_1261), .D(n_1263), .Y(n_1238) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
NOR2xp33_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
INVx2_ASAP7_75t_SL g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1271), .Y(n_1811) );
INVx2_ASAP7_75t_SL g1271 ( .A(n_1272), .Y(n_1271) );
OAI22xp5_ASAP7_75t_L g1498 ( .A1(n_1275), .A2(n_1499), .B1(n_1500), .B2(n_1501), .Y(n_1498) );
HB1xp67_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx2_ASAP7_75t_L g1380 ( .A(n_1284), .Y(n_1380) );
XNOR2x1_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1286), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1338), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1287 ( .A1(n_1288), .A2(n_1289), .B1(n_1332), .B2(n_1333), .Y(n_1287) );
NAND3xp33_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1309), .C(n_1325), .Y(n_1289) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_1291), .A2(n_1296), .B1(n_1300), .B2(n_1302), .C(n_1303), .Y(n_1290) );
BUFx2_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
HB1xp67_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
AOI21xp5_ASAP7_75t_L g1421 ( .A1(n_1300), .A2(n_1411), .B(n_1422), .Y(n_1421) );
AOI221xp5_ASAP7_75t_L g1516 ( .A1(n_1300), .A2(n_1506), .B1(n_1517), .B2(n_1521), .C(n_1524), .Y(n_1516) );
INVx2_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1307 ( .A(n_1308), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1309 ( .A1(n_1310), .A2(n_1317), .B1(n_1319), .B2(n_1321), .C(n_1322), .Y(n_1309) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
AOI221xp5_ASAP7_75t_L g1430 ( .A1(n_1319), .A2(n_1322), .B1(n_1417), .B2(n_1431), .C(n_1436), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1526 ( .A1(n_1319), .A2(n_1322), .B1(n_1512), .B2(n_1527), .C(n_1531), .Y(n_1526) );
BUFx6f_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_SL g1323 ( .A(n_1324), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g1325 ( .A1(n_1326), .A2(n_1327), .B1(n_1329), .B2(n_1330), .Y(n_1325) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_1327), .A2(n_1330), .B1(n_1413), .B2(n_1416), .Y(n_1437) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_1327), .A2(n_1330), .B1(n_1509), .B2(n_1511), .Y(n_1532) );
INVx6_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
INVx4_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AOI21xp33_ASAP7_75t_L g1418 ( .A1(n_1333), .A2(n_1419), .B(n_1420), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_1333), .A2(n_1514), .B1(n_1515), .B2(n_1533), .Y(n_1513) );
INVx5_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
AND2x4_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1337), .Y(n_1334) );
INVx3_ASAP7_75t_L g1356 ( .A(n_1336), .Y(n_1356) );
NOR3xp33_ASAP7_75t_SL g1338 ( .A(n_1339), .B(n_1352), .C(n_1362), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1347), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_1341), .A2(n_1342), .B1(n_1345), .B2(n_1346), .Y(n_1340) );
BUFx2_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
BUFx2_ASAP7_75t_L g1390 ( .A(n_1343), .Y(n_1390) );
BUFx2_ASAP7_75t_L g1486 ( .A(n_1343), .Y(n_1486) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_1346), .A2(n_1389), .B1(n_1390), .B2(n_1391), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g1484 ( .A1(n_1346), .A2(n_1485), .B1(n_1486), .B2(n_1487), .Y(n_1484) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1349), .B1(n_1350), .B2(n_1351), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_1349), .A2(n_1393), .B1(n_1394), .B2(n_1395), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_1349), .A2(n_1351), .B1(n_1489), .B2(n_1490), .Y(n_1488) );
INVx2_ASAP7_75t_SL g1353 ( .A(n_1354), .Y(n_1353) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
NAND2x1p5_ASAP7_75t_L g1358 ( .A(n_1356), .B(n_1359), .Y(n_1358) );
BUFx4f_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
BUFx4f_ASAP7_75t_L g1492 ( .A(n_1358), .Y(n_1492) );
BUFx2_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
BUFx2_ASAP7_75t_L g1397 ( .A(n_1361), .Y(n_1397) );
OAI33xp33_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1366), .A3(n_1370), .B1(n_1376), .B2(n_1377), .B3(n_1379), .Y(n_1362) );
OAI33xp33_ASAP7_75t_L g1398 ( .A1(n_1363), .A2(n_1379), .A3(n_1399), .B1(n_1404), .B2(n_1410), .B3(n_1414), .Y(n_1398) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
OAI33xp33_ASAP7_75t_L g1493 ( .A1(n_1365), .A2(n_1379), .A3(n_1494), .B1(n_1498), .B2(n_1504), .B3(n_1510), .Y(n_1493) );
OAI33xp33_ASAP7_75t_L g1880 ( .A1(n_1365), .A2(n_1881), .A3(n_1884), .B1(n_1885), .B2(n_1887), .B3(n_1890), .Y(n_1880) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_1371), .A2(n_1373), .B1(n_1374), .B2(n_1375), .Y(n_1370) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
OAI22xp33_ASAP7_75t_L g1494 ( .A1(n_1378), .A2(n_1495), .B1(n_1496), .B2(n_1497), .Y(n_1494) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1381), .Y(n_1536) );
XNOR2xp5_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1438), .Y(n_1381) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
XNOR2x1_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1385), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1418), .Y(n_1385) );
NOR3xp33_ASAP7_75t_SL g1386 ( .A(n_1387), .B(n_1396), .C(n_1398), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1392), .Y(n_1387) );
OAI211xp5_ASAP7_75t_L g1425 ( .A1(n_1391), .A2(n_1426), .B(n_1427), .C(n_1428), .Y(n_1425) );
INVx3_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_1405), .A2(n_1406), .B1(n_1407), .B2(n_1408), .Y(n_1404) );
OAI22xp5_ASAP7_75t_L g1410 ( .A1(n_1406), .A2(n_1411), .B1(n_1412), .B2(n_1413), .Y(n_1410) );
OAI22xp5_ASAP7_75t_L g1885 ( .A1(n_1408), .A2(n_1814), .B1(n_1860), .B2(n_1886), .Y(n_1885) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_SL g1423 ( .A(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_1439), .A2(n_1479), .B1(n_1534), .B2(n_1535), .Y(n_1438) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1439), .Y(n_1534) );
NAND4xp25_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1463), .C(n_1476), .D(n_1478), .Y(n_1440) );
OAI221xp5_ASAP7_75t_L g1442 ( .A1(n_1443), .A2(n_1446), .B1(n_1449), .B2(n_1452), .C(n_1455), .Y(n_1442) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1470), .Y(n_1867) );
INVx2_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1479), .Y(n_1535) );
HB1xp67_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1481 ( .A(n_1482), .B(n_1513), .Y(n_1481) );
NOR3xp33_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1491), .C(n_1493), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_1484), .B(n_1488), .Y(n_1483) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g1504 ( .A1(n_1505), .A2(n_1506), .B1(n_1507), .B2(n_1509), .Y(n_1504) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
NAND3xp33_ASAP7_75t_L g1515 ( .A(n_1516), .B(n_1526), .C(n_1532), .Y(n_1515) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
OAI221xp5_ASAP7_75t_SL g1537 ( .A1(n_1538), .A2(n_1780), .B1(n_1782), .B2(n_1830), .C(n_1836), .Y(n_1537) );
AND5x1_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1699), .C(n_1746), .D(n_1759), .E(n_1773), .Y(n_1538) );
OAI31xp33_ASAP7_75t_SL g1539 ( .A1(n_1540), .A2(n_1625), .A3(n_1660), .B(n_1689), .Y(n_1539) );
OAI322xp33_ASAP7_75t_L g1540 ( .A1(n_1541), .A2(n_1571), .A3(n_1589), .B1(n_1593), .B2(n_1599), .C1(n_1612), .C2(n_1614), .Y(n_1540) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
A2O1A1Ixp33_ASAP7_75t_L g1720 ( .A1(n_1542), .A2(n_1601), .B(n_1657), .C(n_1721), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1563), .Y(n_1542) );
NOR2xp33_ASAP7_75t_L g1652 ( .A(n_1543), .B(n_1637), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1543), .B(n_1589), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1543), .B(n_1632), .Y(n_1710) );
NAND2xp5_ASAP7_75t_L g1754 ( .A(n_1543), .B(n_1610), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1772 ( .A(n_1543), .B(n_1564), .Y(n_1772) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1543), .Y(n_1778) );
INVx4_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx3_ASAP7_75t_L g1595 ( .A(n_1544), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1544), .B(n_1634), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1544), .B(n_1632), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1544), .B(n_1640), .Y(n_1726) );
NOR3xp33_ASAP7_75t_L g1732 ( .A(n_1544), .B(n_1598), .C(n_1689), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1544), .B(n_1610), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1544), .B(n_1564), .Y(n_1763) );
NOR2xp33_ASAP7_75t_L g1774 ( .A(n_1544), .B(n_1587), .Y(n_1774) );
AND2x4_ASAP7_75t_L g1544 ( .A(n_1545), .B(n_1557), .Y(n_1544) );
AND2x4_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1552), .Y(n_1546) );
OAI21xp33_ASAP7_75t_SL g1895 ( .A1(n_1547), .A2(n_1893), .B(n_1896), .Y(n_1895) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1548), .B(n_1553), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1551), .Y(n_1548) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1551), .Y(n_1560) );
AND2x4_ASAP7_75t_L g1554 ( .A(n_1552), .B(n_1555), .Y(n_1554) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1581 ( .A(n_1553), .B(n_1556), .Y(n_1581) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1558), .Y(n_1692) );
AND2x4_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1561), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1559), .B(n_1561), .Y(n_1569) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
AND2x4_ASAP7_75t_L g1562 ( .A(n_1560), .B(n_1561), .Y(n_1562) );
INVx2_ASAP7_75t_L g1605 ( .A(n_1562), .Y(n_1605) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1563), .Y(n_1658) );
AOI22xp33_ASAP7_75t_L g1713 ( .A1(n_1563), .A2(n_1714), .B1(n_1716), .B2(n_1719), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1563), .B(n_1602), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1567), .Y(n_1563) );
INVx1_ASAP7_75t_SL g1611 ( .A(n_1564), .Y(n_1611) );
CKINVDCx5p33_ASAP7_75t_R g1619 ( .A(n_1564), .Y(n_1619) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1564), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1564), .B(n_1620), .Y(n_1656) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1564), .Y(n_1683) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1564), .Y(n_1757) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1566), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1567), .B(n_1611), .Y(n_1610) );
CKINVDCx6p67_ASAP7_75t_R g1620 ( .A(n_1567), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1567), .B(n_1637), .Y(n_1642) );
CKINVDCx5p33_ASAP7_75t_R g1678 ( .A(n_1567), .Y(n_1678) );
AOI221xp5_ASAP7_75t_L g1746 ( .A1(n_1567), .A2(n_1703), .B1(n_1747), .B2(n_1749), .C(n_1751), .Y(n_1746) );
OR2x6_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1570), .Y(n_1567) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1587), .Y(n_1571) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1573), .B(n_1590), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1659 ( .A(n_1573), .B(n_1589), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_1573), .B(n_1662), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_1573), .B(n_1655), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1582), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1574), .B(n_1583), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1574), .B(n_1589), .Y(n_1649) );
INVx2_ASAP7_75t_L g1739 ( .A(n_1574), .Y(n_1739) );
NAND2xp5_ASAP7_75t_L g1753 ( .A(n_1574), .B(n_1634), .Y(n_1753) );
NOR2xp33_ASAP7_75t_L g1779 ( .A(n_1574), .B(n_1634), .Y(n_1779) );
INVx2_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1575), .B(n_1583), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1575), .B(n_1582), .Y(n_1632) );
OAI22xp5_ASAP7_75t_L g1576 ( .A1(n_1577), .A2(n_1578), .B1(n_1580), .B2(n_1581), .Y(n_1576) );
OAI22xp33_ASAP7_75t_L g1584 ( .A1(n_1578), .A2(n_1581), .B1(n_1585), .B2(n_1586), .Y(n_1584) );
OAI22xp33_ASAP7_75t_L g1606 ( .A1(n_1578), .A2(n_1607), .B1(n_1608), .B2(n_1609), .Y(n_1606) );
BUFx3_ASAP7_75t_L g1695 ( .A(n_1578), .Y(n_1695) );
BUFx6f_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
HB1xp67_ASAP7_75t_L g1609 ( .A(n_1581), .Y(n_1609) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1581), .Y(n_1698) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1583), .Y(n_1598) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1588), .B(n_1590), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1588), .B(n_1633), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1588), .B(n_1589), .Y(n_1704) );
NOR2x1_ASAP7_75t_L g1597 ( .A(n_1589), .B(n_1598), .Y(n_1597) );
OR2x2_ASAP7_75t_L g1638 ( .A(n_1589), .B(n_1639), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1589), .B(n_1668), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1589), .B(n_1598), .Y(n_1722) );
INVx2_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
BUFx3_ASAP7_75t_L g1634 ( .A(n_1590), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1680 ( .A(n_1590), .B(n_1681), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1590), .B(n_1598), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1768 ( .A(n_1590), .B(n_1632), .Y(n_1768) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
NOR2xp33_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1596), .Y(n_1594) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1595), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1595), .B(n_1640), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1595), .B(n_1649), .Y(n_1648) );
NAND2xp5_ASAP7_75t_L g1674 ( .A(n_1595), .B(n_1613), .Y(n_1674) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1595), .B(n_1677), .Y(n_1676) );
OAI21xp5_ASAP7_75t_SL g1712 ( .A1(n_1595), .A2(n_1713), .B(n_1720), .Y(n_1712) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
OAI21xp33_ASAP7_75t_L g1650 ( .A1(n_1598), .A2(n_1651), .B(n_1653), .Y(n_1650) );
OR2x2_ASAP7_75t_L g1729 ( .A(n_1598), .B(n_1634), .Y(n_1729) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1601), .B(n_1610), .Y(n_1600) );
INVx2_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
INVx2_ASAP7_75t_L g1624 ( .A(n_1602), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1745 ( .A(n_1602), .B(n_1690), .Y(n_1745) );
INVx2_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx2_ASAP7_75t_SL g1637 ( .A(n_1603), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1603), .B(n_1620), .Y(n_1646) );
OR2x2_ASAP7_75t_L g1688 ( .A(n_1603), .B(n_1623), .Y(n_1688) );
INVx2_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
NAND2xp5_ASAP7_75t_L g1645 ( .A(n_1611), .B(n_1646), .Y(n_1645) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1612), .B(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
NOR2xp33_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1621), .Y(n_1614) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
NAND2xp5_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1618), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1617), .B(n_1704), .Y(n_1703) );
OR2x2_ASAP7_75t_L g1728 ( .A(n_1617), .B(n_1729), .Y(n_1728) );
A2O1A1Ixp33_ASAP7_75t_L g1760 ( .A1(n_1617), .A2(n_1715), .B(n_1736), .C(n_1761), .Y(n_1760) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1618), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1620), .Y(n_1618) );
INVx3_ASAP7_75t_L g1623 ( .A(n_1619), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_1619), .B(n_1636), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1619), .B(n_1703), .Y(n_1702) );
NOR2xp33_ASAP7_75t_L g1706 ( .A(n_1619), .B(n_1707), .Y(n_1706) );
OAI32xp33_ASAP7_75t_L g1755 ( .A1(n_1619), .A2(n_1687), .A3(n_1704), .B1(n_1710), .B2(n_1756), .Y(n_1755) );
AND2x4_ASAP7_75t_SL g1636 ( .A(n_1620), .B(n_1637), .Y(n_1636) );
OR2x2_ASAP7_75t_L g1672 ( .A(n_1620), .B(n_1637), .Y(n_1672) );
NOR2xp33_ASAP7_75t_L g1716 ( .A(n_1620), .B(n_1717), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1737 ( .A(n_1620), .B(n_1718), .Y(n_1737) );
NAND3xp33_ASAP7_75t_L g1761 ( .A(n_1620), .B(n_1721), .C(n_1762), .Y(n_1761) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
OAI322xp33_ASAP7_75t_L g1766 ( .A1(n_1622), .A2(n_1635), .A3(n_1685), .B1(n_1688), .B2(n_1717), .C1(n_1767), .C2(n_1769), .Y(n_1766) );
NAND2xp5_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1624), .Y(n_1622) );
NOR2xp33_ASAP7_75t_L g1665 ( .A(n_1623), .B(n_1666), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1748 ( .A(n_1623), .B(n_1637), .Y(n_1748) );
OR2x2_ASAP7_75t_L g1750 ( .A(n_1623), .B(n_1631), .Y(n_1750) );
AOI21xp5_ASAP7_75t_L g1776 ( .A1(n_1623), .A2(n_1770), .B(n_1777), .Y(n_1776) );
NAND2xp5_ASAP7_75t_L g1758 ( .A(n_1624), .B(n_1690), .Y(n_1758) );
OAI221xp5_ASAP7_75t_SL g1625 ( .A1(n_1626), .A2(n_1635), .B1(n_1638), .B2(n_1641), .C(n_1643), .Y(n_1625) );
INVxp67_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1630), .Y(n_1627) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1631 ( .A(n_1632), .B(n_1633), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1632), .B(n_1655), .Y(n_1654) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1632), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1633), .B(n_1640), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1634), .B(n_1710), .Y(n_1709) );
OR2x2_ASAP7_75t_L g1730 ( .A(n_1634), .B(n_1726), .Y(n_1730) );
NOR2xp33_ASAP7_75t_L g1727 ( .A(n_1635), .B(n_1728), .Y(n_1727) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx2_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1642), .B(n_1683), .Y(n_1682) );
AOI21xp5_ASAP7_75t_L g1724 ( .A1(n_1642), .A2(n_1725), .B(n_1727), .Y(n_1724) );
AOI221xp5_ASAP7_75t_L g1643 ( .A1(n_1644), .A2(n_1647), .B1(n_1650), .B2(n_1656), .C(n_1657), .Y(n_1643) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1646), .Y(n_1711) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1656), .Y(n_1765) );
NOR2xp33_ASAP7_75t_L g1657 ( .A(n_1658), .B(n_1659), .Y(n_1657) );
NOR2xp33_ASAP7_75t_L g1764 ( .A(n_1659), .B(n_1765), .Y(n_1764) );
NAND4xp25_ASAP7_75t_L g1660 ( .A(n_1661), .B(n_1664), .C(n_1670), .D(n_1675), .Y(n_1660) );
O2A1O1Ixp33_ASAP7_75t_L g1773 ( .A1(n_1662), .A2(n_1667), .B(n_1774), .C(n_1775), .Y(n_1773) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1665), .Y(n_1664) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1673), .Y(n_1670) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
AOI221xp5_ASAP7_75t_L g1675 ( .A1(n_1676), .A2(n_1678), .B1(n_1679), .B2(n_1682), .C(n_1684), .Y(n_1675) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1677), .Y(n_1707) );
INVx1_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
AOI21xp33_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1686), .B(n_1688), .Y(n_1684) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
OAI221xp5_ASAP7_75t_SL g1723 ( .A1(n_1688), .A2(n_1717), .B1(n_1724), .B2(n_1730), .C(n_1731), .Y(n_1723) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
BUFx3_ASAP7_75t_L g1718 ( .A(n_1690), .Y(n_1718) );
O2A1O1Ixp33_ASAP7_75t_L g1759 ( .A1(n_1690), .A2(n_1760), .B(n_1764), .C(n_1766), .Y(n_1759) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
OAI22xp33_ASAP7_75t_L g1693 ( .A1(n_1694), .A2(n_1695), .B1(n_1696), .B2(n_1697), .Y(n_1693) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1695), .Y(n_1781) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
NOR5xp2_ASAP7_75t_L g1699 ( .A(n_1700), .B(n_1712), .C(n_1723), .D(n_1734), .E(n_1738), .Y(n_1699) );
AOI31xp33_ASAP7_75t_L g1700 ( .A1(n_1701), .A2(n_1705), .A3(n_1708), .B(n_1711), .Y(n_1700) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1704), .Y(n_1715) );
OAI21xp33_ASAP7_75t_L g1731 ( .A1(n_1704), .A2(n_1732), .B(n_1733), .Y(n_1731) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
AOI31xp33_ASAP7_75t_L g1734 ( .A1(n_1708), .A2(n_1735), .A3(n_1736), .B(n_1737), .Y(n_1734) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
INVx2_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1726), .Y(n_1725) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1733), .Y(n_1735) );
O2A1O1Ixp33_ASAP7_75t_L g1738 ( .A1(n_1739), .A2(n_1740), .B(n_1742), .C(n_1744), .Y(n_1738) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
OAI22xp5_ASAP7_75t_L g1775 ( .A1(n_1742), .A2(n_1744), .B1(n_1765), .B2(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
O2A1O1Ixp33_ASAP7_75t_SL g1751 ( .A1(n_1752), .A2(n_1754), .B(n_1755), .C(n_1758), .Y(n_1751) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
NOR2xp33_ASAP7_75t_L g1770 ( .A(n_1753), .B(n_1771), .Y(n_1770) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1768), .Y(n_1767) );
INVxp67_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1778), .B(n_1779), .Y(n_1777) );
INVx1_ASAP7_75t_L g1780 ( .A(n_1781), .Y(n_1780) );
BUFx2_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
BUFx2_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
NAND4xp75_ASAP7_75t_L g1785 ( .A(n_1786), .B(n_1802), .C(n_1828), .D(n_1829), .Y(n_1785) );
AND2x2_ASAP7_75t_SL g1786 ( .A(n_1787), .B(n_1798), .Y(n_1786) );
AOI33xp33_ASAP7_75t_L g1787 ( .A1(n_1788), .A2(n_1789), .A3(n_1792), .B1(n_1794), .B2(n_1795), .B3(n_1797), .Y(n_1787) );
BUFx2_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
OAI221xp5_ASAP7_75t_L g1804 ( .A1(n_1805), .A2(n_1809), .B1(n_1813), .B2(n_1819), .C(n_1822), .Y(n_1804) );
OAI22xp5_ASAP7_75t_L g1813 ( .A1(n_1814), .A2(n_1815), .B1(n_1816), .B2(n_1818), .Y(n_1813) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
AOI21xp5_ASAP7_75t_L g1822 ( .A1(n_1823), .A2(n_1824), .B(n_1825), .Y(n_1822) );
CKINVDCx14_ASAP7_75t_R g1830 ( .A(n_1831), .Y(n_1830) );
INVx4_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1833), .Y(n_1832) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVxp33_ASAP7_75t_SL g1837 ( .A(n_1838), .Y(n_1837) );
HB1xp67_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
NOR2xp33_ASAP7_75t_L g1862 ( .A(n_1863), .B(n_1880), .Y(n_1862) );
OAI22xp5_ASAP7_75t_L g1864 ( .A1(n_1865), .A2(n_1866), .B1(n_1868), .B2(n_1869), .Y(n_1864) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1883), .Y(n_1882) );
BUFx2_ASAP7_75t_L g1891 ( .A(n_1892), .Y(n_1891) );
HB1xp67_ASAP7_75t_L g1894 ( .A(n_1895), .Y(n_1894) );
endmodule