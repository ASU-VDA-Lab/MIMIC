module fake_jpeg_5861_n_165 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g21 ( 
.A(n_0),
.B(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_31),
.B(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_34),
.B(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_29),
.B1(n_20),
.B2(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_3),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_18),
.B(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_29),
.B1(n_20),
.B2(n_17),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_54),
.B1(n_27),
.B2(n_22),
.Y(n_81)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_51),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_62),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_56),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_55),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_34),
.B1(n_33),
.B2(n_38),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_23),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_19),
.B1(n_30),
.B2(n_16),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_63),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_14),
.B1(n_25),
.B2(n_24),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_30),
.B1(n_19),
.B2(n_11),
.Y(n_90)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_78),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_19),
.B(n_30),
.C(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_91),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_94),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_19),
.B1(n_30),
.B2(n_10),
.Y(n_89)
);

NOR4xp25_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_7),
.C(n_8),
.D(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_6),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_6),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_57),
.B(n_58),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_46),
.B(n_50),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_105),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_62),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_95),
.A3(n_88),
.B1(n_77),
.B2(n_78),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_87),
.B1(n_93),
.B2(n_13),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_91),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_49),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_47),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_92),
.B(n_86),
.C(n_95),
.D(n_90),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_107),
.B(n_113),
.C(n_102),
.D(n_101),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_108),
.B(n_110),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_121),
.B(n_112),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_78),
.B1(n_47),
.B2(n_80),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_128),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_76),
.B(n_73),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_72),
.C(n_80),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_97),
.C(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_136),
.C(n_137),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_128),
.B1(n_115),
.B2(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_139),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_114),
.A3(n_125),
.B1(n_117),
.B2(n_126),
.C1(n_105),
.C2(n_96),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_135),
.CI(n_121),
.CON(n_141),
.SN(n_141)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_106),
.C(n_101),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_106),
.C(n_70),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_70),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_145),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_125),
.B1(n_133),
.B2(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_120),
.C(n_118),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_147),
.C(n_48),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_119),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_124),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_148),
.B(n_131),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_151),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_135),
.C(n_9),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_142),
.C(n_144),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_9),
.B(n_13),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_7),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_154),
.B(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_158),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_153),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_143),
.C(n_93),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_159),
.Y(n_165)
);


endmodule