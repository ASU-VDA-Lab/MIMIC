module fake_jpeg_27786_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_18),
.Y(n_56)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_55),
.B1(n_35),
.B2(n_37),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_74),
.B1(n_82),
.B2(n_16),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_16),
.B(n_30),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_67),
.C(n_89),
.Y(n_115)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_76),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_70),
.B(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_32),
.B1(n_39),
.B2(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_41),
.CI(n_39),
.CON(n_80),
.SN(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_83),
.Y(n_104)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_39),
.B1(n_22),
.B2(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_16),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_17),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_46),
.B(n_21),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_19),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

AO22x2_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_34),
.B1(n_36),
.B2(n_33),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_94),
.B1(n_97),
.B2(n_103),
.Y(n_126)
);

NAND2x1p5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_34),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_34),
.Y(n_138)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_118),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_81),
.B1(n_72),
.B2(n_62),
.Y(n_137)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_14),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_112),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_117),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_121),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_79),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_75),
.B(n_79),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_138),
.B(n_118),
.Y(n_155)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_140),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_124),
.B(n_129),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_125),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_133),
.B1(n_95),
.B2(n_98),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_136),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_101),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_17),
.B1(n_23),
.B2(n_27),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_137),
.B1(n_23),
.B2(n_24),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_77),
.B1(n_73),
.B2(n_61),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_88),
.B1(n_85),
.B2(n_63),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_29),
.B1(n_27),
.B2(n_23),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_63),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_72),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_68),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_62),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_22),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_105),
.B(n_30),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_26),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_147),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_129),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_175),
.B(n_135),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_164),
.C(n_168),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_109),
.B1(n_108),
.B2(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_156),
.B1(n_162),
.B2(n_167),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_122),
.B(n_127),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_102),
.B1(n_92),
.B2(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_114),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_26),
.C(n_29),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_25),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_169),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_134),
.B1(n_120),
.B2(n_138),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_121),
.C(n_138),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_179),
.C(n_197),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_138),
.C(n_120),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_0),
.B(n_2),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_192),
.B(n_194),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g210 ( 
.A(n_187),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_124),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_140),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_193),
.B1(n_173),
.B2(n_166),
.Y(n_200)
);

NOR4xp25_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_143),
.C(n_142),
.D(n_145),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_195),
.B1(n_24),
.B2(n_2),
.C(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_130),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_170),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_160),
.B(n_148),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_135),
.C(n_123),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_155),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_209),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_172),
.B1(n_165),
.B2(n_151),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_206),
.B1(n_208),
.B2(n_213),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_152),
.C(n_168),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_178),
.C(n_197),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_154),
.B1(n_156),
.B2(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_167),
.B1(n_159),
.B2(n_161),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_161),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_162),
.B1(n_24),
.B2(n_0),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_194),
.B1(n_192),
.B2(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_0),
.B(n_183),
.Y(n_226)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_193),
.B(n_180),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_195),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_226),
.B1(n_213),
.B2(n_208),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_231),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_185),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_232),
.B(n_201),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_220),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_201),
.C(n_209),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_238),
.C(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_205),
.C(n_203),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_239),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_180),
.C(n_187),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_211),
.B1(n_217),
.B2(n_199),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_225),
.B1(n_216),
.B2(n_221),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_187),
.C(n_199),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_221),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_188),
.B(n_215),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_244),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_250),
.B(n_184),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_227),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_252),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_251),
.Y(n_255)
);

OAI221xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_224),
.B1(n_226),
.B2(n_219),
.C(n_187),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_184),
.B1(n_6),
.B2(n_7),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_255),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_244),
.B(n_240),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_259),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_258),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_238),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_249),
.C(n_251),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_265),
.C(n_5),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_249),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_5),
.C(n_8),
.Y(n_267)
);

A2O1A1O1Ixp25_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_8),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_263),
.B(n_261),
.Y(n_269)
);

OAI321xp33_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_271)
);

AOI31xp33_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_270),
.A3(n_13),
.B(n_15),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_12),
.Y(n_273)
);


endmodule