module real_jpeg_30210_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_313, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_313;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_0),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_0),
.A2(n_58),
.B1(n_62),
.B2(n_64),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_1),
.B(n_62),
.Y(n_91)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_1),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_2),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_133),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_62),
.B1(n_64),
.B2(n_133),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_133),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_3),
.A2(n_40),
.B1(n_55),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_3),
.A2(n_40),
.B1(n_62),
.B2(n_64),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_6),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_6),
.A2(n_33),
.B(n_37),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_161),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_35),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_6),
.A2(n_55),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_6),
.B(n_55),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_6),
.B(n_59),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_6),
.A2(n_90),
.B1(n_250),
.B2(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_6),
.A2(n_36),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_7),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_150),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_150),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_7),
.A2(n_62),
.B1(n_64),
.B2(n_150),
.Y(n_244)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_9),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_46),
.B1(n_62),
.B2(n_64),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_10),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_100),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_100),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_10),
.A2(n_62),
.B1(n_64),
.B2(n_100),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_30),
.B1(n_55),
.B2(n_56),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_11),
.A2(n_30),
.B1(n_62),
.B2(n_64),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_12),
.A2(n_55),
.A3(n_64),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_13),
.A2(n_62),
.B1(n_64),
.B2(n_69),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_69),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_16),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_17),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_17),
.A2(n_36),
.B1(n_37),
.B2(n_157),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_17),
.A2(n_55),
.B1(n_56),
.B2(n_157),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_17),
.A2(n_62),
.B1(n_64),
.B2(n_157),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_101),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_22),
.B(n_101),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_73),
.C(n_79),
.Y(n_22)
);

FAx1_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_73),
.CI(n_79),
.CON(n_134),
.SN(n_134)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_72),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_24),
.A2(n_25),
.B1(n_103),
.B2(n_111),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_43),
.C(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_39),
.B2(n_41),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_26),
.A2(n_31),
.B1(n_41),
.B2(n_98),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_33),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_28),
.A2(n_38),
.B(n_161),
.C(n_162),
.Y(n_160)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_31),
.A2(n_41),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_32),
.A2(n_35),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_32),
.A2(n_35),
.B1(n_99),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_32),
.A2(n_35),
.B1(n_132),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_32),
.A2(n_35),
.B1(n_156),
.B2(n_194),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_49),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_36),
.A2(n_53),
.A3(n_56),
.B1(n_267),
.B2(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_37),
.B(n_161),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_60),
.B1(n_70),
.B2(n_71),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_57),
.B2(n_59),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_48),
.B1(n_52),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_47),
.A2(n_57),
.B1(n_59),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_47),
.A2(n_59),
.B1(n_76),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_47),
.A2(n_59),
.B1(n_125),
.B2(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_47),
.A2(n_59),
.B1(n_188),
.B2(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_48),
.A2(n_52),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_48),
.A2(n_52),
.B1(n_167),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_48),
.A2(n_52),
.B1(n_200),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_53),
.Y(n_276)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_55),
.B(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_71),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_68),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_66),
.B1(n_68),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_61),
.A2(n_66),
.B1(n_85),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_61),
.A2(n_66),
.B1(n_130),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_61),
.A2(n_66),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_61),
.A2(n_66),
.B1(n_225),
.B2(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_61),
.B(n_161),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_61),
.A2(n_66),
.B1(n_192),
.B2(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_62),
.B(n_65),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_62),
.B(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_96),
.B(n_97),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_81),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_82),
.A2(n_83),
.B1(n_89),
.B2(n_96),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_86),
.A2(n_88),
.B1(n_146),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_86),
.A2(n_88),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_96),
.B1(n_97),
.B2(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B(n_95),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_92),
.B1(n_95),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_94),
.B1(n_128),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_90),
.A2(n_94),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_90),
.A2(n_94),
.B1(n_244),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_90),
.A2(n_239),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_91),
.A2(n_143),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_91),
.A2(n_93),
.B1(n_164),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_91),
.A2(n_93),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g278 ( 
.A(n_93),
.Y(n_278)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_94),
.B(n_161),
.Y(n_256)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_135),
.B(n_309),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_134),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_116),
.B(n_134),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_121),
.Y(n_179)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_122),
.A2(n_123),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.C(n_131),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_124),
.B(n_126),
.CI(n_131),
.CON(n_173),
.SN(n_173)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_129),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_134),
.Y(n_310)
);

AOI321xp33_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_175),
.A3(n_180),
.B1(n_303),
.B2(n_308),
.C(n_313),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_137),
.A2(n_304),
.B(n_307),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_170),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_138),
.B(n_170),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_153),
.C(n_169),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_139),
.B(n_169),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_148),
.C(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_144),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.C(n_166),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_154),
.B(n_166),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_159),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_163),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.C(n_174),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_173),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_176),
.B(n_177),
.Y(n_308)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_210),
.C(n_215),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_204),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_182),
.B(n_204),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_195),
.C(n_196),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_183),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_193),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_190),
.C(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_195),
.Y(n_301)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_198),
.B(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_201),
.B(n_203),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_202),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.C(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_211),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_212),
.B(n_213),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_297),
.B(n_302),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_283),
.B(n_296),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_260),
.B(n_282),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_240),
.B(n_259),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_230),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_235),
.C(n_237),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_236),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_238),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_258),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_246),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_252),
.B(n_257),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_262),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_273),
.B1(n_280),
.B2(n_281),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_272),
.C(n_281),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_270),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_273),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_277),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_292),
.C(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);


endmodule