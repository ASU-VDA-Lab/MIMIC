module real_jpeg_8639_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_1),
.B(n_25),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_1),
.B(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_3),
.B(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR4xp25_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_26),
.C(n_29),
.D(n_33),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_10),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_15),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_14),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_21),
.Y(n_18)
);


endmodule