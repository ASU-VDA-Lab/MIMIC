module fake_jpeg_2541_n_86 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_28),
.Y(n_47)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.C(n_47),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_26),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_31),
.C(n_25),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_24),
.C(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_16),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_33),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_58),
.B1(n_56),
.B2(n_44),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_24),
.B(n_5),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_63),
.C(n_4),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_76),
.B1(n_77),
.B2(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_68),
.B(n_9),
.C(n_10),
.Y(n_85)
);

OAI322xp33_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_7),
.A3(n_13),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_22),
.Y(n_86)
);


endmodule