module fake_jpeg_1922_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_46),
.B(n_50),
.Y(n_117)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_52),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_7),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_9),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_16),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_62),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_18),
.B(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_69),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_6),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_82),
.Y(n_126)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_22),
.B(n_30),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_87),
.Y(n_135)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_89),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_31),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_24),
.B1(n_41),
.B2(n_34),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_95),
.A2(n_124),
.B1(n_136),
.B2(n_102),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_96),
.A2(n_97),
.B1(n_108),
.B2(n_114),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_42),
.B1(n_32),
.B2(n_37),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_82),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_48),
.A2(n_32),
.B1(n_39),
.B2(n_37),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_39),
.B1(n_31),
.B2(n_29),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_61),
.A2(n_31),
.B1(n_29),
.B2(n_0),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_125),
.B1(n_128),
.B2(n_133),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_73),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_51),
.A2(n_31),
.B1(n_0),
.B2(n_4),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_51),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_53),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_68),
.A2(n_12),
.B1(n_14),
.B2(n_76),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_53),
.A2(n_65),
.B1(n_85),
.B2(n_81),
.Y(n_137)
);

OAI22x1_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_131),
.B1(n_121),
.B2(n_116),
.Y(n_156)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_74),
.B1(n_72),
.B2(n_92),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_156),
.B1(n_113),
.B2(n_141),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_144),
.B(n_158),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_101),
.A2(n_80),
.A3(n_79),
.B1(n_83),
.B2(n_89),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_151),
.Y(n_180)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_153),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_161),
.Y(n_194)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_132),
.B1(n_111),
.B2(n_99),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_157),
.A2(n_160),
.B1(n_167),
.B2(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_159),
.B(n_165),
.Y(n_198)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_164),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_105),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_100),
.B(n_134),
.Y(n_166)
);

OAI221xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_174),
.C(n_176),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_123),
.B1(n_130),
.B2(n_107),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_94),
.B(n_103),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_106),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_127),
.A2(n_106),
.B1(n_137),
.B2(n_123),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_97),
.B(n_107),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_125),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_133),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_172),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_196),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_128),
.B1(n_141),
.B2(n_130),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_186),
.B1(n_145),
.B2(n_173),
.Y(n_220)
);

OR2x4_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_159),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_198),
.B(n_193),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_178),
.B1(n_144),
.B2(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_150),
.C(n_158),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_202),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_177),
.B1(n_143),
.B2(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_154),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_209),
.Y(n_237)
);

AO22x1_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_149),
.B1(n_161),
.B2(n_170),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_202),
.B(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_215),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_218),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_179),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_223),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_222),
.B1(n_183),
.B2(n_205),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_176),
.B1(n_147),
.B2(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_142),
.B(n_180),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_227),
.B(n_194),
.Y(n_232)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_226),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_200),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_182),
.B1(n_196),
.B2(n_204),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_231),
.B1(n_233),
.B2(n_222),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_202),
.C(n_184),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_225),
.C(n_220),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_181),
.B(n_191),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_185),
.B(n_195),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_195),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_244),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_253),
.B(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_225),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_207),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_262),
.C(n_232),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_258),
.A2(n_231),
.B1(n_233),
.B2(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_246),
.B1(n_255),
.B2(n_223),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_213),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_261),
.B(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_207),
.C(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_268),
.B1(n_271),
.B2(n_273),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_233),
.B1(n_241),
.B2(n_246),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_274),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_241),
.B1(n_245),
.B2(n_240),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_240),
.B1(n_236),
.B2(n_243),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_249),
.A2(n_236),
.B1(n_243),
.B2(n_229),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_254),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_256),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_251),
.Y(n_291)
);

BUFx12_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_280),
.A2(n_281),
.B1(n_284),
.B2(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

OAI22x1_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_254),
.B1(n_251),
.B2(n_236),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_268),
.B1(n_265),
.B2(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_254),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_263),
.C(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_287),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_266),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_263),
.C(n_272),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_290),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_291),
.B(n_283),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_285),
.B(n_276),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_282),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_296),
.B(n_297),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_292),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_300),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_299),
.A2(n_280),
.B1(n_216),
.B2(n_218),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_288),
.C(n_286),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_280),
.B(n_226),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_210),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_306),
.Y(n_307)
);

OAI21x1_ASAP7_75t_SL g308 ( 
.A1(n_307),
.A2(n_305),
.B(n_208),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_214),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_179),
.Y(n_310)
);


endmodule