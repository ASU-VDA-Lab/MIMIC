module fake_jpeg_16954_n_100 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_35),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_2),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_3),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_38),
.B1(n_39),
.B2(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_43),
.B1(n_36),
.B2(n_44),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_40),
.B1(n_37),
.B2(n_4),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_5),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_3),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_40),
.B1(n_19),
.B2(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_72),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_74),
.Y(n_78)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_71),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_4),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_6),
.C(n_7),
.Y(n_80)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_22),
.C(n_8),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_65),
.B1(n_77),
.B2(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_73),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_90),
.C(n_78),
.Y(n_92)
);

OAI322xp33_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_93),
.A3(n_91),
.B1(n_85),
.B2(n_87),
.C1(n_88),
.C2(n_79),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_84),
.C(n_83),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_31),
.B1(n_16),
.B2(n_17),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_15),
.B(n_18),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_23),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_24),
.C(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_29),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_30),
.Y(n_100)
);


endmodule