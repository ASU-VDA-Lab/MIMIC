module fake_jpeg_8498_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_23),
.Y(n_46)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_50),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_28),
.B1(n_32),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_57),
.B1(n_62),
.B2(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_27),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_55),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_19),
.B1(n_63),
.B2(n_18),
.Y(n_101)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_56),
.B(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_28),
.B1(n_32),
.B2(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_67),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_19),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_26),
.B(n_22),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_32),
.B1(n_26),
.B2(n_24),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_30),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_69),
.B(n_83),
.Y(n_133)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_80),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_101),
.B1(n_53),
.B2(n_54),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_37),
.B1(n_19),
.B2(n_41),
.Y(n_74)
);

AOI221xp5_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_76),
.B1(n_104),
.B2(n_89),
.C(n_98),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_36),
.B(n_18),
.C(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_86),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_34),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_33),
.Y(n_88)
);

AOI22x1_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_105),
.B1(n_53),
.B2(n_36),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_92),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_33),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_103),
.Y(n_129)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_18),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_29),
.B(n_24),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_35),
.B(n_31),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_35),
.C(n_31),
.Y(n_125)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_109),
.A2(n_117),
.B1(n_132),
.B2(n_72),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_124),
.B(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_81),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_81),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_100),
.B1(n_78),
.B2(n_97),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_35),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_130),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_90),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_0),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_131),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_35),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g132 ( 
.A1(n_76),
.A2(n_101),
.B1(n_73),
.B2(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_134),
.B(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_162),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_114),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_129),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_158),
.B(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_140),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_84),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_145),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_71),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_92),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_150),
.C(n_113),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_92),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_80),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_153),
.Y(n_166)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_125),
.B1(n_117),
.B2(n_109),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_29),
.B(n_22),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_79),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_121),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_113),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_106),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_182),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_149),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_185),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_153),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_117),
.B1(n_150),
.B2(n_138),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_127),
.B(n_117),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_156),
.B1(n_161),
.B2(n_146),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_199),
.B1(n_208),
.B2(n_209),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_203),
.B1(n_204),
.B2(n_174),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_139),
.Y(n_196)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_128),
.C(n_106),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_202),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_177),
.A2(n_158),
.B(n_154),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_170),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_177),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_168),
.C(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_167),
.C(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_217),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_173),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_206),
.B1(n_163),
.B2(n_195),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_187),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_220),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_172),
.C(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_169),
.B1(n_186),
.B2(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_224),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_164),
.C(n_184),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_226),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_164),
.C(n_171),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_193),
.B(n_205),
.C(n_217),
.D(n_221),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_229),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g229 ( 
.A(n_216),
.B(n_204),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_169),
.B(n_194),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_16),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_0),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_215),
.A2(n_207),
.B(n_178),
.C(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_201),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_112),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_144),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_250),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_225),
.B1(n_220),
.B2(n_213),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_252),
.B1(n_1),
.B2(n_4),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_249),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_251),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_144),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_228),
.B1(n_238),
.B2(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_257),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_237),
.B(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_255),
.C(n_249),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_239),
.B(n_232),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g260 ( 
.A1(n_242),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_7),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g268 ( 
.A(n_261),
.B(n_258),
.CI(n_9),
.CON(n_268),
.SN(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_10),
.Y(n_270)
);

AOI31xp67_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_246),
.A3(n_8),
.B(n_9),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_265),
.B(n_258),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_259),
.B(n_246),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_7),
.C(n_8),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_7),
.C(n_9),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_262),
.C1(n_268),
.C2(n_269),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_11),
.B(n_12),
.Y(n_275)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.C(n_273),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_12),
.B1(n_13),
.B2(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);


endmodule