module fake_jpeg_24546_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_40),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_28),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_45),
.B(n_21),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_18),
.B1(n_23),
.B2(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_30),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_88),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_29),
.B(n_9),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_95),
.B1(n_96),
.B2(n_39),
.Y(n_116)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_40),
.B1(n_57),
.B2(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_108),
.B1(n_74),
.B2(n_34),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_29),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_116),
.B(n_118),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_33),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_40),
.B1(n_36),
.B2(n_51),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_71),
.B1(n_81),
.B2(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_51),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_42),
.B1(n_62),
.B2(n_59),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_61),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_114),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_22),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_39),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_117),
.C(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_41),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_66),
.C(n_55),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_47),
.B1(n_17),
.B2(n_19),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_0),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_0),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_28),
.CI(n_25),
.CON(n_126),
.SN(n_126)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_17),
.B1(n_19),
.B2(n_16),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_17),
.B1(n_32),
.B2(n_22),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_131),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_126),
.A2(n_139),
.B(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_128),
.B(n_130),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_84),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_107),
.B1(n_119),
.B2(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_37),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_70),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_32),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_56),
.B1(n_90),
.B2(n_86),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_148),
.B1(n_119),
.B2(n_120),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_27),
.B(n_33),
.C(n_16),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_32),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_28),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_117),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_115),
.B(n_98),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_24),
.A3(n_26),
.B1(n_30),
.B2(n_25),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_108),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_116),
.B1(n_122),
.B2(n_107),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_157),
.B1(n_164),
.B2(n_170),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_168),
.B1(n_174),
.B2(n_144),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_120),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_165),
.B(n_172),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_118),
.B1(n_123),
.B2(n_113),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_113),
.B(n_115),
.C(n_98),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_101),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_120),
.B1(n_107),
.B2(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_149),
.B1(n_131),
.B2(n_139),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_138),
.C(n_137),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_25),
.C(n_30),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_134),
.B(n_126),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_180),
.B(n_200),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_134),
.B(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_182),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_126),
.B1(n_150),
.B2(n_133),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_189),
.B1(n_191),
.B2(n_156),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_128),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_192),
.C(n_199),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_143),
.B1(n_141),
.B2(n_133),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_202),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_132),
.B1(n_143),
.B2(n_111),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_170),
.B(n_111),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_119),
.B1(n_140),
.B2(n_121),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_101),
.B1(n_27),
.B2(n_33),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_153),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_163),
.B1(n_155),
.B2(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_163),
.B(n_169),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_154),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_203),
.B(n_24),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_27),
.B1(n_16),
.B2(n_92),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_214),
.Y(n_242)
);

XOR2x2_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_172),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_163),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_216),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_156),
.B1(n_166),
.B2(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_161),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_222),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_183),
.A2(n_167),
.B1(n_166),
.B2(n_160),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_218),
.B1(n_198),
.B2(n_187),
.Y(n_244)
);

AO22x1_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_176),
.B1(n_30),
.B2(n_26),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_223),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_26),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_0),
.B(n_1),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_225),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_24),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_8),
.B(n_13),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_199),
.C(n_192),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_241),
.C(n_227),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_245),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_188),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_238),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_194),
.B(n_202),
.C(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_244),
.B1(n_218),
.B2(n_220),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_180),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_215),
.C(n_219),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_181),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_223),
.Y(n_270)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_208),
.B(n_8),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_250),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_208),
.B(n_13),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_15),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_233),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_230),
.C(n_243),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_251),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_207),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_264),
.Y(n_274)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_263),
.B(n_265),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_237),
.B(n_213),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_239),
.B1(n_246),
.B2(n_233),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_212),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_212),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_271),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_252),
.C(n_258),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_216),
.B1(n_242),
.B2(n_240),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_270),
.B1(n_260),
.B2(n_222),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_235),
.B1(n_204),
.B2(n_221),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_297)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_258),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_236),
.B1(n_225),
.B2(n_239),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_229),
.B1(n_271),
.B2(n_228),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_288),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_204),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_1),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_221),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_295),
.C(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_297),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_274),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_0),
.B(n_1),
.Y(n_295)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_275),
.B1(n_6),
.B2(n_7),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_9),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_10),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_12),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_303),
.C(n_286),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_285),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_5),
.C(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_307),
.B(n_313),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_280),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_310),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_275),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_10),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_299),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_292),
.B(n_293),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_302),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_305),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_320),
.B(n_324),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_289),
.B(n_292),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_323),
.A2(n_295),
.B(n_312),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_328),
.B(n_11),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_298),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_327),
.B1(n_330),
.B2(n_5),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_291),
.Y(n_327)
);

AOI21x1_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_290),
.B(n_10),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_11),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_333),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_317),
.C(n_15),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_331),
.B(n_334),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_326),
.B(n_5),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_6),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_6),
.Y(n_341)
);


endmodule