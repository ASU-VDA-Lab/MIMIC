module real_jpeg_24755_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_128;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_48),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_1),
.A2(n_48),
.B1(n_67),
.B2(n_68),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_1),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_66),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_6),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_8),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_8),
.B(n_67),
.C(n_84),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_61),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_8),
.A2(n_69),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_8),
.B(n_98),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_12),
.A2(n_44),
.B1(n_53),
.B2(n_54),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_12),
.A2(n_44),
.B1(n_67),
.B2(n_68),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_13),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_92),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_14),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_206)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_19),
.B(n_112),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_79),
.C(n_100),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_20),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_62),
.B2(n_78),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_45),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_23),
.B(n_45),
.C(n_78),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_37),
.B2(n_42),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_25),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_25),
.A2(n_43),
.B1(n_98),
.B2(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_30),
.B(n_75),
.C(n_77),
.Y(n_74)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_29),
.C(n_34),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_30),
.B1(n_52),
.B2(n_56),
.Y(n_57)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g196 ( 
.A(n_30),
.B(n_76),
.CON(n_196),
.SN(n_196)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_30),
.B(n_53),
.C(n_56),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_36),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_39),
.A2(n_75),
.B(n_76),
.Y(n_97)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_58),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_50),
.B1(n_61),
.B2(n_95),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_49),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_49),
.A2(n_51),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_50),
.A2(n_61),
.B1(n_196),
.B2(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_51)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_52),
.A2(n_54),
.B(n_196),
.C(n_197),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_54),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_54),
.B(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_61),
.B(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_74),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_63),
.B(n_74),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_65),
.A2(n_132),
.B(n_171),
.Y(n_220)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_68),
.B1(n_84),
.B2(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_68),
.B(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_71),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_107),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_69),
.A2(n_129),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_69),
.A2(n_170),
.B1(n_178),
.B2(n_184),
.Y(n_188)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_70),
.Y(n_171)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_70),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_76),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_76),
.B(n_87),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_79),
.A2(n_100),
.B1(n_101),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_79),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_94),
.C(n_96),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_80),
.A2(n_81),
.B1(n_94),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_88),
.B(n_90),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_82),
.A2(n_87),
.B1(n_109),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_82),
.A2(n_87),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_82),
.A2(n_87),
.B1(n_155),
.B2(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_82),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_89),
.B(n_93),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_93),
.A2(n_111),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_94),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_95),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_96),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_108),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_108),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_104),
.A2(n_131),
.B(n_168),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_138),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_125),
.B1(n_136),
.B2(n_137),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_133),
.B2(n_134),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_246),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_241),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_231),
.B(n_240),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_209),
.B(n_230),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_192),
.B(n_208),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_165),
.B(n_191),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_152),
.B1(n_153),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_175),
.B(n_190),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_186),
.B(n_189),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_207),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_207),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_202),
.C(n_205),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_206),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_222),
.B2(n_223),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_225),
.C(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_218),
.C(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_239),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);


endmodule