module fake_jpeg_5981_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_34),
.B1(n_29),
.B2(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_25),
.B1(n_33),
.B2(n_30),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_21),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_62),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_58),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_64),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_27),
.B1(n_17),
.B2(n_31),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_21),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_82),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_63),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_21),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_78),
.B(n_20),
.Y(n_117)
);

BUFx6f_ASAP7_75t_SL g72 ( 
.A(n_63),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

AND2x4_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_21),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_79),
.B(n_88),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_53),
.C(n_45),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_23),
.B(n_26),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_17),
.B(n_31),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_89),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_91),
.B1(n_25),
.B2(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_20),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_44),
.B1(n_32),
.B2(n_22),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_47),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_102),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_68),
.B1(n_64),
.B2(n_66),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_100),
.B1(n_76),
.B2(n_94),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_45),
.B(n_50),
.C(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_114),
.Y(n_136)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_106),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_76),
.B1(n_75),
.B2(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_74),
.B1(n_90),
.B2(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_110),
.Y(n_140)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_27),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_121),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_92),
.C(n_79),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_46),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_53),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_74),
.Y(n_127)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_138),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_86),
.B1(n_90),
.B2(n_78),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_125),
.B1(n_134),
.B2(n_139),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_91),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_91),
.B1(n_76),
.B2(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_143),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_116),
.C(n_112),
.Y(n_168)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_146),
.Y(n_171)
);

AOI31xp33_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_91),
.A3(n_84),
.B(n_73),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_139),
.C(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_92),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_120),
.B1(n_119),
.B2(n_114),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_31),
.B1(n_24),
.B2(n_45),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_150),
.B(n_151),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_165),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_159),
.C(n_32),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_R g158 ( 
.A(n_136),
.B(n_121),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_182),
.B(n_137),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_149),
.A3(n_124),
.B1(n_132),
.B2(n_134),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_160),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_108),
.B(n_111),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_166),
.B(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_106),
.B(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_111),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_183),
.C(n_182),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_46),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_26),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_174),
.Y(n_187)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_77),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_72),
.B1(n_85),
.B2(n_66),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_151),
.B1(n_150),
.B2(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_69),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_82),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_97),
.B(n_46),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_130),
.B1(n_138),
.B2(n_25),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_46),
.B(n_24),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_44),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_156),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_195),
.B1(n_200),
.B2(n_153),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_199),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_194),
.C(n_183),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_158),
.B(n_170),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_130),
.B1(n_47),
.B2(n_32),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_196),
.B(n_26),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_197),
.B(n_206),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_178),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_47),
.B1(n_32),
.B2(n_22),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_32),
.B1(n_26),
.B2(n_23),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_23),
.B1(n_26),
.B2(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_209),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_163),
.A2(n_26),
.B(n_23),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_176),
.B(n_162),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_210),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_220),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_229),
.B1(n_230),
.B2(n_234),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_221),
.C(n_232),
.Y(n_237)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_154),
.A3(n_156),
.B1(n_175),
.B2(n_179),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_168),
.C(n_165),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_225),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_175),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_199),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_198),
.A2(n_175),
.B(n_1),
.C(n_2),
.Y(n_229)
);

OAI22x1_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_173),
.B1(n_160),
.B2(n_180),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_207),
.B1(n_204),
.B2(n_26),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_184),
.C(n_209),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_200),
.Y(n_242)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_205),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_229),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_240),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_208),
.C(n_188),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_239),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_190),
.B(n_195),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_214),
.B1(n_218),
.B2(n_220),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_229),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_190),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_248),
.C(n_250),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_229),
.B1(n_1),
.B2(n_2),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_204),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_23),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_23),
.C(n_1),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_254),
.C(n_219),
.Y(n_259)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_0),
.C(n_1),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_255),
.B(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_262),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_267),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_260),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_248),
.B1(n_240),
.B2(n_236),
.Y(n_278)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_233),
.C(n_226),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_266),
.C(n_271),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_254),
.B1(n_246),
.B2(n_5),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_11),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_269),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_10),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_266),
.B(n_264),
.C(n_238),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_263),
.C(n_259),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_244),
.C(n_237),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_282),
.C(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_250),
.C(n_0),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_3),
.C(n_6),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_286),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_274),
.B1(n_273),
.B2(n_283),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_284),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_7),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_7),
.C(n_8),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_294),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_10),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_10),
.B(n_11),
.Y(n_295)
);

A2O1A1O1Ixp25_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_11),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_298),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_278),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_296),
.B1(n_291),
.B2(n_297),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_15),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_304),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_306),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_288),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_301),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_309),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.C(n_308),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_311),
.B(n_307),
.Y(n_315)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_16),
.C(n_313),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_16),
.Y(n_317)
);


endmodule