module real_jpeg_6656_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_0),
.A2(n_42),
.B1(n_47),
.B2(n_52),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_0),
.A2(n_52),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_0),
.A2(n_52),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_0),
.A2(n_52),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_1),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_1),
.A2(n_56),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_1),
.A2(n_56),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_1),
.A2(n_43),
.B1(n_56),
.B2(n_282),
.Y(n_281)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_3),
.A2(n_256),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_3),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_3),
.A2(n_301),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_3),
.A2(n_301),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_3),
.A2(n_301),
.B1(n_409),
.B2(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_4),
.B(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_4),
.A2(n_265),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_4),
.B(n_196),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_4),
.B(n_375),
.C(n_377),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_L g379 ( 
.A1(n_4),
.A2(n_380),
.B1(n_381),
.B2(n_383),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_4),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_4),
.B(n_152),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_4),
.A2(n_31),
.B1(n_320),
.B2(n_426),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_5),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_5),
.A2(n_286),
.B1(n_296),
.B2(n_312),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_5),
.A2(n_296),
.B1(n_383),
.B2(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_5),
.A2(n_296),
.B1(n_415),
.B2(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_7),
.A2(n_128),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_7),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_7),
.A2(n_67),
.B1(n_131),
.B2(n_188),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_7),
.A2(n_131),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_7),
.A2(n_131),
.B1(n_271),
.B2(n_274),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_115),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_8),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_8),
.A2(n_193),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_8),
.A2(n_193),
.B1(n_403),
.B2(n_406),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_8),
.A2(n_193),
.B1(n_383),
.B2(n_466),
.Y(n_465)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_10),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_10),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_12),
.Y(n_103)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_12),
.Y(n_263)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_15),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_15),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_15),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_15),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_15),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_15),
.Y(n_267)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_15),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_16),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_16),
.A2(n_87),
.B1(n_115),
.B2(n_121),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_16),
.A2(n_87),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_16),
.A2(n_87),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_510),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_500),
.B(n_509),
.Y(n_24)
);

OAI31xp33_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_225),
.A3(n_246),
.B(n_497),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_205),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_27),
.B(n_205),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_124),
.C(n_168),
.Y(n_27)
);

FAx1_ASAP7_75t_SL g365 ( 
.A(n_28),
.B(n_124),
.CI(n_168),
.CON(n_365),
.SN(n_365)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_91),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_29),
.A2(n_30),
.B(n_93),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_53),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_30),
.A2(n_92),
.B1(n_93),
.B2(n_123),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_30),
.A2(n_53),
.B1(n_92),
.B2(n_357),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_39),
.B(n_41),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_31),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_31),
.A2(n_269),
.B1(n_277),
.B2(n_281),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_31),
.A2(n_281),
.B(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_31),
.A2(n_180),
.B(n_402),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_31),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_31),
.A2(n_320),
.B1(n_414),
.B2(n_426),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_31),
.A2(n_41),
.B(n_318),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_34),
.Y(n_276)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_34),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g415 ( 
.A(n_34),
.Y(n_415)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_38),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_38),
.Y(n_435)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_41),
.Y(n_181)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_50),
.Y(n_428)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_51),
.Y(n_405)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_51),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_53),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_64),
.B(n_82),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_55),
.A2(n_65),
.B1(n_83),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_58),
.A2(n_90),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_59),
.Y(n_385)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_59),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_59),
.Y(n_450)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_60),
.Y(n_382)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_64),
.B(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_64),
.A2(n_160),
.B(n_161),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_64),
.A2(n_82),
.B(n_161),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_64),
.A2(n_160),
.B1(n_166),
.B2(n_187),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_64),
.A2(n_481),
.B(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_65),
.A2(n_83),
.B1(n_379),
.B2(n_386),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_65),
.A2(n_83),
.B1(n_386),
.B2(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_65),
.A2(n_83),
.B1(n_396),
.B2(n_465),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_76),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_75),
.Y(n_66)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_67),
.Y(n_373)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_74),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_75),
.Y(n_397)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_79),
.Y(n_273)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_90),
.Y(n_189)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_113),
.B(n_119),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_94),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_94),
.A2(n_196),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_94),
.A2(n_196),
.B1(n_293),
.B2(n_299),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_95),
.A2(n_192),
.B(n_195),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_95),
.A2(n_122),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_95),
.A2(n_122),
.B1(n_192),
.B2(n_300),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_95),
.A2(n_506),
.B(n_507),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_105),
.Y(n_312)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_112),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_115),
.Y(n_298)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_118),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_119),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_122),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_122),
.A2(n_216),
.B(n_221),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_158),
.B(n_167),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_125),
.B(n_158),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_136),
.B1(n_152),
.B2(n_153),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_127),
.A2(n_137),
.B(n_199),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g447 ( 
.A1(n_128),
.A2(n_448),
.A3(n_451),
.B1(n_454),
.B2(n_455),
.Y(n_447)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g463 ( 
.A1(n_129),
.A2(n_380),
.B(n_454),
.Y(n_463)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_130),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_130),
.Y(n_291)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_135),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_136),
.B(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_136),
.A2(n_153),
.B(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_136),
.A2(n_236),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_136),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_136),
.A2(n_152),
.B1(n_348),
.B2(n_463),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_136),
.A2(n_152),
.B(n_504),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_137),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_137),
.A2(n_311),
.B1(n_314),
.B2(n_315),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_137),
.A2(n_311),
.B1(n_314),
.B2(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_139),
.Y(n_457)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_142)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_143),
.Y(n_201)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_145),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_145),
.Y(n_261)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_145),
.Y(n_313)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g453 ( 
.A(n_147),
.Y(n_453)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_200),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_159),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_160),
.B(n_380),
.Y(n_424)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_163),
.Y(n_459)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_164),
.Y(n_469)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_167),
.B(n_206),
.CI(n_224),
.CON(n_205),
.SN(n_205)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_190),
.C(n_197),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_169),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_170),
.A2(n_184),
.B1(n_185),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_170),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_180),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_172),
.A2(n_270),
.B(n_343),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_173),
.Y(n_322)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_175),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_190),
.A2(n_191),
.B1(n_197),
.B2(n_198),
.Y(n_359)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_195),
.B(n_221),
.Y(n_512)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_203),
.B(n_380),
.Y(n_454)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_205),
.B(n_227),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_215),
.B2(n_223),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_214),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_209),
.B(n_233),
.C(n_241),
.Y(n_508)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_212),
.A2(n_237),
.B(n_314),
.Y(n_332)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_223),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_215),
.B(n_228),
.C(n_231),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_226),
.A2(n_498),
.B(n_499),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_241),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_237),
.Y(n_504)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_243),
.Y(n_506)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_366),
.B(n_491),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_351),
.C(n_363),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_336),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_249),
.A2(n_493),
.B(n_494),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_324),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_250),
.B(n_324),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_304),
.C(n_316),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_251),
.B(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_283),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_252),
.B(n_284),
.C(n_292),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_268),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_253),
.B(n_268),
.Y(n_339)
);

OAI32xp33_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_256),
.A3(n_258),
.B1(n_260),
.B2(n_264),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_282),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_292),
.Y(n_283)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_285),
.Y(n_315)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_304),
.B(n_316),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.C(n_310),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_305),
.B(n_306),
.CI(n_310),
.CON(n_338),
.SN(n_338)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_323),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

INVx3_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_327),
.C(n_329),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_334),
.C(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_335),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_349),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_337),
.B(n_349),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_338),
.B(n_489),
.Y(n_488)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_338),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_339),
.B(n_340),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.C(n_346),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_341),
.A2(n_342),
.B1(n_344),
.B2(n_345),
.Y(n_476)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_346),
.B(n_476),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

A2O1A1O1Ixp25_ASAP7_75t_L g491 ( 
.A1(n_351),
.A2(n_363),
.B(n_492),
.C(n_495),
.D(n_496),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_362),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_352),
.B(n_362),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_356),
.C(n_361),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_358),
.B1(n_360),
.B2(n_361),
.Y(n_355)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_356),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_358),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_364),
.B(n_365),
.Y(n_496)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_365),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_486),
.B(n_490),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_471),
.B(n_485),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_443),
.B(n_470),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_410),
.B(n_442),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_391),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_371),
.B(n_391),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_378),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_372),
.B(n_378),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_433),
.Y(n_432)
);

INVx3_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_390),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_401),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_394),
.B1(n_395),
.B2(n_400),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_400),
.C(n_401),
.Y(n_444)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_395),
.Y(n_400)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_402),
.Y(n_417)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_422),
.B(n_441),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_421),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_421),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_413),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_429),
.B(n_440),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_424),
.B(n_425),
.Y(n_440)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_436),
.Y(n_431)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx8_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx4_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_445),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_461),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_462),
.C(n_464),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_460),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_460),
.Y(n_479)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx11_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_464),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_465),
.Y(n_481)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_472),
.B(n_473),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_475),
.B1(n_477),
.B2(n_478),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_480),
.C(n_483),
.Y(n_487)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_479),
.A2(n_480),
.B1(n_483),
.B2(n_484),
.Y(n_478)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_479),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_480),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_487),
.B(n_488),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_502),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_502),
.B(n_512),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_502),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_503),
.B(n_505),
.CI(n_508),
.CON(n_502),
.SN(n_502)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_513),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_512),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);


endmodule