module fake_jpeg_19611_n_277 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_277);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx2_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

OAI22x1_ASAP7_75t_R g64 ( 
.A1(n_44),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_34),
.B1(n_16),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_67),
.B1(n_45),
.B2(n_21),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_16),
.B1(n_30),
.B2(n_14),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_47),
.Y(n_59)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_64),
.B(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_16),
.B1(n_33),
.B2(n_27),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

AND2x4_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_30),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_35),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_45),
.B1(n_38),
.B2(n_36),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_26),
.A3(n_16),
.B1(n_27),
.B2(n_31),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_62),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_76),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_40),
.B1(n_37),
.B2(n_45),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_73),
.B1(n_83),
.B2(n_50),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_28),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_80),
.C(n_85),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_35),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_35),
.C(n_29),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_38),
.B1(n_36),
.B2(n_20),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_35),
.C(n_29),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_68),
.B(n_87),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_89),
.B(n_91),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_62),
.B(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_61),
.B1(n_50),
.B2(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_96),
.B1(n_98),
.B2(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_101),
.B1(n_84),
.B2(n_75),
.Y(n_110)
);

OAI22x1_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_29),
.B1(n_28),
.B2(n_15),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_57),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_105),
.CI(n_78),
.CON(n_109),
.SN(n_109)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_55),
.B1(n_51),
.B2(n_58),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_58),
.B1(n_51),
.B2(n_65),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_79),
.B1(n_69),
.B2(n_81),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_58),
.B1(n_20),
.B2(n_21),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_106),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_29),
.C(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_117),
.B1(n_123),
.B2(n_125),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_114),
.B1(n_93),
.B2(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_87),
.B(n_77),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_119),
.B(n_18),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_87),
.B1(n_85),
.B2(n_69),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_121),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_74),
.B(n_1),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_74),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_18),
.B(n_2),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_127),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_79),
.B1(n_63),
.B2(n_21),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_126),
.B1(n_14),
.B2(n_23),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_89),
.A2(n_22),
.B1(n_42),
.B2(n_25),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_42),
.B1(n_13),
.B2(n_25),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_92),
.B(n_49),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_141),
.B1(n_144),
.B2(n_152),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_104),
.B(n_97),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_130),
.A2(n_139),
.B(n_145),
.Y(n_167)
);

INVxp33_ASAP7_75t_SL g132 ( 
.A(n_107),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_126),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_105),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_135),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_117),
.B(n_98),
.Y(n_135)
);

AOI22x1_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_97),
.B1(n_91),
.B2(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_91),
.B1(n_102),
.B2(n_14),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_24),
.A3(n_19),
.B1(n_18),
.B2(n_42),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_23),
.B1(n_24),
.B2(n_19),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_124),
.B1(n_119),
.B2(n_118),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_146),
.A2(n_150),
.B(n_15),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_15),
.B(n_18),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_15),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_24),
.B1(n_19),
.B2(n_18),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_120),
.B1(n_109),
.B2(n_122),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_157),
.B1(n_135),
.B2(n_141),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_148),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_120),
.B1(n_109),
.B2(n_108),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_125),
.C(n_123),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_174),
.C(n_151),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_170),
.B(n_145),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_18),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_115),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_155),
.A2(n_172),
.B1(n_175),
.B2(n_162),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_173),
.B1(n_165),
.B2(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_193),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_173),
.B1(n_168),
.B2(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_186),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_150),
.C(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_193),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_140),
.C(n_115),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_15),
.C(n_24),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_19),
.C(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_201),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_200),
.B(n_204),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_167),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_166),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_211),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_157),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_11),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_170),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_11),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_184),
.B(n_190),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_222),
.B(n_225),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_203),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_214),
.B1(n_223),
.B2(n_225),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_179),
.B(n_189),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_197),
.B(n_196),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_211),
.A2(n_181),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_0),
.C(n_2),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_229),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_3),
.B(n_4),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_3),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_242),
.B(n_238),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_236),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_5),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_202),
.B1(n_213),
.B2(n_210),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_238),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_201),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_241),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_4),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_4),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_224),
.B(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_216),
.C(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_216),
.C(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_248),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_7),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_237),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_6),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_6),
.C(n_7),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_252),
.B(n_246),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_253),
.C(n_10),
.Y(n_267)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_8),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_8),
.B(n_9),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_248),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_255),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.C(n_257),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_11),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_269),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_271),
.B(n_265),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_254),
.C(n_262),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_266),
.B(n_258),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_273),
.C(n_10),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_9),
.C(n_11),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_9),
.B(n_259),
.Y(n_277)
);


endmodule