module fake_jpeg_234_n_32 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_20),
.B1(n_11),
.B2(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_8),
.B(n_0),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_0),
.C(n_1),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_19),
.B1(n_10),
.B2(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_4),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_12),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_11),
.B1(n_12),
.B2(n_10),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_22),
.C(n_23),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.C(n_29),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_7),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_24),
.B(n_7),
.Y(n_31)
);

AOI321xp33_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_5),
.A3(n_7),
.B1(n_24),
.B2(n_27),
.C(n_30),
.Y(n_32)
);


endmodule