module fake_netlist_1_3234_n_15 (n_1, n_2, n_4, n_3, n_5, n_0, n_15);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_14;
wire n_10;
wire n_7;
wire n_8;
NAND2x1p5_ASAP7_75t_L g6 ( .A(n_1), .B(n_5), .Y(n_6) );
OR2x6_ASAP7_75t_L g7 ( .A(n_4), .B(n_0), .Y(n_7) );
AOI22xp33_ASAP7_75t_L g8 ( .A1(n_1), .A2(n_2), .B1(n_0), .B2(n_4), .Y(n_8) );
INVxp33_ASAP7_75t_L g9 ( .A(n_3), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
AOI22xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_10), .B1(n_11), .B2(n_7), .Y(n_14) );
OAI222xp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_2), .B1(n_3), .B2(n_7), .C1(n_8), .C2(n_6), .Y(n_15) );
endmodule