module fake_netlist_5_1563_n_2017 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2017);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2017;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_55),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_114),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_13),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_69),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_90),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_31),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_6),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_119),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_149),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_58),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_91),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_59),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_14),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_144),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_129),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_54),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_68),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_106),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_19),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_56),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_13),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_36),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_152),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_20),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_82),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_116),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_70),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_143),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_40),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_100),
.Y(n_233)
);

BUFx2_ASAP7_75t_SL g234 ( 
.A(n_69),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_181),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_19),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_63),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_95),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_120),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_65),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_53),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_3),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_167),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_154),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_62),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_59),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_50),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_170),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_125),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_63),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_161),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_164),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_98),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_112),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_93),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_0),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_8),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_75),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_123),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_68),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_131),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_50),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_135),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_30),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_52),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_132),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_180),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_74),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_175),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_128),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_49),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_71),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_65),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_166),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_121),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_88),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_57),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_54),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_3),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_107),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_177),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_92),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_30),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_110),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_18),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_60),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_22),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_124),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_163),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_56),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_146),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_89),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_96),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_182),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_85),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_103),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_35),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_145),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_58),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_39),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_102),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_52),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_43),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_72),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_80),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_47),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_21),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_86),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_2),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_1),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_37),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_29),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_159),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_118),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_2),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_11),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_94),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_7),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_61),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_49),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_66),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_17),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_37),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_39),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_1),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_138),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_158),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_51),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_78),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_122),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_179),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_12),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_140),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_185),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_47),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_162),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_44),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_61),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_51),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_111),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_81),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_151),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_84),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_189),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_97),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_62),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_31),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_12),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_171),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_44),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_46),
.Y(n_359)
);

BUFx10_ASAP7_75t_L g360 ( 
.A(n_101),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_28),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_104),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_64),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_117),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_28),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_187),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_109),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_24),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_33),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_73),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_150),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_4),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_53),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_15),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_137),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_115),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_184),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_5),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_24),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_64),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_242),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_215),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_215),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_284),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_194),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_284),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_292),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_292),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_252),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_265),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_274),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_231),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_193),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_247),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_299),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_236),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_240),
.Y(n_398)
);

BUFx6f_ASAP7_75t_SL g399 ( 
.A(n_203),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_243),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_219),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_315),
.B(n_0),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_312),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_350),
.B(n_4),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_219),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_342),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_248),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_219),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_235),
.B(n_5),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_251),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_357),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_362),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_229),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_254),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_219),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_219),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_226),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_269),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_233),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_226),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_270),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_226),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_276),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_238),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_235),
.B(n_6),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_246),
.B(n_7),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_247),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_226),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_239),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_226),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_245),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_249),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_211),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_245),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_244),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_245),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_245),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_245),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_277),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_253),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_307),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_198),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_255),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_249),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_279),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_307),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_246),
.B(n_257),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_283),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_307),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_307),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_256),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_288),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_259),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_249),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_307),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_257),
.B(n_8),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_263),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_285),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_297),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_266),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_305),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_221),
.B(n_9),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_271),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_327),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_303),
.B(n_9),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_275),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_310),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_314),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_327),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_327),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_318),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_434),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_434),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_327),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_438),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_438),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_327),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_419),
.B(n_329),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_408),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_408),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_421),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_420),
.B(n_329),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_329),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_410),
.B(n_329),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_440),
.Y(n_501)
);

NOR2x1_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_288),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_402),
.B(n_221),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_393),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_441),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_441),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_402),
.B(n_280),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_442),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_395),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_442),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_445),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_SL g517 ( 
.A(n_460),
.B(n_294),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_468),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_473),
.B(n_349),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_473),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_459),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_382),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_395),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_431),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_383),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_384),
.B(n_386),
.Y(n_533)
);

INVx6_ASAP7_75t_L g534 ( 
.A(n_406),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_387),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_388),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_389),
.B(n_349),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_429),
.B(n_329),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_409),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_411),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_430),
.B(n_199),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_446),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_413),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_469),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_404),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_437),
.B(n_367),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_398),
.B(n_199),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_394),
.A2(n_338),
.B(n_280),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_475),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_400),
.B(n_204),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_448),
.B(n_367),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_399),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_400),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_491),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_547),
.B(n_423),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_428),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_545),
.A2(n_417),
.B1(n_439),
.B2(n_433),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_499),
.B(n_348),
.C(n_304),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_407),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_550),
.B(n_444),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_SL g563 ( 
.A1(n_545),
.A2(n_399),
.B1(n_333),
.B2(n_369),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_550),
.B(n_447),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_522),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_522),
.Y(n_566)
);

AO22x2_ASAP7_75t_L g567 ( 
.A1(n_544),
.A2(n_294),
.B1(n_234),
.B2(n_241),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_530),
.B(n_414),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_544),
.A2(n_241),
.B1(n_264),
.B2(n_224),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_455),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_522),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_513),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_522),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_513),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_541),
.B(n_414),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_530),
.B(n_418),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_554),
.B(n_457),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_546),
.B(n_418),
.Y(n_581)
);

OAI21xp33_ASAP7_75t_L g582 ( 
.A1(n_538),
.A2(n_264),
.B(n_224),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_531),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_530),
.B(n_422),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_523),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_499),
.A2(n_340),
.B1(n_373),
.B2(n_380),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_513),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_503),
.B(n_422),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_513),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_542),
.B(n_461),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_523),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_546),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_511),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_513),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_513),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_477),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_496),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_496),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_530),
.B(n_425),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_523),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_523),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_553),
.B(n_464),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_553),
.B(n_467),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_549),
.B(n_436),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_492),
.Y(n_606)
);

BUFx8_ASAP7_75t_SL g607 ( 
.A(n_477),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_542),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_497),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_497),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_480),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_480),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_492),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_492),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_553),
.B(n_470),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_553),
.B(n_425),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_481),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_530),
.B(n_427),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_513),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_549),
.B(n_338),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_541),
.B(n_427),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_549),
.B(n_465),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_549),
.B(n_443),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_537),
.B(n_443),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_545),
.B(n_449),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_481),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_485),
.Y(n_627)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_503),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_494),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_538),
.A2(n_340),
.B1(n_373),
.B2(n_380),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_511),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_531),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_552),
.B(n_196),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_545),
.B(n_449),
.Y(n_635)
);

BUFx6f_ASAP7_75t_SL g636 ( 
.A(n_549),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_485),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_552),
.B(n_196),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_503),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_514),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_503),
.A2(n_308),
.B1(n_232),
.B2(n_237),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_549),
.B(n_452),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_487),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_487),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_531),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_549),
.B(n_452),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_549),
.B(n_462),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_514),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_495),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_529),
.B(n_462),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_503),
.A2(n_250),
.B1(n_260),
.B2(n_320),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_529),
.B(n_463),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_514),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_531),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_L g656 ( 
.A1(n_483),
.A2(n_488),
.B(n_502),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_531),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_514),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_551),
.B(n_463),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_SL g660 ( 
.A(n_489),
.B(n_471),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_495),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_494),
.Y(n_662)
);

INVx5_ASAP7_75t_L g663 ( 
.A(n_503),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_L g664 ( 
.A(n_488),
.B(n_192),
.C(n_191),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_486),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_529),
.B(n_471),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_529),
.B(n_472),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_486),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_551),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_531),
.B(n_472),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_494),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_500),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_500),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_503),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_514),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_510),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_531),
.B(n_475),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_500),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_477),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_500),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_510),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_551),
.B(n_458),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_503),
.A2(n_324),
.B1(n_358),
.B2(n_379),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_502),
.B(n_195),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_508),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_503),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_551),
.B(n_203),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_486),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_508),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_512),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_512),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_551),
.B(n_203),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_503),
.A2(n_261),
.B1(n_354),
.B2(n_378),
.Y(n_693)
);

NOR2x1p5_ASAP7_75t_L g694 ( 
.A(n_552),
.B(n_361),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_518),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_508),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_551),
.B(n_209),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_534),
.B(n_216),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_514),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_518),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_507),
.B(n_516),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_514),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_507),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_507),
.B(n_399),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_520),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_519),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_508),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_656),
.B(n_503),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_706),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_620),
.A2(n_509),
.B1(n_548),
.B2(n_517),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_593),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_620),
.A2(n_509),
.B1(n_548),
.B2(n_517),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_590),
.A2(n_416),
.B1(n_385),
.B2(n_415),
.Y(n_714)
);

NOR3xp33_ASAP7_75t_L g715 ( 
.A(n_558),
.B(n_701),
.C(n_660),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_656),
.B(n_509),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_611),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_706),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_621),
.B(n_509),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_611),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_592),
.B(n_509),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_612),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_592),
.B(n_509),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_620),
.B(n_516),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_555),
.B(n_577),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_669),
.A2(n_577),
.B1(n_597),
.B2(n_555),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_597),
.B(n_509),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_598),
.B(n_509),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_569),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_598),
.B(n_509),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_669),
.B(n_516),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_625),
.B(n_489),
.Y(n_732)
);

INVx8_ASAP7_75t_L g733 ( 
.A(n_628),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_635),
.B(n_490),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_632),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_632),
.B(n_490),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_593),
.B(n_505),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_609),
.B(n_509),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_609),
.B(n_509),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_578),
.A2(n_642),
.B1(n_646),
.B2(n_616),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_612),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_650),
.B(n_390),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_610),
.B(n_548),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_694),
.B(n_533),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_617),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_653),
.B(n_391),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_639),
.B(n_539),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_617),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_639),
.B(n_663),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_626),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_556),
.B(n_392),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_639),
.B(n_539),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_610),
.B(n_535),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_557),
.B(n_396),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_626),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_608),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_666),
.B(n_535),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_627),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_639),
.B(n_539),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_667),
.B(n_535),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_562),
.B(n_403),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_561),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_582),
.A2(n_483),
.B(n_532),
.C(n_528),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_627),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_637),
.B(n_535),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_637),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_643),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_643),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_644),
.B(n_535),
.Y(n_769)
);

INVx4_ASAP7_75t_L g770 ( 
.A(n_628),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_628),
.B(n_205),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_639),
.B(n_539),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_644),
.B(n_649),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_569),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_639),
.B(n_539),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_649),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_628),
.B(n_205),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_661),
.B(n_539),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_661),
.B(n_539),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_694),
.B(n_533),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_676),
.B(n_539),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_676),
.B(n_519),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_704),
.B(n_505),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_561),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_681),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_681),
.Y(n_786)
);

INVxp33_ASAP7_75t_L g787 ( 
.A(n_581),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_559),
.B(n_532),
.C(n_537),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_569),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_559),
.A2(n_519),
.B1(n_301),
.B2(n_273),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_581),
.B(n_533),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_690),
.B(n_519),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_691),
.B(n_519),
.Y(n_794)
);

OR2x6_ASAP7_75t_L g795 ( 
.A(n_698),
.B(n_534),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_691),
.B(n_519),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_564),
.B(n_534),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_624),
.B(n_537),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_663),
.B(n_196),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_624),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_695),
.B(n_476),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_679),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_695),
.B(n_476),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_602),
.B(n_540),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_663),
.B(n_196),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_700),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_568),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_603),
.B(n_540),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_700),
.B(n_476),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_705),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_705),
.B(n_476),
.Y(n_811)
);

NAND2x1p5_ASAP7_75t_L g812 ( 
.A(n_663),
.B(n_218),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_579),
.B(n_476),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_565),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_584),
.B(n_478),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_615),
.B(n_534),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_582),
.A2(n_330),
.B(n_290),
.C(n_311),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_707),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_707),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_572),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_565),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_566),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_663),
.B(n_196),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_605),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_569),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_599),
.B(n_534),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_566),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_618),
.B(n_478),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_623),
.A2(n_647),
.B1(n_698),
.B2(n_684),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_670),
.B(n_478),
.Y(n_830)
);

AND2x4_ASAP7_75t_SL g831 ( 
.A(n_698),
.B(n_209),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_588),
.A2(n_337),
.B1(n_322),
.B2(n_227),
.Y(n_832)
);

INVx8_ASAP7_75t_L g833 ( 
.A(n_628),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_573),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_677),
.B(n_478),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_573),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_580),
.B(n_543),
.C(n_528),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_682),
.B(n_536),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_633),
.B(n_478),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_663),
.B(n_200),
.Y(n_840)
);

INVxp33_ASAP7_75t_L g841 ( 
.A(n_596),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_703),
.B(n_534),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_659),
.B(n_536),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_605),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_674),
.B(n_200),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_655),
.B(n_482),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_563),
.B(n_543),
.C(n_528),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_569),
.B(n_482),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_607),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_606),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_567),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_674),
.B(n_200),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_606),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_665),
.B(n_482),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_665),
.B(n_482),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_665),
.B(n_482),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_665),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_665),
.B(n_484),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_668),
.B(n_688),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_674),
.B(n_200),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_641),
.A2(n_262),
.B1(n_268),
.B2(n_375),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_560),
.A2(n_479),
.B(n_484),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_668),
.B(n_484),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_575),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_604),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_668),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_668),
.B(n_484),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_613),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_567),
.B(n_536),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_613),
.Y(n_870)
);

NOR2xp67_ASAP7_75t_SL g871 ( 
.A(n_674),
.B(n_686),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_674),
.B(n_200),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_668),
.B(n_484),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_674),
.B(n_334),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_622),
.B(n_258),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_688),
.B(n_520),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_575),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_688),
.B(n_498),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_708),
.A2(n_645),
.B(n_560),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_802),
.B(n_664),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_825),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_717),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_SL g883 ( 
.A(n_820),
.B(n_703),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_716),
.A2(n_645),
.B(n_560),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_725),
.B(n_687),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_740),
.A2(n_726),
.B1(n_724),
.B2(n_829),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_875),
.A2(n_697),
.B(n_692),
.C(n_664),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_748),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_748),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_804),
.B(n_688),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_756),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_733),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_724),
.A2(n_636),
.B1(n_698),
.B2(n_652),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_770),
.B(n_686),
.Y(n_894)
);

AND2x2_ASAP7_75t_SL g895 ( 
.A(n_751),
.B(n_571),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_733),
.Y(n_896)
);

AO21x1_ASAP7_75t_L g897 ( 
.A1(n_743),
.A2(n_281),
.B(n_278),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_830),
.A2(n_835),
.B(n_728),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_750),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_712),
.B(n_686),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_750),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_770),
.A2(n_657),
.B(n_645),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_734),
.B(n_567),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_784),
.A2(n_636),
.B1(n_698),
.B2(n_693),
.Y(n_904)
);

OAI21xp33_ASAP7_75t_L g905 ( 
.A1(n_732),
.A2(n_737),
.B(n_787),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_770),
.A2(n_657),
.B(n_686),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_688),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_859),
.A2(n_657),
.B(n_686),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_804),
.B(n_567),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_712),
.B(n_686),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_800),
.A2(n_719),
.B1(n_760),
.B2(n_757),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_762),
.A2(n_636),
.B1(n_683),
.B2(n_583),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_733),
.A2(n_640),
.B(n_594),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_762),
.A2(n_583),
.B1(n_634),
.B2(n_638),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_833),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_808),
.B(n_570),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_808),
.B(n_570),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_727),
.A2(n_291),
.B(n_287),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_833),
.A2(n_640),
.B(n_594),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_807),
.B(n_570),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_833),
.A2(n_640),
.B(n_594),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_833),
.A2(n_640),
.B(n_594),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_720),
.B(n_570),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_798),
.B(n_631),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_787),
.B(n_267),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_722),
.B(n_574),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_862),
.A2(n_576),
.B(n_574),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_825),
.Y(n_928)
);

O2A1O1Ixp5_ASAP7_75t_L g929 ( 
.A1(n_773),
.A2(n_702),
.B(n_699),
.C(n_595),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_730),
.A2(n_300),
.B(n_293),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_SL g931 ( 
.A1(n_738),
.A2(n_377),
.B(n_371),
.C(n_352),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_798),
.B(n_586),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_800),
.A2(n_272),
.B1(n_583),
.B2(n_376),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_774),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_758),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_729),
.A2(n_866),
.B(n_815),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_741),
.B(n_574),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_739),
.A2(n_629),
.B(n_614),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_813),
.A2(n_658),
.B(n_576),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_745),
.B(n_574),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_755),
.B(n_576),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_766),
.B(n_767),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_721),
.A2(n_629),
.B(n_614),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_776),
.B(n_576),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_785),
.B(n_587),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_832),
.A2(n_583),
.B1(n_204),
.B2(n_376),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_793),
.B(n_587),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_806),
.B(n_587),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_L g949 ( 
.A(n_774),
.B(n_634),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_828),
.A2(n_658),
.B(n_589),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_753),
.A2(n_346),
.B(n_319),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_710),
.A2(n_206),
.B1(n_366),
.B2(n_364),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_736),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_774),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_797),
.B(n_206),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_764),
.B(n_587),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_869),
.B(n_589),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_735),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_768),
.B(n_589),
.Y(n_959)
);

AO21x1_ASAP7_75t_L g960 ( 
.A1(n_826),
.A2(n_365),
.B(n_585),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_851),
.A2(n_671),
.B(n_630),
.C(n_696),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_768),
.A2(n_702),
.B(n_699),
.C(n_589),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_786),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_723),
.A2(n_792),
.B(n_782),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_786),
.B(n_595),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_843),
.A2(n_763),
.B(n_788),
.C(n_791),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_791),
.B(n_305),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_810),
.B(n_595),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_810),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_713),
.A2(n_207),
.B1(n_366),
.B2(n_364),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_816),
.B(n_595),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_744),
.B(n_207),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_774),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_869),
.B(n_619),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_851),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_865),
.A2(n_702),
.B(n_699),
.C(n_619),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_L g977 ( 
.A(n_754),
.B(n_213),
.C(n_210),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_742),
.B(n_619),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_714),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_794),
.A2(n_796),
.B(n_777),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_746),
.B(n_619),
.Y(n_981)
);

BUFx8_ASAP7_75t_L g982 ( 
.A(n_744),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_771),
.A2(n_658),
.B(n_651),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_709),
.B(n_711),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_744),
.B(n_210),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_718),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_731),
.A2(n_671),
.B(n_630),
.C(n_696),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_771),
.A2(n_658),
.B(n_651),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_780),
.B(n_648),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_761),
.B(n_213),
.Y(n_990)
);

AO21x1_ASAP7_75t_L g991 ( 
.A1(n_778),
.A2(n_591),
.B(n_585),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_865),
.B(n_214),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_780),
.B(n_731),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_789),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_777),
.A2(n_651),
.B(n_648),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_839),
.A2(n_651),
.B(n_648),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_842),
.B(n_214),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_838),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_780),
.B(n_222),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_789),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_783),
.B(n_222),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_818),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_715),
.A2(n_197),
.B(n_193),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_847),
.B(n_648),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_837),
.B(n_225),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_789),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_801),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_790),
.B(n_654),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_846),
.A2(n_699),
.B(n_654),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_817),
.A2(n_286),
.B(n_223),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_848),
.A2(n_702),
.B(n_654),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_831),
.B(n_225),
.Y(n_1012)
);

NOR2xp67_ASAP7_75t_L g1013 ( 
.A(n_803),
.B(n_282),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_809),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_795),
.A2(n_353),
.B1(n_230),
.B2(n_335),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_824),
.B(n_654),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_854),
.A2(n_675),
.B(n_600),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_831),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_765),
.A2(n_769),
.B(n_811),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_789),
.B(n_228),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_855),
.A2(n_675),
.B(n_600),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_824),
.B(n_675),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_844),
.B(n_675),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_844),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_856),
.A2(n_689),
.B(n_685),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_858),
.A2(n_591),
.B(n_601),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_795),
.B(n_228),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_818),
.A2(n_819),
.B(n_850),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_863),
.A2(n_601),
.B(n_685),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_779),
.A2(n_689),
.B(n_680),
.C(n_678),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_819),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_795),
.B(n_230),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_781),
.A2(n_680),
.B(n_678),
.C(n_673),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_857),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_850),
.B(n_662),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_795),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_817),
.A2(n_673),
.B(n_672),
.C(n_662),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_867),
.A2(n_672),
.B(n_479),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_876),
.A2(n_638),
.B1(n_634),
.B2(n_289),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_853),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_799),
.A2(n_527),
.B(n_526),
.C(n_525),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_853),
.B(n_634),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_868),
.B(n_634),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_868),
.B(n_634),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_814),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_870),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_857),
.B(n_335),
.Y(n_1047)
);

BUFx4f_ASAP7_75t_L g1048 ( 
.A(n_821),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_841),
.B(n_209),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_873),
.A2(n_479),
.B(n_493),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_799),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_870),
.A2(n_638),
.B(n_634),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_857),
.B(n_341),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_861),
.A2(n_638),
.B1(n_370),
.B2(n_334),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_822),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_878),
.A2(n_479),
.B(n_493),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_827),
.B(n_638),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_834),
.B(n_341),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_749),
.A2(n_493),
.B(n_504),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_749),
.A2(n_493),
.B(n_504),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_836),
.B(n_525),
.Y(n_1061)
);

OAI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_864),
.A2(n_202),
.B(n_197),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_812),
.B(n_334),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_877),
.B(n_805),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_747),
.A2(n_493),
.B(n_504),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_874),
.A2(n_526),
.B(n_527),
.C(n_515),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_747),
.A2(n_504),
.B(n_521),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_895),
.B(n_993),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_993),
.B(n_344),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_SL g1070 ( 
.A(n_883),
.B(n_841),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_958),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_905),
.B(n_885),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_907),
.A2(n_752),
.B(n_759),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1034),
.A2(n_752),
.B(n_759),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1036),
.B(n_772),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_982),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_882),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_990),
.B(n_849),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_891),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_887),
.A2(n_874),
.B(n_872),
.C(n_860),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1034),
.A2(n_772),
.B(n_775),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_953),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_934),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_980),
.A2(n_775),
.B(n_823),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_880),
.B(n_344),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_932),
.B(n_805),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_980),
.A2(n_812),
.B(n_871),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_913),
.A2(n_872),
.B(n_860),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_982),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_979),
.B(n_849),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_SL g1091 ( 
.A(n_1003),
.B(n_202),
.C(n_374),
.Y(n_1091)
);

CKINVDCx10_ASAP7_75t_R g1092 ( 
.A(n_1049),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_886),
.A2(n_852),
.B(n_845),
.C(n_840),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_998),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_934),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_881),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_975),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1002),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_967),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_888),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1048),
.B(n_351),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_1036),
.B(n_823),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_992),
.B(n_323),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_919),
.A2(n_852),
.B(n_845),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_977),
.A2(n_506),
.B(n_501),
.C(n_498),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_SL g1106 ( 
.A(n_1018),
.Y(n_1106)
);

AOI22x1_ASAP7_75t_L g1107 ( 
.A1(n_964),
.A2(n_898),
.B1(n_1014),
.B2(n_1007),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_921),
.A2(n_840),
.B(n_334),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1048),
.B(n_351),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_964),
.A2(n_638),
.B(n_498),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_909),
.A2(n_372),
.B1(n_286),
.B2(n_223),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1045),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_942),
.B(n_989),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_924),
.B(n_353),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_925),
.B(n_1012),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_922),
.A2(n_334),
.B(n_370),
.Y(n_1116)
);

NOR2x1_ASAP7_75t_L g1117 ( 
.A(n_1006),
.B(n_954),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_997),
.B(n_295),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_966),
.A2(n_374),
.B1(n_372),
.B2(n_363),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_936),
.A2(n_370),
.B(n_296),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_971),
.A2(n_370),
.B(n_298),
.Y(n_1121)
);

AO21x2_ASAP7_75t_L g1122 ( 
.A1(n_960),
.A2(n_515),
.B(n_506),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_SL g1123 ( 
.A(n_972),
.B(n_363),
.C(n_220),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_934),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1027),
.B(n_302),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_957),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1001),
.B(n_328),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_957),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1031),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_889),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_903),
.B(n_201),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1004),
.A2(n_957),
.B1(n_951),
.B2(n_986),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_985),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_899),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_L g1135 ( 
.A1(n_897),
.A2(n_515),
.B(n_506),
.C(n_501),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_L g1136 ( 
.A1(n_955),
.A2(n_501),
.B(n_521),
.C(n_504),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_999),
.B(n_201),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_L g1138 ( 
.A(n_1032),
.B(n_332),
.C(n_212),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_954),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_L g1140 ( 
.A1(n_991),
.A2(n_918),
.B(n_911),
.C(n_978),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_898),
.A2(n_638),
.B(n_521),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_890),
.A2(n_370),
.B(n_306),
.Y(n_1142)
);

INVx6_ASAP7_75t_L g1143 ( 
.A(n_994),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1047),
.B(n_313),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1062),
.B(n_305),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_963),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_981),
.B(n_208),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_973),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_901),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_916),
.B(n_521),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_SL g1151 ( 
.A(n_1010),
.B(n_332),
.C(n_208),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_920),
.B(n_212),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_881),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_917),
.B(n_521),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_892),
.B(n_524),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1058),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_935),
.B(n_316),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_R g1158 ( 
.A(n_973),
.B(n_321),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_994),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_983),
.A2(n_325),
.B(n_524),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_SL g1161 ( 
.A1(n_1053),
.A2(n_309),
.B(n_360),
.C(n_339),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1005),
.B(n_343),
.C(n_217),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_893),
.A2(n_343),
.B1(n_359),
.B2(n_356),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_983),
.A2(n_524),
.B(n_126),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1015),
.B(n_217),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_912),
.A2(n_345),
.B1(n_359),
.B2(n_356),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_988),
.A2(n_524),
.B(n_83),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1004),
.A2(n_345),
.B(n_220),
.C(n_336),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_928),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_931),
.A2(n_309),
.B(n_339),
.C(n_360),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_L g1171 ( 
.A(n_1020),
.B(n_331),
.C(n_336),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_988),
.A2(n_524),
.B(n_76),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_952),
.A2(n_309),
.B(n_339),
.C(n_360),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_957),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_984),
.B(n_347),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_892),
.B(n_524),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_969),
.A2(n_974),
.B1(n_904),
.B2(n_1008),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1061),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_957),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1061),
.B(n_368),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1024),
.B(n_1040),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1046),
.B(n_205),
.Y(n_1182)
);

INVx6_ASAP7_75t_L g1183 ( 
.A(n_1000),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_894),
.A2(n_524),
.B(n_169),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1000),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_933),
.B(n_347),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_894),
.A2(n_524),
.B(n_168),
.Y(n_1187)
);

NAND2x1p5_ASAP7_75t_L g1188 ( 
.A(n_896),
.B(n_148),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_915),
.A2(n_153),
.B(n_87),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_915),
.B(n_331),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_928),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1055),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_915),
.A2(n_173),
.B(n_190),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_970),
.B(n_368),
.Y(n_1194)
);

OAI21xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1051),
.A2(n_1064),
.B(n_926),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_923),
.B(n_10),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_896),
.B(n_915),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1063),
.Y(n_1198)
);

NOR3xp33_ASAP7_75t_SL g1199 ( 
.A(n_946),
.B(n_368),
.C(n_16),
.Y(n_1199)
);

AOI22x1_ASAP7_75t_L g1200 ( 
.A1(n_996),
.A2(n_205),
.B1(n_188),
.B2(n_183),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_995),
.A2(n_141),
.B(n_178),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1019),
.B(n_205),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_937),
.B(n_205),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_940),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_941),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_944),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1013),
.B(n_205),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_945),
.B(n_205),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_947),
.B(n_176),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_995),
.A2(n_174),
.B(n_147),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_930),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_879),
.A2(n_884),
.B(n_1026),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_902),
.A2(n_139),
.B(n_134),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_948),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_956),
.B(n_130),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_959),
.B(n_127),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_965),
.B(n_79),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1035),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_939),
.A2(n_18),
.B(n_20),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_950),
.A2(n_21),
.B(n_22),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1016),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_968),
.B(n_1028),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_900),
.Y(n_1223)
);

INVx3_ASAP7_75t_SL g1224 ( 
.A(n_1063),
.Y(n_1224)
);

AND2x6_ASAP7_75t_SL g1225 ( 
.A(n_1063),
.B(n_23),
.Y(n_1225)
);

OAI22x1_ASAP7_75t_L g1226 ( 
.A1(n_914),
.A2(n_910),
.B1(n_1039),
.B2(n_1057),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_1022),
.Y(n_1227)
);

INVx1_ASAP7_75t_SL g1228 ( 
.A(n_1082),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1212),
.A2(n_1025),
.B(n_929),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1093),
.A2(n_976),
.B(n_1033),
.C(n_1030),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1087),
.A2(n_906),
.B(n_884),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1077),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1195),
.A2(n_879),
.B(n_908),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1088),
.A2(n_943),
.B(n_996),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1104),
.A2(n_1009),
.B(n_938),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1103),
.B(n_1041),
.C(n_1066),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_SL g1237 ( 
.A1(n_1080),
.A2(n_1217),
.B(n_1068),
.C(n_1086),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1194),
.B(n_961),
.C(n_987),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1099),
.B(n_1023),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1071),
.B(n_1043),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_1185),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1084),
.A2(n_1017),
.B(n_1021),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1115),
.B(n_1054),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1177),
.A2(n_1009),
.A3(n_1026),
.B(n_1017),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_1156),
.B(n_1011),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1197),
.B(n_927),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1112),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1222),
.A2(n_1107),
.B(n_1084),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1140),
.A2(n_962),
.B(n_1029),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1147),
.B(n_1011),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1095),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1177),
.A2(n_1029),
.B(n_1038),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1202),
.A2(n_1038),
.B(n_1021),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1100),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1132),
.A2(n_1042),
.B1(n_1044),
.B2(n_1052),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1186),
.A2(n_949),
.B1(n_1065),
.B2(n_1067),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1070),
.B(n_1060),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1073),
.A2(n_1037),
.B(n_1056),
.Y(n_1258)
);

CKINVDCx11_ASAP7_75t_R g1259 ( 
.A(n_1076),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_SL g1260 ( 
.A1(n_1086),
.A2(n_1065),
.B(n_1067),
.C(n_1060),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_SL g1261 ( 
.A1(n_1105),
.A2(n_1059),
.B(n_1050),
.C(n_1056),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1164),
.A2(n_1050),
.B(n_1059),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1130),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1078),
.B(n_23),
.Y(n_1264)
);

AOI221xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1119),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.C(n_29),
.Y(n_1265)
);

NOR2x1_ASAP7_75t_R g1266 ( 
.A(n_1089),
.B(n_1079),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1152),
.B(n_25),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1185),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1214),
.B(n_1175),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1141),
.A2(n_26),
.B(n_27),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1090),
.B(n_32),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1094),
.B(n_32),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1131),
.B(n_34),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1127),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1141),
.A2(n_38),
.B(n_40),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1173),
.A2(n_38),
.B(n_41),
.C(n_42),
.Y(n_1276)
);

NOR2xp67_ASAP7_75t_SL g1277 ( 
.A(n_1185),
.B(n_41),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1167),
.A2(n_42),
.B(n_45),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1165),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1197),
.Y(n_1280)
);

AOI31xp67_ASAP7_75t_L g1281 ( 
.A1(n_1202),
.A2(n_48),
.A3(n_57),
.B(n_60),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1134),
.A2(n_66),
.B1(n_67),
.B2(n_1149),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1172),
.A2(n_67),
.B(n_1209),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1209),
.A2(n_1072),
.B(n_1215),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1119),
.A2(n_1163),
.B1(n_1137),
.B2(n_1166),
.C(n_1111),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1192),
.B(n_1138),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_L g1287 ( 
.A(n_1199),
.B(n_1091),
.C(n_1170),
.Y(n_1287)
);

INVx3_ASAP7_75t_SL g1288 ( 
.A(n_1224),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1178),
.B(n_1133),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1110),
.A2(n_1135),
.B(n_1203),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1097),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1110),
.A2(n_1154),
.B(n_1150),
.Y(n_1292)
);

AOI221x1_ASAP7_75t_L g1293 ( 
.A1(n_1219),
.A2(n_1220),
.B1(n_1163),
.B2(n_1116),
.C(n_1226),
.Y(n_1293)
);

AOI31xp67_ASAP7_75t_L g1294 ( 
.A1(n_1207),
.A2(n_1208),
.A3(n_1203),
.B(n_1182),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1174),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1215),
.A2(n_1216),
.B(n_1074),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1162),
.A2(n_1114),
.B(n_1151),
.C(n_1171),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_SL g1298 ( 
.A1(n_1216),
.A2(n_1168),
.B(n_1161),
.C(n_1144),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1106),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1095),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1227),
.B(n_1218),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1180),
.B(n_1145),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1150),
.A2(n_1154),
.B(n_1182),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1095),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1081),
.A2(n_1176),
.B(n_1205),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1206),
.B(n_1111),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1069),
.B(n_1085),
.Y(n_1307)
);

AOI211x1_ASAP7_75t_L g1308 ( 
.A1(n_1166),
.A2(n_1181),
.B(n_1157),
.C(n_1125),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1124),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1160),
.A2(n_1187),
.B(n_1184),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1108),
.A2(n_1181),
.B(n_1210),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1075),
.B(n_1174),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1176),
.A2(n_1113),
.B(n_1201),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1123),
.B(n_1146),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1221),
.B(n_1113),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1176),
.A2(n_1113),
.B(n_1213),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1136),
.A2(n_1155),
.B(n_1200),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1225),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1118),
.B(n_1101),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1196),
.A2(n_1157),
.B1(n_1128),
.B2(n_1126),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1204),
.B(n_1129),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1109),
.B(n_1098),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_SL g1323 ( 
.A(n_1211),
.B(n_1158),
.C(n_1190),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1174),
.B(n_1179),
.Y(n_1324)
);

AOI31xp67_ASAP7_75t_L g1325 ( 
.A1(n_1122),
.A2(n_1102),
.A3(n_1075),
.B(n_1120),
.Y(n_1325)
);

INVxp67_ASAP7_75t_SL g1326 ( 
.A(n_1096),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1198),
.B(n_1102),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1204),
.A2(n_1198),
.B1(n_1223),
.B2(n_1179),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1121),
.A2(n_1142),
.B(n_1193),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1153),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1189),
.A2(n_1117),
.B(n_1122),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1179),
.B(n_1204),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1153),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1083),
.A2(n_1159),
.A3(n_1139),
.B(n_1155),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1169),
.B(n_1191),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1188),
.A2(n_1083),
.B(n_1159),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1139),
.A2(n_1188),
.B(n_1223),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1148),
.A2(n_1143),
.B(n_1183),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1148),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1124),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1143),
.A2(n_1183),
.B(n_1092),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1147),
.B(n_734),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1087),
.A2(n_770),
.B(n_907),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1068),
.A2(n_820),
.B1(n_740),
.B2(n_885),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1087),
.A2(n_770),
.B(n_907),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1177),
.A2(n_897),
.A3(n_960),
.B(n_991),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1147),
.B(n_734),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1087),
.A2(n_770),
.B(n_907),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1103),
.A2(n_886),
.B1(n_1220),
.B2(n_1219),
.C(n_990),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1103),
.A2(n_1115),
.B(n_875),
.C(n_990),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1147),
.B(n_734),
.Y(n_1351)
);

AO32x2_ASAP7_75t_L g1352 ( 
.A1(n_1177),
.A2(n_886),
.A3(n_1111),
.B1(n_1119),
.B2(n_1163),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1197),
.B(n_1036),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1147),
.B(n_734),
.Y(n_1354)
);

OAI22x1_ASAP7_75t_L g1355 ( 
.A1(n_1115),
.A2(n_1194),
.B1(n_820),
.B2(n_1103),
.Y(n_1355)
);

AO31x2_ASAP7_75t_L g1356 ( 
.A1(n_1177),
.A2(n_897),
.A3(n_960),
.B(n_991),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1068),
.A2(n_820),
.B1(n_740),
.B2(n_885),
.Y(n_1357)
);

NAND3x1_ASAP7_75t_L g1358 ( 
.A(n_1165),
.B(n_715),
.C(n_751),
.Y(n_1358)
);

INVx3_ASAP7_75t_SL g1359 ( 
.A(n_1076),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1147),
.B(n_734),
.Y(n_1360)
);

OAI22x1_ASAP7_75t_L g1361 ( 
.A1(n_1115),
.A2(n_1194),
.B1(n_820),
.B2(n_1103),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1112),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1077),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1087),
.A2(n_770),
.B(n_907),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1212),
.A2(n_1025),
.B(n_1087),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1103),
.A2(n_1115),
.B(n_875),
.C(n_990),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1140),
.A2(n_886),
.B(n_964),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1087),
.A2(n_770),
.B(n_907),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1177),
.A2(n_897),
.A3(n_960),
.B(n_991),
.Y(n_1369)
);

NOR2x1_ASAP7_75t_R g1370 ( 
.A(n_1089),
.B(n_703),
.Y(n_1370)
);

BUFx5_ASAP7_75t_L g1371 ( 
.A(n_1197),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1103),
.A2(n_1115),
.B(n_875),
.C(n_990),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1103),
.A2(n_1115),
.B(n_875),
.C(n_990),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1095),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1087),
.A2(n_770),
.B(n_907),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_SL g1376 ( 
.A1(n_1093),
.A2(n_887),
.B(n_966),
.C(n_724),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1212),
.A2(n_1025),
.B(n_1087),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1147),
.B(n_734),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1103),
.B(n_990),
.C(n_734),
.Y(n_1379)
);

BUFx8_ASAP7_75t_SL g1380 ( 
.A(n_1079),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_SL g1381 ( 
.A1(n_1093),
.A2(n_887),
.B(n_966),
.C(n_724),
.Y(n_1381)
);

AO21x1_ASAP7_75t_L g1382 ( 
.A1(n_1177),
.A2(n_886),
.B(n_740),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1103),
.A2(n_820),
.B(n_990),
.C(n_734),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1095),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1212),
.A2(n_1222),
.B(n_1202),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_1097),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1140),
.A2(n_886),
.B(n_964),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1178),
.B(n_1112),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1228),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1302),
.B(n_1269),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1342),
.B(n_1347),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1285),
.A2(n_1379),
.B1(n_1360),
.B2(n_1351),
.Y(n_1392)
);

CKINVDCx6p67_ASAP7_75t_R g1393 ( 
.A(n_1359),
.Y(n_1393)
);

BUFx10_ASAP7_75t_L g1394 ( 
.A(n_1388),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1379),
.A2(n_1366),
.B1(n_1350),
.B2(n_1372),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1354),
.A2(n_1378),
.B1(n_1267),
.B2(n_1273),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1367),
.A2(n_1387),
.B(n_1252),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1373),
.B(n_1383),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1315),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1358),
.A2(n_1297),
.B1(n_1307),
.B2(n_1228),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1254),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1314),
.B(n_1264),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1280),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1241),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1259),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1301),
.B(n_1306),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1362),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1241),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1247),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1263),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1388),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1279),
.A2(n_1271),
.B1(n_1382),
.B2(n_1355),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1288),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1279),
.A2(n_1361),
.B1(n_1287),
.B2(n_1323),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1268),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1268),
.Y(n_1416)
);

INVx4_ASAP7_75t_L g1417 ( 
.A(n_1251),
.Y(n_1417)
);

CKINVDCx11_ASAP7_75t_R g1418 ( 
.A(n_1318),
.Y(n_1418)
);

OAI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1282),
.A2(n_1287),
.B1(n_1349),
.B2(n_1357),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1380),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1251),
.Y(n_1421)
);

OAI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1282),
.A2(n_1344),
.B1(n_1243),
.B2(n_1239),
.Y(n_1422)
);

BUFx4f_ASAP7_75t_SL g1423 ( 
.A(n_1299),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1319),
.A2(n_1257),
.B1(n_1320),
.B2(n_1245),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1247),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1367),
.A2(n_1387),
.B1(n_1272),
.B2(n_1265),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1327),
.B(n_1240),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1286),
.A2(n_1289),
.B1(n_1277),
.B2(n_1312),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1291),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1251),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1363),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1265),
.A2(n_1236),
.B1(n_1352),
.B2(n_1250),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1386),
.A2(n_1328),
.B1(n_1322),
.B2(n_1236),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1321),
.B(n_1312),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1238),
.A2(n_1283),
.B1(n_1352),
.B2(n_1284),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1309),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1328),
.A2(n_1293),
.B1(n_1238),
.B2(n_1256),
.Y(n_1437)
);

BUFx10_ASAP7_75t_L g1438 ( 
.A(n_1339),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1300),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1335),
.B(n_1341),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1304),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1330),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1300),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1333),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1270),
.A2(n_1275),
.B1(n_1280),
.B2(n_1332),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1371),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1274),
.B(n_1340),
.Y(n_1447)
);

OAI21xp33_ASAP7_75t_L g1448 ( 
.A1(n_1276),
.A2(n_1256),
.B(n_1290),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1300),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1371),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1305),
.A2(n_1381),
.B(n_1376),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1326),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1374),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_SL g1454 ( 
.A1(n_1352),
.A2(n_1278),
.B1(n_1290),
.B2(n_1252),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1374),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1253),
.A2(n_1255),
.B1(n_1296),
.B2(n_1248),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1384),
.Y(n_1457)
);

BUFx2_ASAP7_75t_R g1458 ( 
.A(n_1324),
.Y(n_1458)
);

CKINVDCx14_ASAP7_75t_R g1459 ( 
.A(n_1384),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1340),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1384),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1253),
.A2(n_1255),
.B1(n_1292),
.B2(n_1303),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1281),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1308),
.B(n_1237),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1295),
.Y(n_1465)
);

BUFx5_ASAP7_75t_L g1466 ( 
.A(n_1260),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1338),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1295),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1337),
.A2(n_1336),
.B1(n_1313),
.B2(n_1316),
.Y(n_1469)
);

CKINVDCx8_ASAP7_75t_R g1470 ( 
.A(n_1370),
.Y(n_1470)
);

CKINVDCx8_ASAP7_75t_R g1471 ( 
.A(n_1266),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1325),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1336),
.Y(n_1473)
);

BUFx2_ASAP7_75t_SL g1474 ( 
.A(n_1329),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1353),
.A2(n_1233),
.B1(n_1262),
.B2(n_1258),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1353),
.Y(n_1476)
);

CKINVDCx11_ASAP7_75t_R g1477 ( 
.A(n_1298),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1334),
.Y(n_1478)
);

CKINVDCx11_ASAP7_75t_R g1479 ( 
.A(n_1334),
.Y(n_1479)
);

AOI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1343),
.A2(n_1368),
.B(n_1345),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1348),
.A2(n_1364),
.B1(n_1375),
.B2(n_1246),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1346),
.B(n_1369),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1235),
.A2(n_1234),
.B1(n_1249),
.B2(n_1329),
.Y(n_1483)
);

CKINVDCx14_ASAP7_75t_R g1484 ( 
.A(n_1246),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1244),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1310),
.A2(n_1249),
.B1(n_1311),
.B2(n_1317),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1242),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1231),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1244),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1244),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1385),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1331),
.A2(n_1294),
.B1(n_1230),
.B2(n_1346),
.Y(n_1492)
);

BUFx8_ASAP7_75t_L g1493 ( 
.A(n_1261),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1365),
.A2(n_1377),
.B1(n_1229),
.B2(n_1356),
.Y(n_1494)
);

BUFx8_ASAP7_75t_L g1495 ( 
.A(n_1346),
.Y(n_1495)
);

CKINVDCx11_ASAP7_75t_R g1496 ( 
.A(n_1356),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1356),
.B(n_1369),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1369),
.A2(n_1285),
.B1(n_1379),
.B2(n_1347),
.Y(n_1498)
);

BUFx2_ASAP7_75t_SL g1499 ( 
.A(n_1241),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1285),
.A2(n_1379),
.B1(n_1347),
.B2(n_1351),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1259),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1232),
.Y(n_1502)
);

INVx6_ASAP7_75t_L g1503 ( 
.A(n_1241),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1285),
.A2(n_1379),
.B1(n_1347),
.B2(n_1351),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1342),
.B(n_1347),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1280),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1241),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1285),
.A2(n_1379),
.B1(n_1347),
.B2(n_1351),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1367),
.Y(n_1509)
);

INVx6_ASAP7_75t_L g1510 ( 
.A(n_1241),
.Y(n_1510)
);

OAI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1379),
.A2(n_1347),
.B1(n_1351),
.B2(n_1342),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1232),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1379),
.A2(n_590),
.B1(n_1347),
.B2(n_1342),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1259),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1259),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1232),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1299),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1232),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1241),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1232),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1379),
.A2(n_1366),
.B1(n_1372),
.B2(n_1350),
.Y(n_1521)
);

BUFx4_ASAP7_75t_R g1522 ( 
.A(n_1380),
.Y(n_1522)
);

OAI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1379),
.A2(n_1347),
.B1(n_1351),
.B2(n_1342),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1379),
.A2(n_1347),
.B1(n_1351),
.B2(n_1342),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1241),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1379),
.A2(n_751),
.B1(n_761),
.B2(n_754),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1285),
.A2(n_1379),
.B1(n_1347),
.B2(n_1351),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1241),
.Y(n_1528)
);

INVx2_ASAP7_75t_R g1529 ( 
.A(n_1241),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1241),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_SL g1531 ( 
.A1(n_1379),
.A2(n_590),
.B1(n_1347),
.B2(n_1342),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1379),
.A2(n_751),
.B1(n_761),
.B2(n_754),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1259),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1379),
.A2(n_1285),
.B1(n_990),
.B2(n_1194),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1232),
.Y(n_1535)
);

BUFx12f_ASAP7_75t_L g1536 ( 
.A(n_1259),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1490),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1514),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1491),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1509),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1392),
.B(n_1500),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1509),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1399),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1489),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1482),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1534),
.A2(n_1532),
.B1(n_1526),
.B2(n_1414),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1480),
.B(n_1474),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1401),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1523),
.Y(n_1549)
);

OR2x6_ASAP7_75t_L g1550 ( 
.A(n_1481),
.B(n_1451),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1395),
.A2(n_1521),
.B(n_1396),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1497),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1399),
.B(n_1427),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1463),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1410),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1475),
.A2(n_1494),
.B(n_1483),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1398),
.A2(n_1513),
.B1(n_1531),
.B2(n_1400),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1485),
.Y(n_1558)
);

AOI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1396),
.A2(n_1419),
.B1(n_1511),
.B2(n_1523),
.C(n_1524),
.Y(n_1559)
);

AO21x2_ASAP7_75t_L g1560 ( 
.A1(n_1437),
.A2(n_1419),
.B(n_1472),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1495),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1389),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1495),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1452),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1431),
.Y(n_1565)
);

OAI221xp5_ASAP7_75t_L g1566 ( 
.A1(n_1392),
.A2(n_1504),
.B1(n_1500),
.B2(n_1508),
.C(n_1527),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1433),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1467),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1397),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1411),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1483),
.A2(n_1435),
.B(n_1448),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1397),
.Y(n_1572)
);

AO21x2_ASAP7_75t_L g1573 ( 
.A1(n_1437),
.A2(n_1492),
.B(n_1487),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1502),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1512),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1516),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1518),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1520),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1535),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1469),
.A2(n_1487),
.B(n_1456),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1464),
.Y(n_1581)
);

AO32x1_ASAP7_75t_L g1582 ( 
.A1(n_1426),
.A2(n_1444),
.A3(n_1442),
.B1(n_1432),
.B2(n_1447),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1498),
.B(n_1432),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1456),
.A2(n_1462),
.B(n_1435),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1466),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1434),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1462),
.A2(n_1445),
.B(n_1450),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1407),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1522),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1498),
.B(n_1426),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1446),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1454),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1488),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1454),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1496),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1513),
.A2(n_1531),
.B1(n_1504),
.B2(n_1527),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1436),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1406),
.B(n_1508),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1486),
.Y(n_1599)
);

NAND2x1p5_ASAP7_75t_L g1600 ( 
.A(n_1440),
.B(n_1403),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1486),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1493),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1524),
.B(n_1391),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1493),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1412),
.A2(n_1424),
.B(n_1414),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_SL g1606 ( 
.A(n_1515),
.B(n_1536),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1413),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1478),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1506),
.B(n_1473),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1479),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1422),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1422),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1519),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1484),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1506),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1412),
.A2(n_1505),
.B(n_1530),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1476),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1429),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1390),
.B(n_1402),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1476),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1476),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1477),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1438),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1428),
.A2(n_1409),
.B(n_1465),
.Y(n_1624)
);

CKINVDCx16_ASAP7_75t_R g1625 ( 
.A(n_1405),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1519),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1438),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1468),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1529),
.Y(n_1629)
);

BUFx4f_ASAP7_75t_SL g1630 ( 
.A(n_1501),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1529),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1519),
.Y(n_1632)
);

AOI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1458),
.A2(n_1499),
.B(n_1503),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_SL g1634 ( 
.A(n_1525),
.B(n_1530),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1525),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1525),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1528),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1393),
.A2(n_1425),
.B1(n_1517),
.B2(n_1441),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1404),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1460),
.B(n_1421),
.Y(n_1640)
);

INVx4_ASAP7_75t_L g1641 ( 
.A(n_1528),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1507),
.B(n_1530),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1530),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1609),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1586),
.B(n_1394),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1561),
.B(n_1449),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_R g1647 ( 
.A(n_1589),
.B(n_1420),
.Y(n_1647)
);

AO32x2_ASAP7_75t_L g1648 ( 
.A1(n_1546),
.A2(n_1417),
.A3(n_1507),
.B1(n_1416),
.B2(n_1459),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1553),
.B(n_1394),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1553),
.B(n_1443),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1551),
.A2(n_1416),
.B(n_1417),
.Y(n_1651)
);

O2A1O1Ixp33_ASAP7_75t_SL g1652 ( 
.A1(n_1559),
.A2(n_1533),
.B(n_1471),
.C(n_1408),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1550),
.B(n_1510),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1550),
.B(n_1510),
.Y(n_1654)
);

A2O1A1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1549),
.A2(n_1461),
.B(n_1453),
.C(n_1457),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1603),
.B(n_1421),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1596),
.A2(n_1510),
.B1(n_1503),
.B2(n_1470),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1609),
.B(n_1455),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1609),
.B(n_1421),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1597),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1556),
.A2(n_1503),
.B(n_1415),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1543),
.B(n_1421),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1596),
.A2(n_1423),
.B1(n_1415),
.B2(n_1430),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1593),
.B(n_1423),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1619),
.B(n_1439),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1598),
.B(n_1415),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_SL g1667 ( 
.A(n_1566),
.B(n_1607),
.Y(n_1667)
);

INVx6_ASAP7_75t_L g1668 ( 
.A(n_1607),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1550),
.B(n_1418),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1574),
.Y(n_1670)
);

OAI211xp5_ASAP7_75t_L g1671 ( 
.A1(n_1557),
.A2(n_1541),
.B(n_1616),
.C(n_1605),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1564),
.B(n_1540),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_R g1673 ( 
.A(n_1538),
.B(n_1625),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1598),
.A2(n_1622),
.B1(n_1595),
.B2(n_1605),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1597),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1590),
.A2(n_1605),
.B1(n_1612),
.B2(n_1611),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1640),
.B(n_1595),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1611),
.A2(n_1612),
.B(n_1567),
.Y(n_1678)
);

BUFx4f_ASAP7_75t_SL g1679 ( 
.A(n_1588),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1630),
.Y(n_1680)
);

A2O1A1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1590),
.A2(n_1583),
.B(n_1584),
.C(n_1608),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1610),
.B(n_1600),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1625),
.B(n_1618),
.Y(n_1683)
);

AO32x2_ASAP7_75t_L g1684 ( 
.A1(n_1591),
.A2(n_1582),
.A3(n_1560),
.B1(n_1626),
.B2(n_1641),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1610),
.B(n_1600),
.Y(n_1685)
);

AO221x1_ASAP7_75t_L g1686 ( 
.A1(n_1592),
.A2(n_1594),
.B1(n_1561),
.B2(n_1563),
.C(n_1544),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1540),
.B(n_1542),
.Y(n_1687)
);

AND2x2_ASAP7_75t_SL g1688 ( 
.A(n_1605),
.B(n_1583),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1548),
.B(n_1555),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1550),
.A2(n_1624),
.B1(n_1622),
.B2(n_1608),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_SL g1691 ( 
.A1(n_1602),
.A2(n_1604),
.B(n_1563),
.C(n_1614),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1581),
.A2(n_1608),
.B1(n_1592),
.B2(n_1594),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1560),
.A2(n_1562),
.B1(n_1581),
.B2(n_1542),
.C(n_1601),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1547),
.A2(n_1582),
.B(n_1571),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1547),
.A2(n_1582),
.B(n_1571),
.Y(n_1695)
);

OA21x2_ASAP7_75t_L g1696 ( 
.A1(n_1584),
.A2(n_1556),
.B(n_1587),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1565),
.B(n_1576),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1599),
.A2(n_1601),
.B(n_1580),
.C(n_1606),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1575),
.B(n_1577),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1560),
.A2(n_1604),
.B1(n_1602),
.B2(n_1571),
.Y(n_1700)
);

NAND2xp33_ASAP7_75t_L g1701 ( 
.A(n_1638),
.B(n_1623),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1588),
.B(n_1570),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1599),
.A2(n_1544),
.B1(n_1579),
.B2(n_1578),
.C(n_1572),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1591),
.B(n_1623),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1578),
.B(n_1579),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1547),
.A2(n_1582),
.B(n_1571),
.Y(n_1706)
);

OR2x6_ASAP7_75t_L g1707 ( 
.A(n_1547),
.B(n_1580),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1582),
.A2(n_1573),
.B(n_1634),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1568),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1545),
.B(n_1552),
.Y(n_1710)
);

AND2x2_ASAP7_75t_SL g1711 ( 
.A(n_1591),
.B(n_1642),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1573),
.A2(n_1634),
.B(n_1585),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1569),
.A2(n_1572),
.B1(n_1545),
.B2(n_1552),
.C(n_1573),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1709),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1688),
.B(n_1569),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1677),
.B(n_1587),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1670),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1672),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1704),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1667),
.B(n_1627),
.C(n_1615),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1676),
.B(n_1554),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1669),
.A2(n_1570),
.B1(n_1621),
.B2(n_1620),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1704),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1669),
.A2(n_1621),
.B1(n_1617),
.B2(n_1620),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1644),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1664),
.B(n_1627),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1705),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1662),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1676),
.B(n_1554),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1699),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1682),
.B(n_1685),
.Y(n_1731)
);

NAND2x1_ASAP7_75t_L g1732 ( 
.A(n_1669),
.B(n_1629),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1671),
.A2(n_1633),
.B1(n_1620),
.B2(n_1617),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1657),
.A2(n_1617),
.B1(n_1613),
.B2(n_1631),
.Y(n_1734)
);

INVxp67_ASAP7_75t_SL g1735 ( 
.A(n_1687),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1666),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1689),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1697),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1710),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1707),
.B(n_1661),
.Y(n_1740)
);

INVx5_ASAP7_75t_L g1741 ( 
.A(n_1707),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1700),
.B(n_1558),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1700),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1703),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1684),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1681),
.B(n_1537),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1684),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1684),
.B(n_1629),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1686),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1678),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1653),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1657),
.A2(n_1663),
.B1(n_1678),
.B2(n_1674),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1692),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1692),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1717),
.Y(n_1755)
);

OAI33xp33_ASAP7_75t_L g1756 ( 
.A1(n_1744),
.A2(n_1656),
.A3(n_1663),
.B1(n_1645),
.B2(n_1628),
.B3(n_1637),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1750),
.B(n_1735),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1748),
.B(n_1696),
.Y(n_1758)
);

OAI321xp33_ASAP7_75t_L g1759 ( 
.A1(n_1733),
.A2(n_1690),
.A3(n_1698),
.B1(n_1693),
.B2(n_1651),
.C(n_1633),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1715),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1744),
.A2(n_1652),
.B1(n_1713),
.B2(n_1701),
.C(n_1695),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1745),
.B(n_1696),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1745),
.B(n_1694),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1748),
.B(n_1706),
.Y(n_1764)
);

AO21x2_ASAP7_75t_L g1765 ( 
.A1(n_1743),
.A2(n_1708),
.B(n_1712),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1716),
.B(n_1698),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1740),
.Y(n_1767)
);

AO21x2_ASAP7_75t_L g1768 ( 
.A1(n_1743),
.A2(n_1747),
.B(n_1729),
.Y(n_1768)
);

OAI33xp33_ASAP7_75t_L g1769 ( 
.A1(n_1749),
.A2(n_1628),
.A3(n_1632),
.B1(n_1636),
.B2(n_1643),
.B3(n_1635),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1714),
.Y(n_1770)
);

OAI31xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1752),
.A2(n_1651),
.A3(n_1683),
.B(n_1648),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1725),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1725),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1714),
.Y(n_1774)
);

INVxp67_ASAP7_75t_SL g1775 ( 
.A(n_1715),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1733),
.A2(n_1654),
.B(n_1711),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1737),
.B(n_1648),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1737),
.B(n_1648),
.Y(n_1778)
);

NAND4xp25_ASAP7_75t_L g1779 ( 
.A(n_1752),
.B(n_1690),
.C(n_1655),
.D(n_1702),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1741),
.B(n_1740),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1732),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1740),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1720),
.A2(n_1668),
.B1(n_1649),
.B2(n_1665),
.Y(n_1783)
);

AOI33xp33_ASAP7_75t_L g1784 ( 
.A1(n_1749),
.A2(n_1691),
.A3(n_1650),
.B1(n_1646),
.B2(n_1658),
.B3(n_1659),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1735),
.B(n_1539),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1721),
.B(n_1729),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1753),
.A2(n_1754),
.B1(n_1721),
.B2(n_1720),
.C(n_1746),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1786),
.B(n_1739),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1786),
.B(n_1736),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1758),
.B(n_1741),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1772),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1758),
.B(n_1741),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1755),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1758),
.B(n_1741),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1786),
.B(n_1736),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1780),
.B(n_1740),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1763),
.B(n_1760),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1772),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1770),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1764),
.B(n_1742),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1763),
.B(n_1760),
.Y(n_1801)
);

NOR3xp33_ASAP7_75t_SL g1802 ( 
.A(n_1759),
.B(n_1680),
.C(n_1726),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1764),
.B(n_1742),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1764),
.B(n_1731),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1767),
.B(n_1731),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1767),
.B(n_1728),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1770),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1763),
.B(n_1738),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1775),
.B(n_1738),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1775),
.B(n_1739),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1757),
.B(n_1727),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1767),
.B(n_1746),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1757),
.B(n_1727),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1767),
.B(n_1730),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1770),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1780),
.B(n_1767),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1773),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1718),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1768),
.B(n_1753),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1781),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1782),
.B(n_1730),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1782),
.B(n_1719),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1782),
.B(n_1719),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1782),
.B(n_1723),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1787),
.B(n_1768),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1768),
.B(n_1754),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1774),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1773),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1768),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1782),
.B(n_1723),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1797),
.B(n_1768),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1797),
.B(n_1801),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1820),
.B(n_1781),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1820),
.B(n_1781),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1800),
.B(n_1766),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1827),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1802),
.A2(n_1761),
.B1(n_1779),
.B2(n_1766),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1800),
.B(n_1766),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1791),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1827),
.Y(n_1840)
);

AOI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1825),
.A2(n_1771),
.B(n_1759),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1818),
.B(n_1784),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1800),
.B(n_1780),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1799),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1793),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1793),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1799),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1793),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_SL g1849 ( 
.A(n_1825),
.B(n_1761),
.C(n_1783),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1818),
.A2(n_1779),
.B1(n_1776),
.B2(n_1783),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1801),
.B(n_1762),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1789),
.B(n_1784),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1807),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1828),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1803),
.B(n_1780),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1814),
.Y(n_1856)
);

AOI21xp33_ASAP7_75t_L g1857 ( 
.A1(n_1820),
.A2(n_1771),
.B(n_1765),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1789),
.B(n_1777),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1798),
.B(n_1776),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1807),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1795),
.B(n_1777),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1795),
.B(n_1777),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1815),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1803),
.B(n_1780),
.Y(n_1864)
);

NAND3xp33_ASAP7_75t_L g1865 ( 
.A(n_1819),
.B(n_1734),
.C(n_1722),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1808),
.B(n_1762),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1796),
.B(n_1781),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1803),
.B(n_1778),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1815),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1798),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1788),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1808),
.B(n_1762),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1788),
.B(n_1785),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1810),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1832),
.B(n_1819),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1867),
.B(n_1796),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1856),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1835),
.B(n_1796),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1841),
.A2(n_1796),
.B1(n_1756),
.B2(n_1751),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1867),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1836),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1856),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1832),
.B(n_1826),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1835),
.B(n_1796),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1840),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1839),
.B(n_1826),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1843),
.Y(n_1887)
);

CKINVDCx20_ASAP7_75t_R g1888 ( 
.A(n_1837),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1838),
.B(n_1812),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1838),
.B(n_1843),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1844),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1842),
.B(n_1668),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1844),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1870),
.Y(n_1894)
);

O2A1O1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1849),
.A2(n_1829),
.B(n_1817),
.C(n_1756),
.Y(n_1895)
);

OR2x6_ASAP7_75t_L g1896 ( 
.A(n_1859),
.B(n_1732),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1850),
.B(n_1804),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1855),
.B(n_1812),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1867),
.B(n_1816),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1855),
.B(n_1812),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1864),
.B(n_1816),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1873),
.B(n_1811),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1847),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1864),
.B(n_1816),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1859),
.A2(n_1734),
.B1(n_1765),
.B2(n_1817),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1852),
.B(n_1804),
.Y(n_1906)
);

NAND4xp25_ASAP7_75t_L g1907 ( 
.A(n_1857),
.B(n_1829),
.C(n_1660),
.D(n_1675),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1854),
.B(n_1804),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1833),
.B(n_1816),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1833),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1874),
.Y(n_1911)
);

AOI31xp33_ASAP7_75t_L g1912 ( 
.A1(n_1894),
.A2(n_1865),
.A3(n_1834),
.B(n_1833),
.Y(n_1912)
);

AOI21xp33_ASAP7_75t_L g1913 ( 
.A1(n_1895),
.A2(n_1871),
.B(n_1834),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1891),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1894),
.B(n_1873),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1891),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1893),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1888),
.B(n_1868),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1890),
.B(n_1834),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1880),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1910),
.B(n_1868),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1880),
.Y(n_1922)
);

OAI21xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1905),
.A2(n_1792),
.B(n_1790),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1890),
.B(n_1816),
.Y(n_1924)
);

NOR2xp67_ASAP7_75t_L g1925 ( 
.A(n_1880),
.B(n_1851),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1880),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1905),
.B(n_1907),
.C(n_1879),
.Y(n_1927)
);

AOI221x1_ASAP7_75t_L g1928 ( 
.A1(n_1907),
.A2(n_1869),
.B1(n_1860),
.B2(n_1863),
.C(n_1853),
.Y(n_1928)
);

NAND2x1_ASAP7_75t_SL g1929 ( 
.A(n_1876),
.B(n_1899),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1899),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1892),
.A2(n_1765),
.B1(n_1794),
.B2(n_1790),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1893),
.Y(n_1932)
);

OAI21xp33_ASAP7_75t_SL g1933 ( 
.A1(n_1897),
.A2(n_1831),
.B(n_1851),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1911),
.B(n_1811),
.Y(n_1934)
);

AOI221x1_ASAP7_75t_L g1935 ( 
.A1(n_1881),
.A2(n_1810),
.B1(n_1861),
.B2(n_1862),
.C(n_1858),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1906),
.B(n_1813),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1881),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1914),
.Y(n_1938)
);

AOI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1927),
.A2(n_1876),
.B1(n_1908),
.B2(n_1896),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1916),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1918),
.B(n_1926),
.Y(n_1941)
);

OAI21xp33_ASAP7_75t_L g1942 ( 
.A1(n_1912),
.A2(n_1887),
.B(n_1884),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1917),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1919),
.B(n_1909),
.Y(n_1944)
);

OAI21xp33_ASAP7_75t_L g1945 ( 
.A1(n_1923),
.A2(n_1921),
.B(n_1933),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1930),
.B(n_1887),
.Y(n_1946)
);

OAI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1928),
.A2(n_1896),
.B1(n_1886),
.B2(n_1831),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1925),
.B(n_1876),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1932),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1928),
.B(n_1885),
.C(n_1896),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1937),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1920),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1930),
.B(n_1889),
.Y(n_1953)
);

OAI322xp33_ASAP7_75t_L g1954 ( 
.A1(n_1915),
.A2(n_1886),
.A3(n_1883),
.B1(n_1875),
.B2(n_1885),
.C1(n_1903),
.C2(n_1902),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1919),
.B(n_1909),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1915),
.B(n_1920),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1922),
.B(n_1934),
.Y(n_1957)
);

NOR4xp25_ASAP7_75t_L g1958 ( 
.A(n_1947),
.B(n_1913),
.C(n_1922),
.D(n_1903),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1952),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1941),
.B(n_1936),
.Y(n_1960)
);

A2O1A1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1945),
.A2(n_1950),
.B(n_1939),
.C(n_1942),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1956),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1946),
.Y(n_1963)
);

HAxp5_ASAP7_75t_SL g1964 ( 
.A(n_1947),
.B(n_1931),
.CON(n_1964),
.SN(n_1964)
);

AOI21xp33_ASAP7_75t_L g1965 ( 
.A1(n_1948),
.A2(n_1896),
.B(n_1882),
.Y(n_1965)
);

AOI211xp5_ASAP7_75t_SL g1966 ( 
.A1(n_1954),
.A2(n_1929),
.B(n_1876),
.C(n_1924),
.Y(n_1966)
);

OAI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1948),
.A2(n_1929),
.B1(n_1896),
.B2(n_1902),
.C(n_1875),
.Y(n_1967)
);

OAI221xp5_ASAP7_75t_L g1968 ( 
.A1(n_1953),
.A2(n_1883),
.B1(n_1877),
.B2(n_1882),
.C(n_1878),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1957),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1961),
.B(n_1955),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1969),
.B(n_1960),
.Y(n_1971)
);

NOR3xp33_ASAP7_75t_L g1972 ( 
.A(n_1961),
.B(n_1951),
.C(n_1940),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_L g1973 ( 
.A(n_1964),
.B(n_1935),
.C(n_1938),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1958),
.A2(n_1935),
.B(n_1955),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1966),
.B(n_1944),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1963),
.B(n_1962),
.Y(n_1976)
);

NOR2x1_ASAP7_75t_L g1977 ( 
.A(n_1959),
.B(n_1943),
.Y(n_1977)
);

OAI21xp33_ASAP7_75t_SL g1978 ( 
.A1(n_1964),
.A2(n_1924),
.B(n_1884),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1968),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1965),
.B(n_1878),
.Y(n_1980)
);

NAND5xp2_ASAP7_75t_L g1981 ( 
.A(n_1967),
.B(n_1949),
.C(n_1889),
.D(n_1901),
.E(n_1904),
.Y(n_1981)
);

AOI211xp5_ASAP7_75t_L g1982 ( 
.A1(n_1973),
.A2(n_1978),
.B(n_1974),
.C(n_1972),
.Y(n_1982)
);

AOI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1970),
.A2(n_1899),
.B(n_1673),
.C(n_1877),
.Y(n_1983)
);

O2A1O1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1979),
.A2(n_1866),
.B(n_1872),
.C(n_1900),
.Y(n_1984)
);

AND4x1_ASAP7_75t_L g1985 ( 
.A(n_1971),
.B(n_1976),
.C(n_1975),
.D(n_1977),
.Y(n_1985)
);

O2A1O1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1981),
.A2(n_1866),
.B(n_1872),
.C(n_1900),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_R g1987 ( 
.A(n_1980),
.B(n_1679),
.Y(n_1987)
);

OAI211xp5_ASAP7_75t_L g1988 ( 
.A1(n_1978),
.A2(n_1647),
.B(n_1901),
.C(n_1904),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1984),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1982),
.A2(n_1899),
.B1(n_1898),
.B2(n_1848),
.C(n_1846),
.Y(n_1990)
);

AOI321xp33_ASAP7_75t_L g1991 ( 
.A1(n_1988),
.A2(n_1898),
.A3(n_1794),
.B1(n_1792),
.B2(n_1790),
.C(n_1724),
.Y(n_1991)
);

AOI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1983),
.A2(n_1848),
.B1(n_1846),
.B2(n_1845),
.C(n_1792),
.Y(n_1992)
);

OAI211xp5_ASAP7_75t_L g1993 ( 
.A1(n_1987),
.A2(n_1794),
.B(n_1845),
.C(n_1809),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1985),
.Y(n_1994)
);

AOI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1986),
.A2(n_1765),
.B1(n_1769),
.B2(n_1823),
.C(n_1822),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1994),
.B(n_1805),
.Y(n_1996)
);

NAND4xp75_ASAP7_75t_L g1997 ( 
.A(n_1989),
.B(n_1830),
.C(n_1822),
.D(n_1824),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1990),
.B(n_1822),
.Y(n_1998)
);

AOI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1993),
.A2(n_1830),
.B1(n_1824),
.B2(n_1823),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1991),
.Y(n_2000)
);

XNOR2xp5_ASAP7_75t_L g2001 ( 
.A(n_1992),
.B(n_1646),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_2000),
.B(n_1995),
.Y(n_2002)
);

XNOR2xp5_ASAP7_75t_L g2003 ( 
.A(n_1996),
.B(n_1642),
.Y(n_2003)
);

A2O1A1Ixp33_ASAP7_75t_L g2004 ( 
.A1(n_1998),
.A2(n_1830),
.B(n_1824),
.C(n_1823),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_2003),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_2005),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_2006),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_2006),
.Y(n_2008)
);

OR2x6_ASAP7_75t_L g2009 ( 
.A(n_2007),
.B(n_2002),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_2008),
.B(n_2001),
.Y(n_2010)
);

OAI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_2010),
.A2(n_1997),
.B(n_2004),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_2009),
.B(n_1999),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_2012),
.A2(n_1813),
.B(n_1809),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_2013),
.A2(n_2011),
.B1(n_1806),
.B2(n_1814),
.Y(n_2014)
);

OAI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_2014),
.A2(n_1613),
.B1(n_1626),
.B2(n_1641),
.Y(n_2015)
);

OAI221xp5_ASAP7_75t_R g2016 ( 
.A1(n_2015),
.A2(n_1769),
.B1(n_1806),
.B2(n_1765),
.C(n_1821),
.Y(n_2016)
);

AOI211xp5_ASAP7_75t_L g2017 ( 
.A1(n_2016),
.A2(n_1613),
.B(n_1642),
.C(n_1639),
.Y(n_2017)
);


endmodule