module fake_jpeg_20063_n_290 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_15),
.B1(n_21),
.B2(n_23),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_40),
.B1(n_32),
.B2(n_15),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_15),
.B1(n_23),
.B2(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_50),
.B1(n_65),
.B2(n_54),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_49),
.Y(n_80)
);

NAND2x1_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_32),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_38),
.B(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_33),
.B(n_27),
.C(n_32),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_20),
.B1(n_12),
.B2(n_23),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_61),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_21),
.B1(n_16),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_37),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_67),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_48),
.B(n_50),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_45),
.B1(n_37),
.B2(n_44),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_45),
.B1(n_37),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_45),
.B1(n_35),
.B2(n_43),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_35),
.B1(n_43),
.B2(n_24),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_56),
.B1(n_59),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_83),
.B1(n_58),
.B2(n_12),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_25),
.C(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_25),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_43),
.B1(n_26),
.B2(n_20),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_91),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_30),
.C(n_28),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_61),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_98),
.B(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_26),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_56),
.B1(n_49),
.B2(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_68),
.B1(n_84),
.B2(n_63),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_58),
.B1(n_57),
.B2(n_12),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_25),
.C(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_100),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_30),
.B(n_25),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_79),
.B1(n_76),
.B2(n_73),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_42),
.B1(n_17),
.B2(n_24),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_42),
.B1(n_17),
.B2(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_18),
.B1(n_19),
.B2(n_42),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_84),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_25),
.Y(n_106)
);

AOI22x1_ASAP7_75t_R g110 ( 
.A1(n_106),
.A2(n_25),
.B1(n_30),
.B2(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_75),
.B1(n_71),
.B2(n_85),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_131),
.B1(n_87),
.B2(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_92),
.B1(n_109),
.B2(n_132),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_111),
.B(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_85),
.B1(n_68),
.B2(n_75),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_119),
.A2(n_18),
.B1(n_28),
.B2(n_29),
.Y(n_162)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_77),
.C(n_85),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_34),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_68),
.B1(n_71),
.B2(n_19),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_124),
.Y(n_134)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_98),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_87),
.B(n_98),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_104),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_100),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_31),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_103),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_63),
.B1(n_34),
.B2(n_31),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_132),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_133),
.A2(n_141),
.B(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_140),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_146),
.B1(n_116),
.B2(n_131),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_127),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_153),
.B1(n_162),
.B2(n_120),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_34),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_19),
.B(n_18),
.C(n_22),
.D(n_28),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_124),
.Y(n_176)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_31),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_22),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_19),
.B(n_18),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_29),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_29),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_111),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_118),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_121),
.C(n_125),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_174),
.C(n_183),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_135),
.B(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_167),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_114),
.B(n_113),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_188),
.B1(n_143),
.B2(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_115),
.C(n_123),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_189),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_123),
.B1(n_114),
.B2(n_130),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_114),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_160),
.B(n_136),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_184),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_28),
.B1(n_14),
.B2(n_22),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_22),
.C(n_14),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_138),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_22),
.C(n_14),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_142),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_194),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_179),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_206),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_177),
.B(n_142),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_203),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_157),
.B(n_158),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_134),
.B(n_168),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_207),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_147),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_175),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_178),
.B1(n_146),
.B2(n_182),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_154),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_211),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVxp33_ASAP7_75t_SL g213 ( 
.A(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_188),
.B1(n_149),
.B2(n_150),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_216),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_150),
.B1(n_166),
.B2(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_183),
.C(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_227),
.C(n_195),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_180),
.B1(n_185),
.B2(n_135),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_224),
.Y(n_242)
);

FAx1_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_176),
.CI(n_148),
.CON(n_223),
.SN(n_223)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_189),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_202),
.B1(n_3),
.B2(n_4),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_14),
.C(n_2),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_198),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_1),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_211),
.C(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_206),
.C(n_195),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_196),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_236),
.Y(n_249)
);

FAx1_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_210),
.CI(n_199),
.CON(n_236),
.SN(n_236)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_241),
.B1(n_223),
.B2(n_217),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_226),
.B1(n_4),
.B2(n_5),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_225),
.B(n_1),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_225),
.C(n_217),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_248),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_219),
.B(n_213),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_252),
.Y(n_263)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_231),
.B(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_223),
.B1(n_4),
.B2(n_5),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_264),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_260),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_244),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_236),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_265),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_3),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_6),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_249),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_273),
.B(n_266),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_6),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_7),
.C(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_10),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_7),
.B(n_8),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_276),
.A2(n_277),
.B(n_268),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_8),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_279),
.A2(n_267),
.B(n_11),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_280),
.C(n_269),
.Y(n_287)
);

OAI211xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_286),
.B(n_282),
.C(n_281),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_288),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_10),
.B(n_11),
.Y(n_290)
);


endmodule