module fake_jpeg_31669_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_32),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_38),
.B1(n_48),
.B2(n_47),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_51),
.B1(n_44),
.B2(n_50),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_68),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_7),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_3),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_38),
.B1(n_49),
.B2(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_40),
.B1(n_21),
.B2(n_5),
.Y(n_67)
);

NOR2x1_ASAP7_75t_R g68 ( 
.A(n_53),
.B(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_3),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_9),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_11),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_15),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_86),
.Y(n_100)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_28),
.B(n_29),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_24),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_90),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_89),
.B(n_92),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_88),
.B(n_100),
.C(n_94),
.D(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_99),
.C(n_88),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_102),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_105),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_108),
.A2(n_87),
.B(n_95),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_31),
.Y(n_111)
);


endmodule