module fake_jpeg_2695_n_439 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_439);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_439;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_15),
.B(n_14),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_32),
.B(n_37),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_51),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_53),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_80),
.Y(n_113)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_34),
.B(n_15),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_13),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_13),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_2),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_92),
.B(n_5),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_101),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_35),
.B1(n_43),
.B2(n_17),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_119),
.B1(n_127),
.B2(n_129),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_37),
.B1(n_25),
.B2(n_22),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_117),
.A2(n_118),
.B(n_125),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_25),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_20),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_18),
.B1(n_17),
.B2(n_32),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_132),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_71),
.A2(n_26),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_62),
.B(n_2),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_113),
.B1(n_119),
.B2(n_88),
.Y(n_169)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_48),
.Y(n_136)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_46),
.Y(n_139)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_60),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_55),
.B1(n_85),
.B2(n_74),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_143),
.B(n_164),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_67),
.B1(n_76),
.B2(n_61),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_144),
.A2(n_146),
.B1(n_162),
.B2(n_169),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_51),
.B1(n_79),
.B2(n_66),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_81),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_147),
.B(n_165),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_49),
.B1(n_57),
.B2(n_56),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_149),
.B(n_195),
.Y(n_216)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_152),
.Y(n_232)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_105),
.A2(n_45),
.B1(n_54),
.B2(n_53),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_155),
.A2(n_156),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_100),
.B1(n_127),
.B2(n_135),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_60),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_47),
.B1(n_80),
.B2(n_50),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_101),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_99),
.B(n_4),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_87),
.B(n_50),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_102),
.B(n_4),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_114),
.Y(n_173)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_106),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_175),
.A2(n_138),
.B1(n_137),
.B2(n_122),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_10),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_108),
.B(n_5),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_177),
.B(n_182),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_186),
.Y(n_208)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_130),
.B(n_6),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_189),
.C(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_95),
.B(n_6),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_120),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_89),
.B(n_8),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_95),
.B(n_8),
.Y(n_189)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_97),
.B(n_9),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_114),
.A2(n_9),
.B(n_10),
.C(n_98),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_149),
.B1(n_147),
.B2(n_146),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_198),
.A2(n_207),
.B1(n_210),
.B2(n_215),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_199),
.B(n_190),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_154),
.A2(n_116),
.B1(n_137),
.B2(n_121),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_98),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_211),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_158),
.A2(n_116),
.B1(n_122),
.B2(n_114),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_217),
.A2(n_225),
.B1(n_237),
.B2(n_205),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_174),
.B(n_10),
.CI(n_183),
.CON(n_221),
.SN(n_221)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_221),
.B(n_223),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_223),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_189),
.B1(n_182),
.B2(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_180),
.A2(n_165),
.B1(n_176),
.B2(n_179),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_230),
.A2(n_184),
.B1(n_185),
.B2(n_160),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_180),
.C(n_145),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_167),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_157),
.B(n_145),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_235),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_163),
.A2(n_187),
.B(n_153),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_236),
.A2(n_240),
.B(n_219),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_172),
.A2(n_151),
.B1(n_148),
.B2(n_161),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_148),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_163),
.A2(n_192),
.B(n_191),
.C(n_187),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_240),
.A2(n_220),
.B(n_204),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_242),
.B(n_249),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_152),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_253),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_244),
.B(n_245),
.Y(n_308)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_181),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_201),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_150),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_150),
.B1(n_181),
.B2(n_216),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_262),
.B1(n_263),
.B2(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_237),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_267),
.Y(n_292)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_216),
.A2(n_224),
.B1(n_222),
.B2(n_213),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_224),
.B1(n_215),
.B2(n_198),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_196),
.B(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_265),
.B(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_230),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_259),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_200),
.Y(n_269)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_272),
.A2(n_277),
.B(n_219),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_223),
.A2(n_226),
.B1(n_220),
.B2(n_210),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_282),
.B1(n_214),
.B2(n_233),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_279),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_281),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_203),
.B(n_202),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_234),
.A2(n_233),
.B1(n_214),
.B2(n_221),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_273),
.B(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_287),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_262),
.B(n_221),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_293),
.C(n_315),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_290),
.A2(n_295),
.B1(n_309),
.B2(n_312),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_232),
.C(n_241),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_294),
.A2(n_300),
.B(n_301),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_202),
.B1(n_232),
.B2(n_231),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_253),
.B1(n_243),
.B2(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_269),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_272),
.B(n_273),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_257),
.A2(n_276),
.B(n_275),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_302),
.A2(n_279),
.B(n_297),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_271),
.B(n_258),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_305),
.A2(n_307),
.B(n_311),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_256),
.A2(n_282),
.B(n_268),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_274),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_246),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_280),
.A2(n_260),
.B1(n_250),
.B2(n_251),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_246),
.B(n_254),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_286),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_332),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_264),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_323),
.B(n_328),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_324),
.Y(n_359)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_325),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_SL g326 ( 
.A(n_302),
.B(n_305),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_326),
.B(n_316),
.Y(n_369)
);

BUFx12_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_327),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_247),
.C(n_261),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_289),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_329),
.B(n_335),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_247),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_330),
.B(n_331),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_255),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_286),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_285),
.A2(n_274),
.B1(n_279),
.B2(n_248),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_337),
.B1(n_296),
.B2(n_301),
.Y(n_347)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_334),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_336),
.A2(n_339),
.B1(n_342),
.B2(n_343),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_285),
.A2(n_290),
.B1(n_297),
.B2(n_301),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_340),
.A2(n_341),
.B(n_344),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_292),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_287),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_347),
.A2(n_368),
.B1(n_322),
.B2(n_332),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_338),
.A2(n_294),
.B(n_291),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_354),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_334),
.A2(n_295),
.B1(n_291),
.B2(n_312),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_351),
.A2(n_365),
.B1(n_319),
.B2(n_313),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_308),
.C(n_293),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_345),
.C(n_344),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_318),
.A2(n_309),
.B1(n_284),
.B2(n_310),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_321),
.B(n_308),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_357),
.B(n_369),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_318),
.A2(n_335),
.B(n_338),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_363),
.C(n_306),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_340),
.A2(n_298),
.B(n_306),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_337),
.A2(n_287),
.B1(n_284),
.B2(n_317),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_288),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_327),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_341),
.A2(n_315),
.B1(n_313),
.B2(n_316),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_374),
.Y(n_393)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_368),
.Y(n_371)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_352),
.Y(n_372)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_SL g373 ( 
.A(n_366),
.B(n_325),
.C(n_343),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_373),
.B(n_376),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_345),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_352),
.Y(n_376)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_333),
.C(n_320),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_382),
.C(n_385),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_379),
.A2(n_383),
.B1(n_387),
.B2(n_388),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_380),
.A2(n_350),
.B(n_351),
.Y(n_398)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_384),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_367),
.A2(n_339),
.B1(n_324),
.B2(n_327),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_327),
.C(n_346),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_363),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_386),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_355),
.Y(n_387)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_355),
.C(n_362),
.Y(n_388)
);

A2O1A1O1Ixp25_ASAP7_75t_L g394 ( 
.A1(n_385),
.A2(n_346),
.B(n_360),
.C(n_362),
.D(n_347),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_394),
.A2(n_389),
.B(n_382),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_364),
.C(n_349),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_400),
.C(n_402),
.Y(n_412)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_354),
.C(n_365),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_356),
.C(n_358),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_356),
.Y(n_403)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_403),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_358),
.B1(n_359),
.B2(n_389),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_389),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_416),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_359),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_410),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_409),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_402),
.B(n_375),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_393),
.B(n_375),
.Y(n_413)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_413),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_399),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_415),
.B(n_397),
.C(n_391),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_396),
.Y(n_416)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_417),
.Y(n_426)
);

BUFx4f_ASAP7_75t_SL g421 ( 
.A(n_414),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_421),
.B(n_392),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_396),
.C(n_400),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_423),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_401),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_420),
.C(n_418),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_427),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_411),
.C(n_408),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_392),
.B(n_403),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_428),
.A2(n_424),
.B(n_394),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_431),
.B(n_421),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_434),
.A2(n_432),
.B(n_398),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_433),
.C(n_429),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_436),
.A2(n_426),
.B(n_405),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_405),
.B(n_406),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_421),
.Y(n_439)
);


endmodule