module fake_jpeg_24796_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_15),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_21),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_15),
.B1(n_25),
.B2(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_59),
.B1(n_15),
.B2(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_15),
.B1(n_25),
.B2(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_95)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_76),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_71),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_75),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_80),
.Y(n_101)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_86),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_45),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_96),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_74),
.B(n_77),
.C(n_42),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_102),
.B(n_27),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_28),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_99),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_26),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_52),
.B1(n_57),
.B2(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_52),
.B1(n_36),
.B2(n_37),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_85),
.B1(n_71),
.B2(n_82),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_33),
.B(n_36),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_79),
.C(n_37),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_46),
.B1(n_27),
.B2(n_51),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_80),
.B(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_45),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_67),
.Y(n_123)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_129),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_130),
.B(n_131),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_116),
.B(n_120),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_121),
.B(n_123),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_126),
.B(n_96),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_107),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_11),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_132),
.C(n_100),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_51),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_88),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_107),
.B(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_63),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_116),
.B1(n_135),
.B2(n_134),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_95),
.B1(n_90),
.B2(n_91),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_146),
.B1(n_126),
.B2(n_134),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_159),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_94),
.B(n_101),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_142),
.B(n_149),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_137),
.B(n_132),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_105),
.B1(n_103),
.B2(n_109),
.Y(n_146)
);

OAI22x1_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_107),
.B1(n_110),
.B2(n_90),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_161),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_106),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_127),
.B(n_19),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_111),
.C(n_101),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_164),
.C(n_18),
.Y(n_188)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_107),
.B1(n_86),
.B2(n_70),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_97),
.C(n_92),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_177),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_125),
.Y(n_170)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_150),
.B1(n_145),
.B2(n_155),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_183),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_130),
.B(n_122),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_147),
.B1(n_151),
.B2(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_127),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_184),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_30),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_141),
.B(n_114),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_181),
.B(n_190),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_119),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_169),
.C(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_63),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_67),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_168),
.B1(n_175),
.B2(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_151),
.B1(n_142),
.B2(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_182),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_159),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_18),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_191),
.B1(n_179),
.B2(n_181),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_145),
.B1(n_150),
.B2(n_103),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_213),
.C(n_186),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_92),
.C(n_50),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_188),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_70),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_119),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_26),
.Y(n_258)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_223),
.C(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_186),
.C(n_180),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_171),
.B(n_172),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_227),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_170),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_182),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_211),
.C(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_192),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_193),
.B(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_105),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_196),
.B1(n_199),
.B2(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_194),
.B(n_12),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_214),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_103),
.C(n_105),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_239),
.C(n_210),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_199),
.C(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_230),
.B1(n_220),
.B2(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_194),
.CI(n_222),
.CON(n_245),
.SN(n_245)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_8),
.Y(n_274)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_20),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_210),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_251),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_212),
.B1(n_208),
.B2(n_204),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_219),
.B1(n_30),
.B2(n_28),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_24),
.B(n_2),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_8),
.B(n_11),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_26),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_24),
.C(n_26),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_10),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_30),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_238),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_277),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_272),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_24),
.B1(n_10),
.B2(n_14),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_268),
.C(n_260),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_245),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_274),
.B(n_279),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_26),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_7),
.C(n_11),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_249),
.C(n_246),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_288),
.C(n_290),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_246),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_291),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_243),
.B(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_263),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_251),
.B(n_252),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_254),
.C(n_242),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_245),
.C(n_259),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_258),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_255),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_7),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_279),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_265),
.C(n_263),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_281),
.C(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_305),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_7),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_26),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_307),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_30),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_28),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_309),
.A2(n_310),
.B(n_313),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_294),
.B(n_20),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_20),
.B(n_17),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_301),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_295),
.A2(n_20),
.B(n_17),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_17),
.C(n_28),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_300),
.A2(n_1),
.B(n_2),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_311),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_296),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_301),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_284),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_324),
.CI(n_321),
.CON(n_328),
.SN(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_325),
.B(n_327),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_328),
.C(n_323),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_323),
.B(n_3),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_1),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_3),
.B(n_5),
.Y(n_333)
);


endmodule