module real_jpeg_27710_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_1),
.A2(n_18),
.B(n_20),
.C(n_21),
.D(n_29),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_1),
.B(n_25),
.Y(n_79)
);

A2O1A1O1Ixp25_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_25),
.B(n_37),
.C(n_79),
.D(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_1),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_1),
.A2(n_56),
.B(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_36),
.B1(n_42),
.B2(n_45),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_4),
.A2(n_42),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_5),
.A2(n_31),
.B1(n_42),
.B2(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_25),
.B(n_38),
.C(n_41),
.Y(n_37)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_10),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_75),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_62),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_15),
.B(n_62),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_16),
.Y(n_110)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_33),
.CI(n_48),
.CON(n_16),
.SN(n_16)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_28)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI32xp33_ASAP7_75t_L g59 ( 
.A1(n_19),
.A2(n_20),
.A3(n_25),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_24),
.B(n_26),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g78 ( 
.A1(n_24),
.A2(n_40),
.A3(n_45),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_41),
.B2(n_46),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_64),
.B(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_42),
.Y(n_80)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2x1_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_45),
.B(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_99),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.C(n_70),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_68),
.B1(n_69),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_86),
.B(n_108),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_81),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_96),
.B(n_107),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_94),
.B(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_102),
.B(n_106),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);


endmodule