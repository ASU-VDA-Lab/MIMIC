module fake_jpeg_15678_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.C(n_1),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_22),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_60),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_21),
.B1(n_23),
.B2(n_33),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_21),
.B1(n_19),
.B2(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_33),
.B1(n_27),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_29),
.B1(n_27),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_17),
.B1(n_28),
.B2(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_69),
.Y(n_101)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_35),
.B(n_31),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_24),
.B(n_25),
.Y(n_100)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_31),
.B1(n_20),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_86),
.B1(n_91),
.B2(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_19),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_77),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_34),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_89),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_32),
.B1(n_28),
.B2(n_41),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_98)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_34),
.B1(n_14),
.B2(n_15),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_44),
.B1(n_43),
.B2(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_34),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_18),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_62),
.B(n_65),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_77),
.B1(n_71),
.B2(n_76),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_40),
.B1(n_36),
.B2(n_42),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_113),
.B1(n_99),
.B2(n_121),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_40),
.B1(n_29),
.B2(n_27),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_120),
.B1(n_124),
.B2(n_68),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_18),
.B1(n_13),
.B2(n_12),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_128),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_38),
.C(n_25),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_79),
.C(n_67),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_24),
.B1(n_18),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_24),
.B1(n_18),
.B2(n_4),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_0),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_130),
.A2(n_135),
.B1(n_146),
.B2(n_147),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_133),
.B(n_134),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_97),
.C(n_66),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_115),
.C(n_124),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_101),
.B(n_13),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_143),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_12),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_63),
.B(n_81),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_89),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_77),
.B1(n_92),
.B2(n_84),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_88),
.B1(n_72),
.B2(n_4),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_150),
.B1(n_121),
.B2(n_118),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_72),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_106),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_148),
.B1(n_150),
.B2(n_135),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_113),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_116),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_128),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_100),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_104),
.B1(n_125),
.B2(n_119),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_104),
.A3(n_117),
.B1(n_111),
.B2(n_119),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_158),
.B(n_169),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_174),
.B(n_129),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_180),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_176),
.C(n_186),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_110),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_131),
.B(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_116),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_152),
.B1(n_156),
.B2(n_147),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_134),
.A2(n_105),
.B1(n_122),
.B2(n_123),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_183),
.A2(n_129),
.B1(n_1),
.B2(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_122),
.C(n_123),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_116),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_0),
.C(n_1),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_176),
.B1(n_184),
.B2(n_185),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_130),
.B1(n_151),
.B2(n_146),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_180),
.B1(n_172),
.B2(n_183),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_153),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_182),
.B(n_170),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_143),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_203),
.C(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_129),
.B1(n_139),
.B2(n_4),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_163),
.B1(n_175),
.B2(n_162),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_18),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_214),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_1),
.Y(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_11),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_165),
.B(n_5),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_217),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_157),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_5),
.C(n_6),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_7),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_158),
.B(n_5),
.CI(n_6),
.CON(n_217),
.SN(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_7),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_222),
.B1(n_229),
.B2(n_242),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_227),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_160),
.B1(n_187),
.B2(n_9),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_210),
.C(n_216),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_237),
.Y(n_246)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_7),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_171),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_189),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_195),
.B1(n_198),
.B2(n_194),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_206),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_248),
.B(n_254),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_255),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_251),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_253),
.C(n_257),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_206),
.C(n_192),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_192),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_197),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_227),
.B(n_207),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_259),
.C(n_260),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_203),
.C(n_212),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_190),
.C(n_193),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_188),
.C(n_200),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_263),
.C(n_230),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_217),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_270),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_219),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_224),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_242),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_272),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_231),
.Y(n_272)
);

A2O1A1O1Ixp25_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_204),
.B(n_240),
.C(n_217),
.D(n_228),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_277),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_236),
.CI(n_228),
.CON(n_276),
.SN(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_244),
.Y(n_288)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_245),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_226),
.B1(n_231),
.B2(n_209),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_240),
.B(n_230),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_272),
.B1(n_269),
.B2(n_266),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_239),
.B(n_235),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_280),
.A2(n_226),
.B(n_202),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_253),
.C(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_289),
.Y(n_308)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_276),
.B1(n_273),
.B2(n_282),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_278),
.B(n_238),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_295),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_281),
.B(n_267),
.Y(n_300)
);

NAND2x1_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_243),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_268),
.B(n_276),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_259),
.C(n_252),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_233),
.C(n_208),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_279),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_304),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_283),
.C(n_287),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_280),
.B(n_271),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_302),
.B(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_283),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_274),
.B1(n_282),
.B2(n_10),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_274),
.B1(n_9),
.B2(n_10),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_297),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_310),
.C(n_317),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_294),
.B(n_290),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_316),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_305),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_296),
.B(n_284),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_319),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_314),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_324),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_323),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_320),
.Y(n_330)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

AOI321xp33_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_318),
.A3(n_327),
.B1(n_326),
.B2(n_313),
.C(n_295),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_329),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_333),
.Y(n_334)
);


endmodule