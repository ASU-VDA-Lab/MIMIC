module real_jpeg_23438_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_39),
.B1(n_42),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_1),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_2),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_70),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_4),
.A2(n_27),
.B1(n_39),
.B2(n_42),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_27),
.B1(n_65),
.B2(n_66),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_39),
.B1(n_42),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_7),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_7),
.A2(n_48),
.B1(n_65),
.B2(n_66),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_11),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_12),
.B(n_30),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_12),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_12),
.B(n_38),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_12),
.B(n_51),
.C(n_52),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_12),
.A2(n_39),
.B1(n_42),
.B2(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_12),
.B(n_106),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_156),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_12),
.B(n_65),
.C(n_78),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_12),
.A2(n_67),
.B(n_218),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_14),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_83),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_14),
.A2(n_39),
.B1(n_42),
.B2(n_83),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_15),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_15),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_15),
.A2(n_44),
.B1(n_65),
.B2(n_66),
.Y(n_217)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_16),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_20),
.B(n_115),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.C(n_96),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_21),
.A2(n_22),
.B1(n_84),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_25),
.B(n_45),
.C(n_60),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_38),
.B2(n_43),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_26),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_28),
.A2(n_35),
.A3(n_42),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_29),
.Y(n_155)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_32),
.B(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_32),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_32),
.A2(n_133),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_34),
.B(n_39),
.Y(n_114)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_37),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_37),
.B(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_39),
.B(n_181),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_43),
.Y(n_130)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_54),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_47),
.A2(n_49),
.B1(n_58),
.B2(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_49),
.A2(n_54),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_51),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_51),
.B(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_55),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_57),
.A2(n_104),
.B1(n_106),
.B2(n_146),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_58),
.A2(n_105),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_74),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_61),
.B(n_74),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_89),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_68),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_66),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_66),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_69),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_67),
.A2(n_71),
.B(n_86),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_67),
.A2(n_111),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_67),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_67),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_71),
.B(n_156),
.Y(n_242)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_75),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_75),
.A2(n_206),
.B(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_92),
.B1(n_93),
.B2(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_76),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_76),
.A2(n_93),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_80),
.A2(n_81),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_80),
.A2(n_149),
.B(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_80),
.B(n_156),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_84),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_89),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_93),
.B(n_150),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_96),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.C(n_107),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_97),
.B(n_102),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_107),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_112),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_109),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_135),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_134),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B(n_132),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_173),
.B(n_260),
.C(n_265),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_167),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_158),
.C(n_159),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_141),
.A2(n_142),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_151),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_147),
.C(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B(n_157),
.Y(n_152)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_158),
.B(n_159),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_254),
.B(n_259),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_207),
.B(n_253),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_196),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_196),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.C(n_193),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_182),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B(n_187),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_186),
.A2(n_230),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_189),
.A2(n_193),
.B1(n_194),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_203),
.C(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_247),
.B(n_252),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_226),
.B(n_246),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_220),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_220),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_235),
.B(n_245),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_233),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_244),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_258),
.Y(n_259)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);


endmodule