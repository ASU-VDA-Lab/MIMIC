module fake_netlist_1_4391_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
BUFx6f_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
HB1xp67_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
AOI221xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_4), .B1(n_5), .B2(n_1), .C(n_2), .Y(n_8) );
HB1xp67_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_9), .B(n_4), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_4), .B(n_2), .Y(n_11) );
endmodule