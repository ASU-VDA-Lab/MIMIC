module real_aes_2802_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_449;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_0), .B(n_487), .Y(n_501) );
AOI22xp5_ASAP7_75t_SL g780 ( .A1(n_1), .A2(n_781), .B1(n_784), .B2(n_785), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_1), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_2), .A2(n_486), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_3), .B(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_4), .B(n_276), .Y(n_512) );
INVx1_ASAP7_75t_L g150 ( .A(n_5), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_6), .B(n_169), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_7), .B(n_276), .Y(n_541) );
INVx1_ASAP7_75t_L g178 ( .A(n_8), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g792 ( .A(n_9), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_10), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g582 ( .A(n_11), .B(n_273), .Y(n_582) );
INVx2_ASAP7_75t_L g139 ( .A(n_12), .Y(n_139) );
AOI221x1_ASAP7_75t_L g485 ( .A1(n_13), .A2(n_26), .B1(n_486), .B2(n_487), .C(n_488), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_14), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_15), .B(n_487), .Y(n_578) );
INVx1_ASAP7_75t_L g274 ( .A(n_16), .Y(n_274) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_17), .A2(n_175), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_18), .B(n_221), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_19), .B(n_276), .Y(n_565) );
AO21x1_ASAP7_75t_L g507 ( .A1(n_20), .A2(n_487), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g118 ( .A(n_21), .Y(n_118) );
NOR2xp33_ASAP7_75t_SL g789 ( .A(n_21), .B(n_119), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_22), .Y(n_120) );
INVx1_ASAP7_75t_L g271 ( .A(n_23), .Y(n_271) );
INVx1_ASAP7_75t_SL g236 ( .A(n_24), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_25), .B(n_156), .Y(n_257) );
AOI33xp33_ASAP7_75t_L g207 ( .A1(n_27), .A2(n_56), .A3(n_145), .B1(n_154), .B2(n_208), .B3(n_209), .Y(n_207) );
NAND2x1_ASAP7_75t_L g499 ( .A(n_28), .B(n_276), .Y(n_499) );
NAND2x1_ASAP7_75t_L g540 ( .A(n_29), .B(n_273), .Y(n_540) );
INVx1_ASAP7_75t_L g187 ( .A(n_30), .Y(n_187) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_31), .A2(n_89), .B(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g170 ( .A(n_31), .B(n_89), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_32), .B(n_164), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_33), .B(n_273), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_34), .A2(n_94), .B1(n_762), .B2(n_763), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_34), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_35), .B(n_276), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_36), .B(n_273), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_37), .A2(n_486), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g144 ( .A(n_38), .Y(n_144) );
AND2x2_ASAP7_75t_L g162 ( .A(n_38), .B(n_150), .Y(n_162) );
AND2x2_ASAP7_75t_L g168 ( .A(n_38), .B(n_147), .Y(n_168) );
OR2x6_ASAP7_75t_L g116 ( .A(n_39), .B(n_117), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g790 ( .A(n_39), .B(n_114), .C(n_791), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_40), .A2(n_760), .B1(n_765), .B2(n_770), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_41), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_42), .A2(n_53), .B1(n_782), .B2(n_783), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_42), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_43), .B(n_487), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_44), .B(n_164), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_45), .A2(n_137), .B1(n_169), .B2(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_46), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_47), .B(n_156), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_48), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_49), .B(n_273), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_50), .B(n_175), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_51), .B(n_156), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_52), .A2(n_486), .B(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_53), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_54), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_55), .B(n_273), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_57), .B(n_156), .Y(n_219) );
INVx1_ASAP7_75t_L g149 ( .A(n_58), .Y(n_149) );
INVx1_ASAP7_75t_L g158 ( .A(n_58), .Y(n_158) );
AND2x2_ASAP7_75t_L g220 ( .A(n_59), .B(n_221), .Y(n_220) );
AOI221xp5_ASAP7_75t_L g176 ( .A1(n_60), .A2(n_77), .B1(n_142), .B2(n_164), .C(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_61), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_62), .B(n_276), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_63), .B(n_137), .Y(n_197) );
AOI21xp5_ASAP7_75t_SL g141 ( .A1(n_64), .A2(n_142), .B(n_151), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_65), .A2(n_486), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g268 ( .A(n_66), .Y(n_268) );
AO21x1_ASAP7_75t_L g509 ( .A1(n_67), .A2(n_486), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_68), .B(n_487), .Y(n_530) );
INVx1_ASAP7_75t_L g218 ( .A(n_69), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_70), .B(n_487), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_71), .A2(n_142), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g523 ( .A(n_72), .B(n_222), .Y(n_523) );
INVx1_ASAP7_75t_L g147 ( .A(n_73), .Y(n_147) );
INVx1_ASAP7_75t_L g160 ( .A(n_73), .Y(n_160) );
AND2x2_ASAP7_75t_L g543 ( .A(n_74), .B(n_136), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_75), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_76), .B(n_164), .Y(n_210) );
AND2x2_ASAP7_75t_L g238 ( .A(n_78), .B(n_136), .Y(n_238) );
INVx1_ASAP7_75t_L g269 ( .A(n_79), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_80), .A2(n_142), .B(n_235), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_81), .A2(n_142), .B(n_202), .C(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
AND2x2_ASAP7_75t_L g528 ( .A(n_83), .B(n_136), .Y(n_528) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_84), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_85), .B(n_487), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_86), .A2(n_142), .B1(n_205), .B2(n_206), .Y(n_204) );
XNOR2xp5_ASAP7_75t_L g760 ( .A(n_87), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g508 ( .A(n_88), .B(n_169), .Y(n_508) );
AND2x2_ASAP7_75t_L g502 ( .A(n_90), .B(n_136), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_91), .B(n_273), .Y(n_566) );
INVx1_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_93), .B(n_276), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_94), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_95), .B(n_273), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_96), .A2(n_486), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g211 ( .A(n_97), .B(n_136), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_98), .B(n_276), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_99), .A2(n_185), .B(n_186), .C(n_189), .Y(n_184) );
BUFx2_ASAP7_75t_L g123 ( .A(n_100), .Y(n_123) );
BUFx2_ASAP7_75t_SL g776 ( .A(n_100), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_101), .A2(n_486), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_102), .B(n_156), .Y(n_155) );
AOI21xp33_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_786), .B(n_793), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI21x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_124), .B(n_774), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_121), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_108), .A2(n_778), .B(n_779), .Y(n_777) );
NOR2xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_120), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_112), .Y(n_778) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OR2x6_ASAP7_75t_SL g473 ( .A(n_114), .B(n_115), .Y(n_473) );
AND2x6_ASAP7_75t_SL g477 ( .A(n_114), .B(n_116), .Y(n_477) );
OR2x2_ASAP7_75t_L g773 ( .A(n_114), .B(n_116), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_760), .B(n_764), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_471), .B1(n_474), .B2(n_478), .Y(n_126) );
INVx2_ASAP7_75t_L g769 ( .A(n_127), .Y(n_769) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NAND3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_361), .C(n_426), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_315), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_260), .B(n_288), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_223), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_171), .Y(n_132) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_133), .A2(n_363), .B(n_374), .Y(n_362) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_133), .B(n_304), .Y(n_397) );
AND2x2_ASAP7_75t_L g412 ( .A(n_133), .B(n_413), .Y(n_412) );
OR2x6_ASAP7_75t_L g422 ( .A(n_133), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g424 ( .A(n_133), .B(n_414), .Y(n_424) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g298 ( .A(n_134), .Y(n_298) );
AND2x2_ASAP7_75t_L g311 ( .A(n_134), .B(n_312), .Y(n_311) );
INVx4_ASAP7_75t_L g330 ( .A(n_134), .Y(n_330) );
AND2x2_ASAP7_75t_L g333 ( .A(n_134), .B(n_249), .Y(n_333) );
NOR2x1_ASAP7_75t_SL g336 ( .A(n_134), .B(n_264), .Y(n_336) );
AND2x4_ASAP7_75t_L g348 ( .A(n_134), .B(n_346), .Y(n_348) );
OR2x2_ASAP7_75t_L g358 ( .A(n_134), .B(n_230), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_134), .B(n_370), .Y(n_375) );
OR2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_136), .A2(n_184), .B1(n_190), .B2(n_191), .Y(n_183) );
INVx3_ASAP7_75t_L g191 ( .A(n_136), .Y(n_191) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_137), .B(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_138), .Y(n_175) );
AND2x4_ASAP7_75t_L g169 ( .A(n_139), .B(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_139), .B(n_170), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_163), .B(n_169), .Y(n_140) );
INVxp67_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
NOR2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx1_ASAP7_75t_L g209 ( .A(n_145), .Y(n_209) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x6_ASAP7_75t_L g153 ( .A(n_146), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g273 ( .A(n_147), .B(n_157), .Y(n_273) );
AND2x6_ASAP7_75t_L g486 ( .A(n_148), .B(n_168), .Y(n_486) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
INVx2_ASAP7_75t_L g154 ( .A(n_149), .Y(n_154) );
AND2x4_ASAP7_75t_L g276 ( .A(n_149), .B(n_159), .Y(n_276) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_155), .C(n_161), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_153), .A2(n_161), .B(n_178), .C(n_179), .Y(n_177) );
INVxp67_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_153), .A2(n_161), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_153), .A2(n_161), .B(n_236), .C(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g259 ( .A(n_153), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_153), .A2(n_188), .B1(n_268), .B2(n_269), .Y(n_267) );
AND2x2_ASAP7_75t_L g165 ( .A(n_154), .B(n_166), .Y(n_165) );
INVxp33_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
INVx1_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
AND2x4_ASAP7_75t_L g487 ( .A(n_156), .B(n_162), .Y(n_487) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_161), .A2(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_161), .B(n_169), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_161), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_161), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_161), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_161), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_161), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_161), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_161), .A2(n_565), .B(n_566), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_161), .A2(n_581), .B(n_582), .Y(n_580) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
INVx1_ASAP7_75t_L g198 ( .A(n_164), .Y(n_198) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_167), .Y(n_164) );
INVx1_ASAP7_75t_L g252 ( .A(n_165), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_167), .Y(n_253) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_169), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_SL g561 ( .A(n_169), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_169), .A2(n_578), .B(n_579), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_171), .A2(n_304), .B1(n_399), .B2(n_400), .Y(n_398) );
INVx1_ASAP7_75t_SL g442 ( .A(n_171), .Y(n_442) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_199), .Y(n_171) );
INVx2_ASAP7_75t_L g373 ( .A(n_172), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_172), .B(n_319), .Y(n_445) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_181), .Y(n_172) );
BUFx3_ASAP7_75t_L g291 ( .A(n_173), .Y(n_291) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g284 ( .A(n_174), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_174), .B(n_201), .Y(n_306) );
AND2x4_ASAP7_75t_L g323 ( .A(n_174), .B(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_L g339 ( .A(n_174), .Y(n_339) );
INVx2_ASAP7_75t_L g396 ( .A(n_174), .Y(n_396) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_180), .Y(n_174) );
INVx2_ASAP7_75t_SL g202 ( .A(n_175), .Y(n_202) );
AND2x2_ASAP7_75t_L g314 ( .A(n_181), .B(n_280), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g360 ( .A(n_181), .B(n_283), .Y(n_360) );
AND2x2_ASAP7_75t_L g379 ( .A(n_181), .B(n_283), .Y(n_379) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g241 ( .A(n_182), .Y(n_241) );
INVx1_ASAP7_75t_L g322 ( .A(n_182), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_182), .B(n_213), .Y(n_341) );
AND2x4_ASAP7_75t_L g395 ( .A(n_182), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_192), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_191), .A2(n_214), .B(n_220), .Y(n_213) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_191), .A2(n_214), .B(n_220), .Y(n_283) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_191), .A2(n_496), .B(n_502), .Y(n_495) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_191), .A2(n_517), .B(n_523), .Y(n_516) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_191), .A2(n_517), .B(n_523), .Y(n_550) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_191), .A2(n_496), .B(n_502), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g354 ( .A(n_199), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_199), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_212), .Y(n_199) );
AND2x2_ASAP7_75t_L g338 ( .A(n_200), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g378 ( .A(n_200), .Y(n_378) );
AND2x2_ASAP7_75t_L g383 ( .A(n_200), .B(n_283), .Y(n_383) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_201), .B(n_213), .Y(n_243) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_201) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_204), .B(n_210), .Y(n_203) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g319 ( .A(n_212), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_212), .B(n_291), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_212), .B(n_241), .Y(n_458) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_213), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_221), .Y(n_231) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_221), .A2(n_485), .B(n_491), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_221), .A2(n_530), .B(n_531), .Y(n_529) );
OA21x2_ASAP7_75t_L g630 ( .A1(n_221), .A2(n_485), .B(n_491), .Y(n_630) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OAI21xp33_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_239), .B(n_244), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_226), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g296 ( .A(n_227), .Y(n_296) );
AND2x2_ASAP7_75t_L g310 ( .A(n_227), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g344 ( .A(n_227), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g410 ( .A(n_227), .B(n_328), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g456 ( .A(n_227), .B(n_457), .C(n_458), .Y(n_456) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_228), .Y(n_287) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g303 ( .A(n_230), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_230), .B(n_264), .Y(n_309) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_230), .Y(n_320) );
AND2x2_ASAP7_75t_L g365 ( .A(n_230), .B(n_263), .Y(n_365) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_230), .Y(n_388) );
INVx1_ASAP7_75t_L g405 ( .A(n_230), .Y(n_405) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_238), .Y(n_230) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_231), .A2(n_537), .B(n_543), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g447 ( .A(n_239), .Y(n_447) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_240), .B(n_318), .Y(n_419) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g281 ( .A(n_241), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AOI211x1_ASAP7_75t_L g315 ( .A1(n_245), .A2(n_316), .B(n_325), .C(n_342), .Y(n_315) );
INVx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_246), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g368 ( .A(n_246), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g304 ( .A(n_248), .B(n_263), .Y(n_304) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x4_ASAP7_75t_L g262 ( .A(n_249), .B(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_249), .Y(n_329) );
INVx1_ASAP7_75t_L g346 ( .A(n_249), .Y(n_346) );
AND2x2_ASAP7_75t_L g414 ( .A(n_249), .B(n_264), .Y(n_414) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_255), .Y(n_249) );
NOR3xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .C(n_254), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_278), .B(n_285), .Y(n_260) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_261), .B(n_330), .Y(n_433) );
INVx2_ASAP7_75t_L g465 ( .A(n_261), .Y(n_465) );
INVx4_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g297 ( .A(n_262), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g370 ( .A(n_263), .Y(n_370) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g312 ( .A(n_264), .Y(n_312) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B(n_277), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_274), .B2(n_275), .Y(n_270) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
OR2x2_ASAP7_75t_L g372 ( .A(n_279), .B(n_373), .Y(n_372) );
NAND2x1_ASAP7_75t_SL g394 ( .A(n_279), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g294 ( .A(n_280), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g324 ( .A(n_280), .Y(n_324) );
INVx1_ASAP7_75t_L g448 ( .A(n_281), .Y(n_448) );
AND2x2_ASAP7_75t_L g313 ( .A(n_282), .B(n_314), .Y(n_313) );
NOR2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g295 ( .A(n_283), .Y(n_295) );
INVxp33_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g352 ( .A(n_287), .B(n_345), .Y(n_352) );
OAI211xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_292), .B(n_299), .C(n_307), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g376 ( .A(n_290), .B(n_377), .Y(n_376) );
NOR2xp67_ASAP7_75t_SL g381 ( .A(n_290), .B(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_291), .B(n_378), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_297), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
AND2x2_ASAP7_75t_L g425 ( .A(n_294), .B(n_395), .Y(n_425) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_297), .A2(n_444), .B1(n_446), .B2(n_449), .C1(n_450), .C2(n_453), .Y(n_443) );
INVx1_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_305), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_303), .Y(n_334) );
AND2x4_ASAP7_75t_SL g369 ( .A(n_303), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g423 ( .A(n_304), .Y(n_423) );
AND2x2_ASAP7_75t_L g468 ( .A(n_304), .B(n_320), .Y(n_468) );
AND2x2_ASAP7_75t_L g349 ( .A(n_305), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g462 ( .A(n_306), .B(n_341), .Y(n_462) );
OAI21xp33_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_310), .B(n_313), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_308), .A2(n_328), .B(n_369), .Y(n_429) );
AND2x2_ASAP7_75t_L g453 ( .A(n_309), .B(n_330), .Y(n_453) );
NOR2xp33_ASAP7_75t_SL g463 ( .A(n_309), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g401 ( .A(n_312), .Y(n_401) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_312), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g436 ( .A(n_314), .Y(n_436) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_321), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g439 ( .A(n_319), .B(n_323), .Y(n_439) );
BUFx2_ASAP7_75t_L g327 ( .A(n_320), .Y(n_327) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g350 ( .A(n_322), .Y(n_350) );
INVx2_ASAP7_75t_L g356 ( .A(n_322), .Y(n_356) );
AND2x2_ASAP7_75t_L g392 ( .A(n_322), .B(n_383), .Y(n_392) );
AND2x4_ASAP7_75t_L g359 ( .A(n_323), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g399 ( .A(n_323), .B(n_356), .Y(n_399) );
AND2x2_ASAP7_75t_L g450 ( .A(n_323), .B(n_451), .Y(n_450) );
AOI31xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_331), .A3(n_335), .B(n_337), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g347 ( .A(n_327), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_SL g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g345 ( .A(n_330), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_333), .A2(n_385), .B1(n_416), .B2(n_419), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_333), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g470 ( .A(n_333), .B(n_386), .Y(n_470) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g385 ( .A(n_336), .B(n_386), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AND2x2_ASAP7_75t_L g408 ( .A(n_338), .B(n_379), .Y(n_408) );
INVx1_ASAP7_75t_L g418 ( .A(n_340), .Y(n_418) );
INVx2_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_351), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B(n_349), .Y(n_343) );
INVx1_ASAP7_75t_L g441 ( .A(n_344), .Y(n_441) );
AND2x2_ASAP7_75t_L g449 ( .A(n_345), .B(n_401), .Y(n_449) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_345), .Y(n_455) );
AND2x2_ASAP7_75t_L g400 ( .A(n_348), .B(n_401), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_353), .B1(n_357), .B2(n_359), .Y(n_351) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_355), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_354), .A2(n_373), .B1(n_467), .B2(n_469), .Y(n_466) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g366 ( .A(n_359), .Y(n_366) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_389), .Y(n_361) );
OAI21xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B(n_367), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_365), .A2(n_368), .B(n_371), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_368), .A2(n_392), .B1(n_393), .B2(n_397), .Y(n_391) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_380), .B2(n_384), .Y(n_374) );
INVx1_ASAP7_75t_L g409 ( .A(n_377), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g389 ( .A(n_390), .B(n_402), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_398), .Y(n_390) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
NAND2xp33_ASAP7_75t_SL g444 ( .A(n_394), .B(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g417 ( .A(n_395), .Y(n_417) );
INVx3_ASAP7_75t_L g431 ( .A(n_399), .Y(n_431) );
INVxp67_ASAP7_75t_L g460 ( .A(n_400), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_403), .B(n_411), .C(n_415), .D(n_420), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_408), .B1(n_409), .B2(n_410), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g413 ( .A(n_405), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g461 ( .A(n_409), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_424), .B(n_425), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND3x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_443), .C(n_454), .Y(n_426) );
AOI221x1_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_432), .B2(n_434), .C(n_440), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp33_ASAP7_75t_SL g434 ( .A(n_435), .B(n_438), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
NAND2xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_459), .C(n_466), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_459) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_472), .Y(n_768) );
CKINVDCx11_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
CKINVDCx6p67_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
CKINVDCx11_ASAP7_75t_R g766 ( .A(n_475), .Y(n_766) );
INVx3_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g767 ( .A(n_478), .Y(n_767) );
XNOR2x2_ASAP7_75t_SL g779 ( .A(n_478), .B(n_780), .Y(n_779) );
NAND4xp75_ASAP7_75t_L g478 ( .A(n_479), .B(n_670), .C(n_710), .D(n_739), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_632), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_589), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_524), .B(n_544), .Y(n_481) );
AND2x2_ASAP7_75t_SL g482 ( .A(n_483), .B(n_492), .Y(n_482) );
AND2x4_ASAP7_75t_L g588 ( .A(n_483), .B(n_549), .Y(n_588) );
INVx1_ASAP7_75t_SL g641 ( .A(n_483), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_483), .A2(n_677), .B(n_680), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_SL g680 ( .A1(n_483), .A2(n_681), .B(n_682), .C(n_683), .Y(n_680) );
NAND2x1_ASAP7_75t_L g721 ( .A(n_483), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_483), .B(n_682), .Y(n_743) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g547 ( .A(n_484), .Y(n_547) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_484), .Y(n_620) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_503), .Y(n_492) );
AND2x2_ASAP7_75t_L g612 ( .A(n_493), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g693 ( .A(n_493), .B(n_549), .Y(n_693) );
INVx1_ASAP7_75t_L g753 ( .A(n_493), .Y(n_753) );
BUFx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g597 ( .A(n_494), .B(n_515), .Y(n_597) );
AND2x2_ASAP7_75t_L g722 ( .A(n_494), .B(n_516), .Y(n_722) );
AND2x2_ASAP7_75t_L g727 ( .A(n_494), .B(n_687), .Y(n_727) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVxp67_ASAP7_75t_L g603 ( .A(n_495), .Y(n_603) );
BUFx3_ASAP7_75t_L g636 ( .A(n_495), .Y(n_636) );
AND2x2_ASAP7_75t_L g682 ( .A(n_495), .B(n_516), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
AND2x2_ASAP7_75t_L g667 ( .A(n_503), .B(n_546), .Y(n_667) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
AND2x4_ASAP7_75t_L g549 ( .A(n_504), .B(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g659 ( .A(n_504), .B(n_643), .Y(n_659) );
AND2x2_ASAP7_75t_SL g702 ( .A(n_504), .B(n_630), .Y(n_702) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g638 ( .A(n_505), .Y(n_638) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g599 ( .A(n_506), .Y(n_599) );
OAI21x1_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_509), .B(n_513), .Y(n_506) );
INVx1_ASAP7_75t_L g514 ( .A(n_508), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_515), .B(n_599), .Y(n_602) );
AND2x2_ASAP7_75t_L g687 ( .A(n_515), .B(n_630), .Y(n_687) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g684 ( .A(n_516), .B(n_547), .Y(n_684) );
AND2x2_ASAP7_75t_L g704 ( .A(n_516), .B(n_630), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_518), .B(n_522), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_524), .B(n_593), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_524), .A2(n_716), .B1(n_717), .B2(n_718), .C(n_720), .Y(n_715) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI332xp33_ASAP7_75t_L g749 ( .A1(n_525), .A2(n_609), .A3(n_616), .B1(n_675), .B2(n_750), .B3(n_751), .C1(n_752), .C2(n_754), .Y(n_749) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_526), .B(n_535), .Y(n_525) );
AND2x2_ASAP7_75t_L g555 ( .A(n_526), .B(n_536), .Y(n_555) );
AND2x2_ASAP7_75t_L g572 ( .A(n_526), .B(n_573), .Y(n_572) );
INVx4_ASAP7_75t_L g584 ( .A(n_526), .Y(n_584) );
AND2x2_ASAP7_75t_SL g644 ( .A(n_526), .B(n_585), .Y(n_644) );
INVx5_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NOR2x1_ASAP7_75t_SL g606 ( .A(n_527), .B(n_573), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_527), .B(n_535), .Y(n_610) );
AND2x2_ASAP7_75t_L g617 ( .A(n_527), .B(n_536), .Y(n_617) );
BUFx2_ASAP7_75t_L g652 ( .A(n_527), .Y(n_652) );
AND2x2_ASAP7_75t_L g707 ( .A(n_527), .B(n_576), .Y(n_707) );
OR2x6_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
OR2x2_ASAP7_75t_L g575 ( .A(n_535), .B(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g585 ( .A(n_535), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g625 ( .A(n_535), .Y(n_625) );
AND2x2_ASAP7_75t_L g695 ( .A(n_535), .B(n_594), .Y(n_695) );
AND2x2_ASAP7_75t_L g708 ( .A(n_535), .B(n_709), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_535), .B(n_709), .Y(n_726) );
INVx4_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_536), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
OAI32xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_551), .A3(n_556), .B1(n_570), .B2(n_587), .Y(n_544) );
INVx2_ASAP7_75t_L g653 ( .A(n_545), .Y(n_653) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
INVx1_ASAP7_75t_L g664 ( .A(n_546), .Y(n_664) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g598 ( .A(n_547), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g731 ( .A(n_547), .B(n_636), .Y(n_731) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g643 ( .A(n_550), .Y(n_643) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx2_ASAP7_75t_L g631 ( .A(n_553), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_553), .B(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_SL g642 ( .A(n_554), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g719 ( .A(n_554), .Y(n_719) );
AND2x2_ASAP7_75t_L g737 ( .A(n_554), .B(n_599), .Y(n_737) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NOR2xp67_ASAP7_75t_SL g681 ( .A(n_557), .B(n_610), .Y(n_681) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_558), .B(n_592), .Y(n_679) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g755 ( .A(n_559), .B(n_625), .Y(n_755) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g586 ( .A(n_560), .Y(n_586) );
INVx2_ASAP7_75t_L g627 ( .A(n_560), .Y(n_627) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_568), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_561), .B(n_569), .Y(n_568) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_561), .A2(n_562), .B(n_568), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_583), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_571), .B(n_629), .Y(n_714) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND3x2_ASAP7_75t_L g669 ( .A(n_572), .B(n_616), .C(n_625), .Y(n_669) );
AND2x2_ASAP7_75t_L g593 ( .A(n_573), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_573), .B(n_576), .Y(n_650) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g604 ( .A(n_575), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g594 ( .A(n_576), .Y(n_594) );
INVx1_ASAP7_75t_L g609 ( .A(n_576), .Y(n_609) );
BUFx3_ASAP7_75t_L g616 ( .A(n_576), .Y(n_616) );
AND2x2_ASAP7_75t_L g626 ( .A(n_576), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x4_ASAP7_75t_L g635 ( .A(n_584), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_584), .B(n_594), .Y(n_678) );
AND2x2_ASAP7_75t_L g634 ( .A(n_585), .B(n_609), .Y(n_634) );
INVx2_ASAP7_75t_L g661 ( .A(n_585), .Y(n_661) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
AOI211xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_595), .B(n_600), .C(n_621), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_590), .A2(n_717), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_593), .B(n_652), .Y(n_651) );
AOI211xp5_ASAP7_75t_SL g671 ( .A1(n_593), .A2(n_672), .B(n_676), .C(n_685), .Y(n_671) );
AND2x2_ASAP7_75t_L g657 ( .A(n_594), .B(n_617), .Y(n_657) );
OR2x2_ASAP7_75t_L g660 ( .A(n_594), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_597), .B(n_702), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_598), .B(n_643), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_598), .A2(n_624), .B1(n_704), .B2(n_707), .C(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g629 ( .A(n_599), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g675 ( .A(n_599), .B(n_630), .Y(n_675) );
OAI221xp5_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_604), .B1(n_607), .B2(n_611), .C(n_614), .Y(n_600) );
AND2x2_ASAP7_75t_L g746 ( .A(n_601), .B(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g613 ( .A(n_602), .Y(n_613) );
INVx1_ASAP7_75t_L g699 ( .A(n_603), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_604), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g618 ( .A(n_606), .B(n_609), .Y(n_618) );
AND2x2_ASAP7_75t_L g694 ( .A(n_606), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g619 ( .A(n_613), .B(n_620), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_618), .B(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g738 ( .A(n_615), .Y(n_738) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g717 ( .A(n_616), .B(n_644), .Y(n_717) );
AND2x2_ASAP7_75t_SL g690 ( .A(n_617), .B(n_626), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B(n_628), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_622), .A2(n_656), .B1(n_659), .B2(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g728 ( .A(n_622), .Y(n_728) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g648 ( .A(n_625), .Y(n_648) );
INVx1_ASAP7_75t_L g709 ( .A(n_627), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_629), .B(n_699), .Y(n_750) );
AND2x2_ASAP7_75t_L g718 ( .A(n_630), .B(n_719), .Y(n_718) );
OAI211xp5_ASAP7_75t_L g711 ( .A1(n_631), .A2(n_712), .B(n_715), .C(n_723), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_654), .Y(n_632) );
AOI322xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .A3(n_637), .B1(n_639), .B2(n_644), .C1(n_645), .C2(n_653), .Y(n_633) );
CKINVDCx16_ASAP7_75t_R g751 ( .A(n_635), .Y(n_751) );
AND2x2_ASAP7_75t_L g701 ( .A(n_636), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g735 ( .A(n_636), .Y(n_735) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_SL g686 ( .A(n_638), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_SL g692 ( .A(n_638), .B(n_684), .Y(n_692) );
AND2x2_ASAP7_75t_L g716 ( .A(n_638), .B(n_682), .Y(n_716) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g688 ( .A(n_642), .Y(n_688) );
NAND2xp33_ASAP7_75t_SL g645 ( .A(n_646), .B(n_651), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_SL g691 ( .A1(n_647), .A2(n_692), .B1(n_693), .B2(n_694), .C(n_696), .Y(n_691) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g758 ( .A(n_650), .Y(n_758) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_658), .C(n_662), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g733 ( .A(n_657), .Y(n_733) );
INVx1_ASAP7_75t_L g665 ( .A(n_659), .Y(n_665) );
OR2x2_ASAP7_75t_L g752 ( .A(n_659), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g748 ( .A(n_660), .Y(n_748) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_668), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_664), .B(n_682), .Y(n_759) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_691), .Y(n_670) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_674), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OR2x2_ASAP7_75t_L g725 ( .A(n_678), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_688), .B(n_689), .Y(n_685) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
AOI31xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_700), .A3(n_703), .B(n_705), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_702), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_727), .B1(n_728), .B2(n_729), .C(n_732), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B1(n_736), .B2(n_738), .Y(n_732) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_749), .C(n_756), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_741), .B(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_748), .Y(n_744) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI22x1_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g784 ( .A(n_781), .Y(n_784) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_786), .Y(n_795) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_SL g788 ( .A(n_789), .B(n_790), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
endmodule