module fake_jpeg_8955_n_302 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_288;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_27),
.B1(n_26),
.B2(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_53),
.B1(n_62),
.B2(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_26),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_64),
.B(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_27),
.B1(n_26),
.B2(n_32),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_28),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_33),
.B1(n_31),
.B2(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_23),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_75),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_36),
.B1(n_33),
.B2(n_31),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_85),
.B1(n_50),
.B2(n_30),
.Y(n_102)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_71),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_77),
.B(n_81),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_39),
.B1(n_43),
.B2(n_37),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_66),
.B1(n_63),
.B2(n_49),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_33),
.B1(n_19),
.B2(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_39),
.B1(n_35),
.B2(n_40),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_65),
.B1(n_60),
.B2(n_48),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_19),
.B1(n_28),
.B2(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_90),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_22),
.B1(n_21),
.B2(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_37),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_115),
.B1(n_78),
.B2(n_68),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_83),
.B1(n_34),
.B2(n_17),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_R g139 ( 
.A(n_102),
.B(n_118),
.Y(n_139)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_39),
.B(n_47),
.C(n_35),
.D(n_49),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_40),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_35),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_120),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_35),
.B1(n_34),
.B2(n_17),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_72),
.B1(n_84),
.B2(n_71),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_74),
.C(n_80),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_25),
.C(n_34),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_37),
.B1(n_59),
.B2(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_121),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_37),
.B(n_24),
.C(n_35),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_44),
.A3(n_40),
.B1(n_67),
.B2(n_20),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_40),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_136),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_24),
.B(n_25),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_106),
.B(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_134),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_86),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_89),
.Y(n_131)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_55),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_147),
.B1(n_100),
.B2(n_113),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_143),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_25),
.B(n_68),
.C(n_72),
.Y(n_141)
);

AO22x2_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_118),
.B1(n_99),
.B2(n_101),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_83),
.C(n_20),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_2),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_34),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_2),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_10),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_127),
.B1(n_145),
.B2(n_133),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_150),
.B(n_103),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_157),
.B(n_163),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_170),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_115),
.B1(n_97),
.B2(n_126),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_162),
.B1(n_164),
.B2(n_168),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_109),
.B1(n_99),
.B2(n_117),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_109),
.B1(n_99),
.B2(n_108),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_172),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_128),
.A2(n_96),
.B1(n_112),
.B2(n_120),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_11),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_103),
.B1(n_112),
.B2(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_176),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_119),
.B1(n_20),
.B2(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_142),
.B1(n_146),
.B2(n_145),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_124),
.C(n_148),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_199),
.C(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_188),
.Y(n_216)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_197),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_194),
.A2(n_204),
.B(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_163),
.B1(n_175),
.B2(n_176),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx3_ASAP7_75t_SL g202 ( 
.A(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_167),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_208),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_159),
.B1(n_162),
.B2(n_168),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_209),
.A2(n_211),
.B1(n_214),
.B2(n_224),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_175),
.B(n_158),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_164),
.B1(n_171),
.B2(n_163),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_170),
.B(n_163),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_213),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_187),
.B1(n_181),
.B2(n_204),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_130),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_11),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_222),
.C(n_182),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_165),
.C(n_152),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_189),
.A2(n_163),
.B1(n_153),
.B2(n_134),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_205),
.B1(n_198),
.B2(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_153),
.B1(n_130),
.B2(n_5),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_213),
.A2(n_182),
.B(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_235),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_206),
.C(n_183),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_245),
.C(n_218),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_185),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_238),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_240),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_9),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_8),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_8),
.B(n_14),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_224),
.B1(n_211),
.B2(n_223),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_8),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_212),
.B(n_6),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_225),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_229),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_246),
.B1(n_243),
.B2(n_215),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_235),
.B(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_240),
.C(n_245),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_229),
.C(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_234),
.C(n_214),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_253),
.C(n_255),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_268),
.B(n_209),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_228),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_272),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_228),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_230),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_254),
.Y(n_275)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_283),
.C(n_248),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_272),
.A3(n_271),
.B1(n_266),
.B2(n_265),
.C1(n_217),
.C2(n_248),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_217),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_281),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_274),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_261),
.B1(n_207),
.B2(n_225),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_261),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_248),
.B(n_7),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_286),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_291),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_280),
.C(n_7),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_280),
.B(n_282),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_292),
.B(n_293),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_7),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_3),
.A3(n_12),
.B1(n_13),
.B2(n_16),
.C1(n_298),
.C2(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_12),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_13),
.Y(n_302)
);


endmodule