module real_aes_1258_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_0), .B(n_152), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_1), .A2(n_146), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_2), .B(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_3), .B(n_163), .Y(n_238) );
INVx1_ASAP7_75t_L g151 ( .A(n_4), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_5), .B(n_163), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_6), .B(n_215), .Y(n_503) );
INVx1_ASAP7_75t_L g546 ( .A(n_7), .Y(n_546) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_8), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_9), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_10), .Y(n_805) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_11), .B(n_161), .Y(n_214) );
INVx2_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
AOI221x1_ASAP7_75t_L g145 ( .A1(n_13), .A2(n_26), .B1(n_146), .B2(n_152), .C(n_159), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_14), .B(n_441), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_16), .B(n_152), .Y(n_210) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_17), .A2(n_208), .B(n_209), .Y(n_207) );
INVx1_ASAP7_75t_L g512 ( .A(n_18), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_19), .B(n_141), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_20), .B(n_163), .Y(n_222) );
AO21x1_ASAP7_75t_L g233 ( .A1(n_21), .A2(n_152), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g510 ( .A(n_23), .Y(n_510) );
INVx1_ASAP7_75t_SL g496 ( .A(n_24), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_25), .B(n_153), .Y(n_474) );
NAND2x1_ASAP7_75t_L g171 ( .A(n_27), .B(n_163), .Y(n_171) );
AOI33xp33_ASAP7_75t_L g527 ( .A1(n_28), .A2(n_56), .A3(n_462), .B1(n_471), .B2(n_528), .B3(n_529), .Y(n_527) );
NAND2x1_ASAP7_75t_L g201 ( .A(n_29), .B(n_161), .Y(n_201) );
INVx1_ASAP7_75t_L g554 ( .A(n_30), .Y(n_554) );
OR2x2_ASAP7_75t_L g144 ( .A(n_31), .B(n_90), .Y(n_144) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_31), .A2(n_90), .B(n_143), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_32), .B(n_487), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_33), .B(n_161), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_34), .A2(n_35), .B1(n_787), .B2(n_788), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_34), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_35), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_36), .B(n_163), .Y(n_213) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_37), .A2(n_38), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_37), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_38), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_39), .B(n_161), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_40), .A2(n_146), .B(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g147 ( .A(n_41), .B(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g158 ( .A(n_41), .B(n_151), .Y(n_158) );
INVx1_ASAP7_75t_L g470 ( .A(n_41), .Y(n_470) );
OR2x6_ASAP7_75t_L g112 ( .A(n_42), .B(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_43), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_44), .B(n_152), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_45), .B(n_487), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_46), .A2(n_176), .B1(n_215), .B2(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_47), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_48), .B(n_153), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_49), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_50), .B(n_161), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_51), .B(n_208), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_52), .B(n_153), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_53), .A2(n_146), .B(n_200), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_54), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_55), .B(n_161), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_57), .B(n_153), .Y(n_538) );
INVx1_ASAP7_75t_L g150 ( .A(n_58), .Y(n_150) );
INVx1_ASAP7_75t_L g155 ( .A(n_58), .Y(n_155) );
AND2x2_ASAP7_75t_L g539 ( .A(n_59), .B(n_141), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_60), .A2(n_77), .B1(n_468), .B2(n_487), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_61), .B(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_62), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_63), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_64), .B(n_176), .Y(n_562) );
AOI21xp5_ASAP7_75t_SL g482 ( .A1(n_65), .A2(n_468), .B(n_483), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_66), .A2(n_146), .B(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g506 ( .A(n_67), .Y(n_506) );
AO21x1_ASAP7_75t_L g235 ( .A1(n_68), .A2(n_146), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_69), .B(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g537 ( .A(n_70), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_71), .B(n_152), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_72), .A2(n_468), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g186 ( .A(n_73), .B(n_142), .Y(n_186) );
INVx1_ASAP7_75t_L g148 ( .A(n_74), .Y(n_148) );
INVx1_ASAP7_75t_L g157 ( .A(n_74), .Y(n_157) );
AND2x2_ASAP7_75t_L g205 ( .A(n_75), .B(n_175), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_76), .B(n_487), .Y(n_530) );
AND2x2_ASAP7_75t_L g498 ( .A(n_78), .B(n_175), .Y(n_498) );
INVx1_ASAP7_75t_L g507 ( .A(n_79), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_80), .A2(n_468), .B(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g784 ( .A1(n_81), .A2(n_785), .B1(n_786), .B2(n_789), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_81), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_82), .A2(n_468), .B(n_473), .C(n_478), .Y(n_467) );
INVx1_ASAP7_75t_L g115 ( .A(n_83), .Y(n_115) );
AND2x2_ASAP7_75t_L g190 ( .A(n_84), .B(n_175), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_85), .B(n_152), .Y(n_224) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_86), .B(n_175), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_87), .A2(n_468), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_88), .A2(n_128), .B1(n_438), .B2(n_439), .Y(n_127) );
INVx1_ASAP7_75t_L g438 ( .A(n_88), .Y(n_438) );
AND2x2_ASAP7_75t_L g234 ( .A(n_89), .B(n_215), .Y(n_234) );
AND2x2_ASAP7_75t_L g178 ( .A(n_91), .B(n_175), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_92), .B(n_161), .Y(n_223) );
INVx1_ASAP7_75t_L g484 ( .A(n_93), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_94), .B(n_163), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_95), .B(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_96), .A2(n_146), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g531 ( .A(n_97), .B(n_175), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_98), .B(n_163), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_99), .A2(n_552), .B(n_553), .C(n_555), .Y(n_551) );
BUFx2_ASAP7_75t_SL g123 ( .A(n_100), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_101), .A2(n_146), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_102), .B(n_153), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_119), .B(n_804), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_104), .B(n_805), .Y(n_804) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_107), .B(n_116), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx3_ASAP7_75t_L g444 ( .A(n_109), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x6_ASAP7_75t_SL g780 ( .A(n_110), .B(n_111), .Y(n_780) );
AND2x6_ASAP7_75t_SL g783 ( .A(n_110), .B(n_112), .Y(n_783) );
OR2x2_ASAP7_75t_L g802 ( .A(n_110), .B(n_112), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AO21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_445), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
CKINVDCx11_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
AOI31xp33_ASAP7_75t_L g445 ( .A1(n_122), .A2(n_446), .A3(n_790), .B(n_799), .Y(n_445) );
CKINVDCx8_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_127), .B(n_440), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g439 ( .A(n_128), .Y(n_439) );
XOR2x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
INVx3_ASAP7_75t_L g781 ( .A(n_132), .Y(n_781) );
OAI22xp5_ASAP7_75t_SL g791 ( .A1(n_132), .A2(n_792), .B1(n_794), .B2(n_795), .Y(n_791) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_350), .Y(n_132) );
AND4x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_262), .C(n_289), .D(n_324), .Y(n_133) );
AOI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_187), .B1(n_227), .B2(n_242), .C(n_246), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_166), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_137), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g303 ( .A(n_138), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g358 ( .A(n_138), .B(n_313), .Y(n_358) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g261 ( .A(n_139), .B(n_179), .Y(n_261) );
AND2x4_ASAP7_75t_L g297 ( .A(n_139), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g311 ( .A(n_139), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g228 ( .A(n_140), .Y(n_228) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_140), .Y(n_400) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B(n_165), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_141), .A2(n_192), .B(n_193), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_141), .Y(n_204) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_141), .A2(n_145), .B(n_165), .Y(n_274) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x4_ASAP7_75t_L g215 ( .A(n_143), .B(n_144), .Y(n_215) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
BUFx3_ASAP7_75t_L g465 ( .A(n_147), .Y(n_465) );
AND2x6_ASAP7_75t_L g161 ( .A(n_148), .B(n_154), .Y(n_161) );
INVx2_ASAP7_75t_L g472 ( .A(n_148), .Y(n_472) );
AND2x4_ASAP7_75t_L g468 ( .A(n_149), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x4_ASAP7_75t_L g163 ( .A(n_150), .B(n_156), .Y(n_163) );
INVx2_ASAP7_75t_L g462 ( .A(n_150), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_151), .Y(n_463) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_158), .Y(n_152) );
INVx1_ASAP7_75t_L g508 ( .A(n_153), .Y(n_508) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx5_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_158), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_164), .Y(n_159) );
INVxp67_ASAP7_75t_L g511 ( .A(n_161), .Y(n_511) );
INVxp67_ASAP7_75t_L g513 ( .A(n_163), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_164), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_164), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_164), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_164), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_164), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_164), .A2(n_474), .B(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_164), .A2(n_477), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_164), .A2(n_477), .B(n_496), .C(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_164), .B(n_215), .Y(n_514) );
INVx1_ASAP7_75t_L g525 ( .A(n_164), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_164), .A2(n_477), .B(n_537), .C(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g545 ( .A1(n_164), .A2(n_477), .B(n_546), .C(n_547), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_SL g255 ( .A1(n_166), .A2(n_228), .B(n_256), .C(n_260), .Y(n_255) );
AND2x2_ASAP7_75t_L g276 ( .A(n_166), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_166), .B(n_228), .Y(n_416) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
INVx2_ASAP7_75t_L g296 ( .A(n_167), .Y(n_296) );
BUFx3_ASAP7_75t_L g312 ( .A(n_167), .Y(n_312) );
INVxp67_ASAP7_75t_L g316 ( .A(n_167), .Y(n_316) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_174), .B(n_178), .Y(n_167) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_168), .A2(n_174), .B(n_178), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_173), .Y(n_168) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_174), .A2(n_180), .B(n_186), .Y(n_179) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_174), .A2(n_180), .B(n_186), .Y(n_241) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_174), .A2(n_533), .B(n_539), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_174), .A2(n_175), .B1(n_551), .B2(n_556), .Y(n_550) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_174), .A2(n_533), .B(n_539), .Y(n_569) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_176), .B(n_559), .Y(n_558) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx4f_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
INVx2_ASAP7_75t_L g295 ( .A(n_179), .Y(n_295) );
AND2x2_ASAP7_75t_L g301 ( .A(n_179), .B(n_274), .Y(n_301) );
AND2x2_ASAP7_75t_L g327 ( .A(n_179), .B(n_296), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_181), .B(n_185), .Y(n_180) );
AOI211xp5_ASAP7_75t_L g324 ( .A1(n_187), .A2(n_325), .B(n_328), .C(n_338), .Y(n_324) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_188), .B(n_206), .Y(n_187) );
OAI321xp33_ASAP7_75t_L g299 ( .A1(n_188), .A2(n_247), .A3(n_300), .B1(n_302), .B2(n_303), .C(n_305), .Y(n_299) );
AND2x2_ASAP7_75t_L g420 ( .A(n_188), .B(n_395), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_188), .Y(n_423) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_197), .Y(n_188) );
INVx5_ASAP7_75t_L g245 ( .A(n_189), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_189), .B(n_259), .Y(n_258) );
NOR2x1_ASAP7_75t_SL g290 ( .A(n_189), .B(n_291), .Y(n_290) );
BUFx2_ASAP7_75t_L g335 ( .A(n_189), .Y(n_335) );
AND2x2_ASAP7_75t_L g437 ( .A(n_189), .B(n_207), .Y(n_437) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
AND2x2_ASAP7_75t_L g244 ( .A(n_197), .B(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_197), .Y(n_254) );
INVx4_ASAP7_75t_L g259 ( .A(n_197), .Y(n_259) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_204), .B(n_205), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_203), .Y(n_198) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_204), .A2(n_492), .B(n_498), .Y(n_491) );
INVx1_ASAP7_75t_L g302 ( .A(n_206), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_R g405 ( .A1(n_206), .A2(n_244), .B(n_276), .C(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g425 ( .A(n_206), .B(n_250), .Y(n_425) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
INVx1_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
INVx2_ASAP7_75t_L g249 ( .A(n_207), .Y(n_249) );
OR2x2_ASAP7_75t_L g268 ( .A(n_207), .B(n_259), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_207), .B(n_291), .Y(n_337) );
BUFx3_ASAP7_75t_L g344 ( .A(n_207), .Y(n_344) );
INVx2_ASAP7_75t_SL g478 ( .A(n_208), .Y(n_478) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_208), .A2(n_544), .B(n_548), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_215), .Y(n_209) );
INVx1_ASAP7_75t_SL g218 ( .A(n_215), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_215), .B(n_240), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_215), .A2(n_482), .B(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g307 ( .A(n_216), .Y(n_307) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_216), .Y(n_320) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g253 ( .A(n_217), .Y(n_253) );
INVx1_ASAP7_75t_L g362 ( .A(n_217), .Y(n_362) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_218), .B(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
AND2x2_ASAP7_75t_L g263 ( .A(n_227), .B(n_264), .Y(n_263) );
OAI31xp33_ASAP7_75t_L g414 ( .A1(n_227), .A2(n_415), .A3(n_417), .B(n_420), .Y(n_414) );
INVx1_ASAP7_75t_SL g432 ( .A(n_227), .Y(n_432) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AOI21xp33_ASAP7_75t_L g246 ( .A1(n_228), .A2(n_247), .B(n_255), .Y(n_246) );
NAND2x1_ASAP7_75t_L g326 ( .A(n_228), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g355 ( .A(n_228), .Y(n_355) );
INVx2_ASAP7_75t_L g304 ( .A(n_229), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_229), .B(n_287), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_229), .B(n_286), .Y(n_396) );
NOR2xp33_ASAP7_75t_SL g404 ( .A(n_229), .B(n_355), .Y(n_404) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_241), .Y(n_229) );
AND2x2_ASAP7_75t_SL g273 ( .A(n_230), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g284 ( .A(n_230), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g313 ( .A(n_230), .B(n_295), .Y(n_313) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
BUFx2_ASAP7_75t_L g277 ( .A(n_231), .Y(n_277) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g298 ( .A(n_232), .Y(n_298) );
OAI21x1_ASAP7_75t_SL g232 ( .A1(n_233), .A2(n_235), .B(n_239), .Y(n_232) );
INVx1_ASAP7_75t_L g240 ( .A(n_234), .Y(n_240) );
INVx2_ASAP7_75t_L g285 ( .A(n_241), .Y(n_285) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_241), .Y(n_345) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g281 ( .A(n_243), .Y(n_281) );
AND2x2_ASAP7_75t_L g360 ( .A(n_243), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g271 ( .A(n_244), .B(n_265), .Y(n_271) );
INVx2_ASAP7_75t_SL g319 ( .A(n_244), .Y(n_319) );
INVx4_ASAP7_75t_L g250 ( .A(n_245), .Y(n_250) );
AND2x2_ASAP7_75t_L g348 ( .A(n_245), .B(n_291), .Y(n_348) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_245), .B(n_361), .Y(n_366) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_245), .B(n_259), .Y(n_383) );
INVx1_ASAP7_75t_L g389 ( .A(n_247), .Y(n_389) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx1_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
OR2x2_ASAP7_75t_L g321 ( .A(n_248), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
OR2x2_ASAP7_75t_L g373 ( .A(n_249), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g403 ( .A(n_249), .B(n_291), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_250), .B(n_253), .Y(n_279) );
AND2x2_ASAP7_75t_L g371 ( .A(n_250), .B(n_361), .Y(n_371) );
AND2x4_ASAP7_75t_L g433 ( .A(n_250), .B(n_312), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx2_ASAP7_75t_L g257 ( .A(n_252), .Y(n_257) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp67_ASAP7_75t_SL g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OAI322xp33_ASAP7_75t_SL g269 ( .A1(n_257), .A2(n_270), .A3(n_272), .B1(n_275), .B2(n_278), .C1(n_280), .C2(n_282), .Y(n_269) );
INVx1_ASAP7_75t_L g427 ( .A(n_257), .Y(n_427) );
OR2x2_ASAP7_75t_L g280 ( .A(n_258), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g306 ( .A(n_259), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_259), .B(n_307), .Y(n_322) );
INVx2_ASAP7_75t_L g349 ( .A(n_259), .Y(n_349) );
AND2x4_ASAP7_75t_L g361 ( .A(n_259), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_261), .B(n_277), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B(n_269), .Y(n_262) );
AND2x2_ASAP7_75t_L g330 ( .A(n_264), .B(n_297), .Y(n_330) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_265), .B(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_266), .B(n_285), .Y(n_370) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g278 ( .A(n_268), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_271), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g406 ( .A(n_273), .B(n_370), .Y(n_406) );
NOR4xp25_ASAP7_75t_L g410 ( .A(n_273), .B(n_287), .C(n_327), .D(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g287 ( .A(n_274), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g323 ( .A(n_274), .B(n_298), .Y(n_323) );
AND2x4_ASAP7_75t_L g387 ( .A(n_274), .B(n_298), .Y(n_387) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_277), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
OR2x2_ASAP7_75t_L g376 ( .A(n_284), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g430 ( .A(n_284), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_285), .B(n_297), .Y(n_331) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AOI211xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_292), .B(n_299), .C(n_314), .Y(n_289) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_295), .B(n_298), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_296), .B(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g378 ( .A(n_296), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_297), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g393 ( .A(n_297), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B(n_309), .Y(n_305) );
AND2x4_ASAP7_75t_L g342 ( .A(n_306), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g436 ( .A(n_306), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_SL g340 ( .A(n_312), .Y(n_340) );
AND2x2_ASAP7_75t_L g399 ( .A(n_313), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g413 ( .A(n_313), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_317), .B(n_321), .C(n_323), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_315), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g391 ( .A(n_316), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g412 ( .A(n_316), .B(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OR2x2_ASAP7_75t_L g401 ( .A(n_319), .B(n_343), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_322), .A2(n_329), .B1(n_331), .B2(n_332), .Y(n_328) );
INVx1_ASAP7_75t_SL g419 ( .A(n_323), .Y(n_419) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_334), .B(n_343), .Y(n_385) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_337), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B1(n_345), .B2(n_346), .Y(n_338) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI21xp5_ASAP7_75t_SL g352 ( .A1(n_343), .A2(n_353), .B(n_356), .Y(n_352) );
AND2x2_ASAP7_75t_L g381 ( .A(n_343), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND3x2_ASAP7_75t_L g347 ( .A(n_344), .B(n_348), .C(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g409 ( .A(n_344), .B(n_366), .Y(n_409) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g394 ( .A(n_349), .B(n_395), .Y(n_394) );
NOR2xp67_ASAP7_75t_L g350 ( .A(n_351), .B(n_407), .Y(n_350) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_367), .C(n_388), .D(n_405), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B1(n_363), .B2(n_365), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_359), .A2(n_373), .B1(n_393), .B2(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g374 ( .A(n_361), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_363), .A2(n_386), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_372), .B2(n_375), .C(n_379), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_384), .B1(n_385), .B2(n_386), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_382), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_382), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_394), .B2(n_396), .C(n_397), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_391), .B(n_393), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .B1(n_402), .B2(n_404), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI211xp5_ASAP7_75t_SL g422 ( .A1(n_403), .A2(n_423), .B(n_424), .C(n_426), .Y(n_422) );
OAI211xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_414), .C(n_421), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_428), .B1(n_431), .B2(n_433), .C(n_434), .Y(n_421) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g803 ( .A(n_440), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
CKINVDCx11_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_447), .B(n_784), .Y(n_446) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVxp67_ASAP7_75t_L g794 ( .A(n_450), .Y(n_794) );
NAND4xp75_ASAP7_75t_L g450 ( .A(n_451), .B(n_631), .C(n_697), .D(n_760), .Y(n_450) );
NOR2x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_594), .Y(n_451) );
OR3x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_564), .C(n_591), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_499), .B(n_520), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_488), .Y(n_455) );
AND2x2_ASAP7_75t_L g694 ( .A(n_456), .B(n_664), .Y(n_694) );
INVx1_ASAP7_75t_L g767 ( .A(n_456), .Y(n_767) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_479), .Y(n_456) );
INVx2_ASAP7_75t_L g519 ( .A(n_457), .Y(n_519) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_457), .Y(n_582) );
AND2x2_ASAP7_75t_L g586 ( .A(n_457), .B(n_502), .Y(n_586) );
AND2x4_ASAP7_75t_L g602 ( .A(n_457), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g606 ( .A(n_457), .Y(n_606) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_467), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .C(n_466), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g487 ( .A(n_461), .B(n_465), .Y(n_487) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
OR2x6_ASAP7_75t_L g477 ( .A(n_462), .B(n_472), .Y(n_477) );
INVxp33_ASAP7_75t_L g528 ( .A(n_462), .Y(n_528) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVxp67_ASAP7_75t_L g561 ( .A(n_468), .Y(n_561) );
NOR2x1p5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g529 ( .A(n_471), .Y(n_529) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_477), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_505) );
INVxp67_ASAP7_75t_L g552 ( .A(n_477), .Y(n_552) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_478), .A2(n_523), .B(n_531), .Y(n_522) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_478), .A2(n_523), .B(n_531), .Y(n_570) );
AND2x2_ASAP7_75t_L g500 ( .A(n_479), .B(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g583 ( .A(n_479), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_479), .B(n_573), .Y(n_587) );
INVx2_ASAP7_75t_L g601 ( .A(n_479), .Y(n_601) );
AND2x4_ASAP7_75t_L g605 ( .A(n_479), .B(n_606), .Y(n_605) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_479), .Y(n_640) );
OR2x2_ASAP7_75t_L g646 ( .A(n_479), .B(n_491), .Y(n_646) );
NOR2x1_ASAP7_75t_SL g675 ( .A(n_479), .B(n_502), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_479), .B(n_749), .Y(n_777) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g563 ( .A(n_487), .Y(n_563) );
AND2x2_ASAP7_75t_L g674 ( .A(n_488), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2x1_ASAP7_75t_L g708 ( .A(n_489), .B(n_501), .Y(n_708) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g516 ( .A(n_491), .Y(n_516) );
INVx2_ASAP7_75t_L g574 ( .A(n_491), .Y(n_574) );
AND2x2_ASAP7_75t_L g597 ( .A(n_491), .B(n_502), .Y(n_597) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_491), .Y(n_624) );
INVx1_ASAP7_75t_L g665 ( .A(n_491), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_515), .Y(n_499) );
AND2x2_ASAP7_75t_L g677 ( .A(n_500), .B(n_572), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_501), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g744 ( .A(n_501), .Y(n_744) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g603 ( .A(n_502), .Y(n_603) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_509), .B(n_514), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_508), .B(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_509) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_515), .A2(n_681), .B(n_685), .C(n_691), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_516), .B(n_517), .Y(n_515) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_517), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_SL g727 ( .A(n_517), .Y(n_727) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g649 ( .A(n_519), .B(n_603), .Y(n_649) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_540), .Y(n_520) );
AOI32xp33_ASAP7_75t_L g685 ( .A1(n_521), .A2(n_669), .A3(n_686), .B1(n_687), .B2(n_689), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_532), .Y(n_521) );
INVx2_ASAP7_75t_L g611 ( .A(n_522), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_522), .B(n_543), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_524), .B(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g623 ( .A(n_532), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_532), .B(n_549), .Y(n_654) );
AND2x2_ASAP7_75t_L g659 ( .A(n_532), .B(n_660), .Y(n_659) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_532), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
OR2x2_ASAP7_75t_L g642 ( .A(n_540), .B(n_643), .Y(n_642) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g593 ( .A(n_541), .B(n_567), .Y(n_593) );
AND2x2_ASAP7_75t_L g742 ( .A(n_541), .B(n_740), .Y(n_742) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g579 ( .A(n_543), .Y(n_579) );
AND2x4_ASAP7_75t_L g618 ( .A(n_543), .B(n_619), .Y(n_618) );
INVxp67_ASAP7_75t_L g652 ( .A(n_543), .Y(n_652) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_543), .Y(n_660) );
AND2x2_ASAP7_75t_L g669 ( .A(n_543), .B(n_549), .Y(n_669) );
INVx1_ASAP7_75t_L g753 ( .A(n_543), .Y(n_753) );
INVx2_ASAP7_75t_L g590 ( .A(n_549), .Y(n_590) );
INVx1_ASAP7_75t_L g617 ( .A(n_549), .Y(n_617) );
INVx1_ASAP7_75t_L g684 ( .A(n_549), .Y(n_684) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_557), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI32xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_575), .A3(n_580), .B1(n_584), .B2(n_588), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_566), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_567), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g668 ( .A(n_567), .B(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g693 ( .A(n_567), .Y(n_693) );
AND2x2_ASAP7_75t_L g774 ( .A(n_567), .B(n_616), .Y(n_774) );
AND2x4_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g589 ( .A(n_569), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g688 ( .A(n_569), .B(n_611), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_569), .B(n_590), .Y(n_710) );
NOR2x1_ASAP7_75t_L g752 ( .A(n_569), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g619 ( .A(n_570), .Y(n_619) );
INVx1_ASAP7_75t_L g643 ( .A(n_570), .Y(n_643) );
AND2x2_ASAP7_75t_L g658 ( .A(n_570), .B(n_590), .Y(n_658) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g686 ( .A(n_572), .B(n_675), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_572), .B(n_605), .Y(n_756) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_573), .Y(n_725) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_574), .Y(n_707) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g608 ( .A(n_577), .B(n_609), .Y(n_608) );
NOR2xp67_ASAP7_75t_L g692 ( .A(n_577), .B(n_693), .Y(n_692) );
NOR2xp67_ASAP7_75t_SL g779 ( .A(n_577), .B(n_717), .Y(n_779) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g636 ( .A(n_579), .B(n_590), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_580), .B(n_646), .Y(n_704) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_SL g670 ( .A(n_581), .B(n_597), .Y(n_670) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_583), .B(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g735 ( .A(n_583), .B(n_606), .Y(n_735) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_583), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_584), .B(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
OR2x2_ASAP7_75t_L g706 ( .A(n_585), .B(n_707), .Y(n_706) );
NOR2x1_ASAP7_75t_L g771 ( .A(n_585), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g695 ( .A(n_586), .B(n_640), .Y(n_695) );
INVxp33_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_589), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g769 ( .A(n_589), .B(n_651), .Y(n_769) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_612), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B(n_607), .Y(n_595) );
AND2x2_ASAP7_75t_L g730 ( .A(n_597), .B(n_605), .Y(n_730) );
NAND2xp33_ASAP7_75t_R g598 ( .A(n_599), .B(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g772 ( .A(n_601), .Y(n_772) );
INVx4_ASAP7_75t_L g630 ( .A(n_602), .Y(n_630) );
INVx1_ASAP7_75t_L g749 ( .A(n_603), .Y(n_749) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g743 ( .A(n_605), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_SL g747 ( .A(n_605), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_608), .A2(n_673), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g637 ( .A(n_611), .B(n_623), .Y(n_637) );
AND2x2_ASAP7_75t_L g651 ( .A(n_611), .B(n_652), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_620), .B(n_625), .C(n_628), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g699 ( .A(n_615), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g627 ( .A(n_616), .Y(n_627) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g687 ( .A(n_617), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g696 ( .A(n_617), .B(n_618), .Y(n_696) );
INVx1_ASAP7_75t_L g728 ( .A(n_617), .Y(n_728) );
AND2x4_ASAP7_75t_L g709 ( .A(n_618), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g731 ( .A(n_618), .B(n_622), .Y(n_731) );
AND2x2_ASAP7_75t_L g739 ( .A(n_618), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g714 ( .A(n_622), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_622), .B(n_636), .Y(n_716) );
AND2x2_ASAP7_75t_L g719 ( .A(n_622), .B(n_669), .Y(n_719) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_623), .B(n_684), .Y(n_733) );
AND2x2_ASAP7_75t_L g661 ( .A(n_624), .B(n_649), .Y(n_661) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g757 ( .A(n_627), .B(n_637), .Y(n_757) );
BUFx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_629), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g641 ( .A(n_630), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_630), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_671), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_655), .Y(n_632) );
OAI222xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_638), .B1(n_642), .B2(n_644), .C1(n_647), .C2(n_650), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_SL g648 ( .A(n_640), .B(n_649), .Y(n_648) );
OR2x6_ASAP7_75t_L g720 ( .A(n_640), .B(n_690), .Y(n_720) );
NAND5xp2_ASAP7_75t_L g723 ( .A(n_640), .B(n_643), .C(n_659), .D(n_724), .E(n_726), .Y(n_723) );
NAND2x1_ASAP7_75t_L g759 ( .A(n_641), .B(n_645), .Y(n_759) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_646), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_648), .A2(n_739), .B1(n_742), .B2(n_743), .Y(n_738) );
INVx2_ASAP7_75t_L g690 ( .A(n_649), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_649), .B(n_665), .Y(n_702) );
INVx3_ASAP7_75t_L g737 ( .A(n_650), .Y(n_737) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
AND2x2_ASAP7_75t_L g682 ( .A(n_651), .B(n_683), .Y(n_682) );
BUFx2_ASAP7_75t_L g715 ( .A(n_651), .Y(n_715) );
INVx2_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g678 ( .A(n_654), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_656), .B(n_667), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_661), .B(n_662), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g666 ( .A(n_658), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_661), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_SL g748 ( .A(n_665), .B(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_680), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_676), .B(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g717 ( .A(n_688), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_691) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_721), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_703), .C(n_711), .Y(n_698) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OA21x2_ASAP7_75t_SL g703 ( .A1(n_704), .A2(n_705), .B(n_709), .Y(n_703) );
NAND2xp33_ASAP7_75t_SL g705 ( .A(n_706), .B(n_708), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_718), .B(n_720), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_716), .C(n_717), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_715), .A2(n_755), .B1(n_757), .B2(n_758), .Y(n_754) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_745), .Y(n_721) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_723), .B(n_729), .C(n_736), .D(n_738), .Y(n_722) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g734 ( .A(n_725), .B(n_735), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g765 ( .A(n_728), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_732), .B2(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_734), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_750), .B(n_754), .Y(n_745) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_775), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_765), .B(n_766), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_770), .B2(n_773), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
CKINVDCx11_ASAP7_75t_R g793 ( .A(n_780), .Y(n_793) );
CKINVDCx11_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_783), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_784), .Y(n_798) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_791), .B(n_798), .Y(n_790) );
INVx1_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
INVx4_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
INVx3_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_803), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
endmodule