module fake_jpeg_3175_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_61),
.B(n_67),
.Y(n_154)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_66),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_0),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_68),
.Y(n_212)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_20),
.B(n_2),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_70),
.B(n_73),
.Y(n_157)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_74),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_21),
.B(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_75),
.B(n_111),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_30),
.B(n_11),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_78),
.B(n_83),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_34),
.B(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_84),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_34),
.B(n_11),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_107),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_96),
.B(n_123),
.Y(n_184)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_100),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

NAND2x1_ASAP7_75t_SL g210 ( 
.A(n_101),
.B(n_102),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_113),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_108),
.B(n_109),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

CKINVDCx6p67_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_17),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_116),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_46),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_118),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_119),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_51),
.Y(n_153)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_121),
.B(n_124),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_52),
.B(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_26),
.B(n_2),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_26),
.B(n_50),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_125),
.B(n_146),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_51),
.B1(n_38),
.B2(n_24),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_126),
.A2(n_203),
.A3(n_171),
.B1(n_160),
.B2(n_130),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_67),
.A2(n_35),
.B1(n_37),
.B2(n_50),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_128),
.A2(n_137),
.B1(n_144),
.B2(n_147),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_70),
.A2(n_28),
.B1(n_35),
.B2(n_37),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_51),
.B1(n_28),
.B2(n_40),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_90),
.A2(n_24),
.B1(n_36),
.B2(n_39),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_153),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_75),
.A2(n_40),
.B1(n_49),
.B2(n_42),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_156),
.A2(n_180),
.B1(n_155),
.B2(n_143),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_49),
.B(n_42),
.C(n_31),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_158),
.A2(n_134),
.B(n_167),
.C(n_184),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_95),
.A2(n_39),
.B1(n_36),
.B2(n_31),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_161),
.A2(n_168),
.B1(n_196),
.B2(n_176),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_57),
.B(n_53),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_163),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_83),
.B(n_15),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_164),
.B(n_174),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_106),
.A2(n_33),
.B1(n_53),
.B2(n_4),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_101),
.A2(n_53),
.B1(n_33),
.B2(n_48),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_170),
.A2(n_178),
.B1(n_204),
.B2(n_209),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_63),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_102),
.A2(n_53),
.B1(n_48),
.B2(n_4),
.Y(n_178)
);

CKINVDCx12_ASAP7_75t_R g179 ( 
.A(n_122),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_65),
.A2(n_53),
.B1(n_3),
.B2(n_5),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_66),
.B(n_12),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_186),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_74),
.A2(n_53),
.B(n_15),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_79),
.B(n_16),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_187),
.B(n_188),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_85),
.B(n_17),
.C(n_3),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_88),
.B(n_2),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_191),
.B(n_199),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_89),
.B(n_3),
.C(n_5),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_210),
.C(n_196),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_103),
.A2(n_5),
.B1(n_7),
.B2(n_108),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_109),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_114),
.B(n_7),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_213),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_116),
.A2(n_7),
.B1(n_67),
.B2(n_124),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_7),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_205),
.B(n_207),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_67),
.A2(n_124),
.B1(n_70),
.B2(n_75),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_93),
.B(n_123),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_163),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_215),
.B(n_250),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_154),
.B(n_157),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_216),
.B(n_234),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_218),
.Y(n_310)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_220),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_144),
.A2(n_169),
.B1(n_178),
.B2(n_170),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_221),
.A2(n_276),
.B1(n_214),
.B2(n_277),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_149),
.B1(n_150),
.B2(n_129),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_149),
.A2(n_150),
.B1(n_131),
.B2(n_172),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_226),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_149),
.A2(n_172),
.B1(n_159),
.B2(n_132),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_227),
.A2(n_236),
.B1(n_240),
.B2(n_241),
.Y(n_301)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_230),
.B(n_235),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_232),
.B(n_251),
.Y(n_293)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_138),
.Y(n_233)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_158),
.B(n_148),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_165),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_132),
.A2(n_159),
.B1(n_142),
.B2(n_141),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_152),
.Y(n_239)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_126),
.B1(n_147),
.B2(n_197),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_142),
.A2(n_126),
.B1(n_173),
.B2(n_136),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_136),
.A2(n_208),
.B1(n_145),
.B2(n_195),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_243),
.A2(n_246),
.B1(n_247),
.B2(n_253),
.Y(n_324)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_208),
.A2(n_195),
.B1(n_198),
.B2(n_175),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_175),
.A2(n_200),
.B1(n_203),
.B2(n_168),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_249),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_139),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_252),
.B(n_262),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_140),
.B(n_177),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_151),
.B(n_135),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_255),
.B(n_282),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_155),
.A2(n_139),
.B1(n_143),
.B2(n_161),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_256),
.B(n_258),
.Y(n_317)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_203),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_259),
.B(n_260),
.Y(n_334)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_189),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_263),
.B(n_279),
.Y(n_319)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_266),
.Y(n_314)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_127),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_268),
.Y(n_316)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_166),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_130),
.A2(n_194),
.B1(n_133),
.B2(n_166),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_269),
.A2(n_275),
.B1(n_256),
.B2(n_218),
.Y(n_330)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_270),
.B(n_272),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_181),
.A2(n_192),
.B1(n_211),
.B2(n_133),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_271),
.A2(n_288),
.B1(n_267),
.B2(n_272),
.Y(n_323)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_274),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_162),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_162),
.A2(n_180),
.B1(n_156),
.B2(n_120),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_162),
.A2(n_204),
.B1(n_209),
.B2(n_185),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_185),
.B(n_67),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_277),
.B(n_238),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_154),
.B(n_185),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_190),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_190),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_280),
.B(n_286),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_154),
.B(n_185),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_231),
.Y(n_309)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_165),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_285),
.Y(n_297)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_201),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_190),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_204),
.A2(n_180),
.B1(n_209),
.B2(n_185),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_249),
.B(n_234),
.C(n_259),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_289),
.A2(n_335),
.B(n_317),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_290),
.A2(n_323),
.B1(n_322),
.B2(n_306),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_221),
.A2(n_214),
.B1(n_288),
.B2(n_253),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_291),
.A2(n_296),
.B1(n_298),
.B2(n_271),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_261),
.B1(n_215),
.B2(n_250),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_215),
.A2(n_248),
.B1(n_278),
.B2(n_283),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_303),
.B(n_309),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_216),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_307),
.B(n_308),
.C(n_298),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_224),
.B(n_244),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_225),
.A2(n_252),
.B(n_281),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_315),
.A2(n_333),
.B(n_325),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_239),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_331),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_264),
.B(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_321),
.B(n_302),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_233),
.B(n_286),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_219),
.B(n_262),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_332),
.B(n_316),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_258),
.A2(n_217),
.B(n_235),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_258),
.A2(n_230),
.B(n_228),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_280),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_340),
.B(n_361),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_341),
.B(n_344),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_292),
.B(n_229),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_342),
.B(n_345),
.Y(n_406)
);

OAI31xp33_ASAP7_75t_SL g343 ( 
.A1(n_289),
.A2(n_296),
.A3(n_290),
.B(n_315),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_370),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_287),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_292),
.B(n_260),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_291),
.A2(n_237),
.B1(n_268),
.B2(n_270),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_355),
.Y(n_378)
);

INVx11_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_309),
.B(n_265),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_350),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_274),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_319),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_357),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_334),
.A2(n_266),
.B1(n_273),
.B2(n_257),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_242),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_336),
.C(n_333),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_285),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_364),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_302),
.A2(n_338),
.B1(n_326),
.B2(n_334),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_369),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_338),
.A2(n_301),
.B1(n_329),
.B2(n_324),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_363),
.A2(n_376),
.B(n_377),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_308),
.B(n_312),
.Y(n_364)
);

BUFx12f_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_366),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_312),
.B(n_313),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_373),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_306),
.B1(n_317),
.B2(n_318),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_335),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_371),
.B(n_300),
.Y(n_398)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_293),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_375),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_306),
.A2(n_317),
.B1(n_323),
.B2(n_322),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_402),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_387),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_371),
.A2(n_329),
.B1(n_320),
.B2(n_327),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_398),
.B1(n_355),
.B2(n_375),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_344),
.Y(n_387)
);

OA22x2_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_337),
.B1(n_300),
.B2(n_304),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_390),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_374),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_342),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_400),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_377),
.A2(n_328),
.B(n_297),
.C(n_314),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_394),
.B(n_370),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_313),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_399),
.B(n_294),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_349),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_294),
.C(n_299),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_407),
.B(n_356),
.C(n_369),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_383),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_414),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_411),
.C(n_425),
.Y(n_448)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_412),
.Y(n_438)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_384),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_408),
.Y(n_416)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_384),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_420),
.B(n_421),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_397),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_422),
.A2(n_437),
.B1(n_400),
.B2(n_393),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_397),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_423),
.Y(n_458)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_429),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_340),
.C(n_376),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_343),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_430),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_345),
.C(n_354),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_431),
.C(n_433),
.Y(n_459)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_401),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_354),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_339),
.C(n_351),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_434),
.B1(n_406),
.B2(n_423),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_341),
.C(n_360),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_391),
.A2(n_352),
.B1(n_353),
.B2(n_348),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_403),
.Y(n_435)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_435),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_390),
.B(n_365),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_436),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_405),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_440),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_405),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_379),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_454),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_392),
.B(n_391),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_449),
.A2(n_427),
.B1(n_415),
.B2(n_398),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_416),
.A2(n_408),
.B(n_394),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_457),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_392),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_392),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_461),
.C(n_433),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_382),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_415),
.A2(n_398),
.B(n_387),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_462),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_472),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_430),
.C(n_386),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_465),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_386),
.C(n_382),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_449),
.B1(n_438),
.B2(n_450),
.Y(n_489)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_455),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_445),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_470),
.Y(n_483)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_452),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_462),
.A2(n_422),
.B1(n_417),
.B2(n_434),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_471),
.A2(n_476),
.B1(n_466),
.B2(n_472),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_385),
.C(n_435),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_452),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_347),
.B1(n_451),
.B2(n_403),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_458),
.A2(n_395),
.B1(n_381),
.B2(n_378),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_429),
.C(n_424),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_439),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_441),
.B(n_406),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_479),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_480),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_495),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_SL g486 ( 
.A(n_481),
.B(n_460),
.C(n_447),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_486),
.B(n_440),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_478),
.A2(n_449),
.B(n_444),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_488),
.A2(n_494),
.B(n_463),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_388),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_471),
.A2(n_451),
.B1(n_456),
.B2(n_443),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_492),
.B1(n_493),
.B2(n_419),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_476),
.A2(n_456),
.B(n_459),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_464),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_503),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_477),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_499),
.B(n_508),
.Y(n_517)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_483),
.Y(n_500)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_500),
.Y(n_514)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_485),
.Y(n_501)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_504),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_488),
.A2(n_465),
.B(n_475),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_489),
.A2(n_475),
.B(n_461),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_506),
.B1(n_494),
.B2(n_491),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_486),
.B1(n_496),
.B2(n_482),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_474),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_498),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_505),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_516),
.Y(n_523)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_511),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_495),
.C(n_490),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_516),
.B(n_497),
.C(n_503),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_518),
.B(n_522),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_517),
.B(n_504),
.Y(n_520)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_520),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_512),
.Y(n_525)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_523),
.A2(n_515),
.B(n_511),
.Y(n_524)
);

AOI21xp33_ASAP7_75t_L g529 ( 
.A1(n_524),
.A2(n_519),
.B(n_513),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_525),
.A2(n_514),
.B(n_520),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_528),
.A2(n_529),
.B(n_527),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_531),
.C(n_526),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_528),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_532),
.B(n_513),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_533),
.B(n_474),
.Y(n_534)
);


endmodule