module fake_jpeg_21895_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_0),
.CON(n_39),
.SN(n_39)
);

AO22x1_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_47),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_52),
.B1(n_22),
.B2(n_17),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_27),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_23),
.B(n_22),
.C(n_17),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_51),
.A2(n_21),
.B1(n_28),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_60),
.B1(n_64),
.B2(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_38),
.C(n_36),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_5),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_67),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_81),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_37),
.B1(n_33),
.B2(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_78),
.B1(n_82),
.B2(n_67),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_42),
.B(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_1),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_6),
.Y(n_104)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_22),
.B1(n_17),
.B2(n_16),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_49),
.Y(n_83)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_86),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_90),
.B1(n_95),
.B2(n_84),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_22),
.B1(n_17),
.B2(n_16),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_75),
.B1(n_59),
.B2(n_83),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_110),
.C(n_95),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_75),
.B(n_86),
.Y(n_114)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_73),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_6),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_115),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_65),
.B1(n_61),
.B2(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_119),
.B1(n_126),
.B2(n_134),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_117),
.B(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_123),
.B1(n_97),
.B2(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_74),
.B(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_83),
.B1(n_77),
.B2(n_71),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_79),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_7),
.B(n_8),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_133),
.B(n_135),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_7),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_90),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_7),
.B(n_8),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_56),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_120),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_148),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_150),
.C(n_155),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_97),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_149),
.B(n_115),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_93),
.B(n_111),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_93),
.C(n_92),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_92),
.C(n_99),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_103),
.C(n_104),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_128),
.C(n_113),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_174),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_173),
.B(n_177),
.Y(n_181)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_116),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_132),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_175),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_126),
.C(n_125),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_147),
.B1(n_154),
.B2(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_130),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_141),
.B1(n_152),
.B2(n_139),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_179),
.B1(n_167),
.B2(n_166),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_134),
.B1(n_145),
.B2(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_140),
.B1(n_145),
.B2(n_143),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_171),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_140),
.B1(n_143),
.B2(n_138),
.Y(n_187)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_147),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_161),
.C(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_197),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_161),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_195),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_180),
.B1(n_167),
.B2(n_189),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_160),
.B(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_196),
.B(n_200),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_155),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_187),
.C(n_185),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_166),
.C(n_150),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_202),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_188),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_182),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_195),
.B1(n_197),
.B2(n_192),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_198),
.A2(n_189),
.B1(n_172),
.B2(n_158),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_144),
.B1(n_153),
.B2(n_111),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_SL g215 ( 
.A(n_212),
.B(n_193),
.Y(n_215)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_211),
.B(n_153),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_217),
.B(n_216),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_135),
.B(n_107),
.Y(n_219)
);

OAI321xp33_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_209),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.C(n_218),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_222),
.C(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_204),
.C(n_210),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_222),
.C(n_227),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_230),
.A2(n_231),
.B(n_10),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_11),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_14),
.Y(n_234)
);


endmodule