module fake_ibex_1997_n_4949 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_961, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_960, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4949);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_960;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4949;

wire n_4557;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_962;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_3208;
wire n_4569;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_2253;
wire n_4479;
wire n_3858;
wire n_4173;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_3060;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_3293;
wire n_2550;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_4757;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3529;
wire n_3222;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_1471;
wire n_3441;
wire n_4559;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_4851;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_1127;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_2422;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_2223;
wire n_3876;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_3096;
wire n_1278;
wire n_2059;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_985;
wire n_4611;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_4895;
wire n_3354;
wire n_4069;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_2574;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_4686;
wire n_4682;
wire n_2914;
wire n_1833;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_4733;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_4412;
wire n_4266;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_3857;
wire n_2357;
wire n_4354;
wire n_2937;
wire n_3728;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_4539;
wire n_1205;
wire n_2969;
wire n_3550;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_3502;
wire n_3935;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_4926;
wire n_4688;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_3484;
wire n_2485;
wire n_4477;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_3726;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_4491;
wire n_4672;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_4433;
wire n_3030;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4393;
wire n_3777;
wire n_4553;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_3633;
wire n_1731;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3788;
wire n_3448;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_2829;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_965;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_3787;
wire n_3445;
wire n_2080;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_2142;
wire n_3703;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_1729;
wire n_998;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_4579;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_4636;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_2442;
wire n_1067;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_1662;
wire n_3443;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_1660;
wire n_4000;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_3712;
wire n_2143;
wire n_4637;
wire n_4021;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_3327;
wire n_1114;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_1885;
wire n_1989;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_1175;
wire n_4408;
wire n_1221;
wire n_3875;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_4565;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_4574;
wire n_4242;
wire n_4748;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_4562;
wire n_1584;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_4196;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_3036;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_3332;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_1442;
wire n_2168;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_3861;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_1640;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_4590;
wire n_4602;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_1743;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_4159;
wire n_4372;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_3819;
wire n_3334;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_963;
wire n_2139;
wire n_3693;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_3641;
wire n_4887;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_3722;
wire n_3802;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_4806;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_1269;
wire n_2773;
wire n_3097;
wire n_2906;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_2859;
wire n_2564;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_2114;
wire n_1609;
wire n_3530;
wire n_1132;
wire n_4548;
wire n_1803;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_2660;
wire n_4604;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_3282;
wire n_1003;
wire n_2708;
wire n_2748;
wire n_2224;
wire n_2233;
wire n_2499;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_1553;
wire n_3542;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_1189;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_2852;
wire n_2132;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_3785;
wire n_3525;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_2481;
wire n_4409;
wire n_1264;
wire n_2808;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_4152;
wire n_1352;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_2908;
wire n_4561;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_3328;
wire n_2763;
wire n_994;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_3028;
wire n_3228;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_2086;
wire n_4832;
wire n_3666;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2108;
wire n_2535;
wire n_2945;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_3302;
wire n_1673;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_2894;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_2315;
wire n_3623;
wire n_2157;
wire n_3446;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_1105;
wire n_2898;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_4670;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_4053;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_1693;
wire n_2081;
wire n_2993;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_3989;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_967;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_3430;
wire n_1685;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_1398;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2855;
wire n_2653;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_4088;
wire n_2136;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_2262;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_1080;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4668;
wire n_2383;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_2230;
wire n_3033;
wire n_2151;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_1606;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_2826;
wire n_2112;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_4671;
wire n_1326;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_3618;
wire n_2727;
wire n_2719;
wire n_2213;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_3847;
wire n_2203;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_2646;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_4136;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1360;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_1452;
wire n_4570;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_2819;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_4407;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_3680;
wire n_3624;
wire n_2467;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1566;
wire n_1464;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_4929;
wire n_1608;
wire n_3776;
wire n_1009;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_4427;
wire n_3505;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_2525;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4297;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_2986;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_964;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_3867;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_3588;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_2271;
wire n_2356;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_2187;
wire n_2105;
wire n_2642;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_4048;
wire n_4084;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_2849;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_4860;
wire n_4438;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_2665;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_2581;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_3454;
wire n_4143;
wire n_4410;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_1433;
wire n_1907;
wire n_3994;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_4487;
wire n_1165;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_3042;
wire n_2561;
wire n_2491;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_4811;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_1419;
wire n_4738;
wire n_980;
wire n_1193;
wire n_3557;
wire n_3380;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_4086;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_966;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_1791;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_1164;
wire n_3749;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_168),
.Y(n_962)
);

BUFx10_ASAP7_75t_L g963 ( 
.A(n_384),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_845),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_935),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_649),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_67),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_112),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_641),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_687),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_896),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_669),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_947),
.Y(n_973)
);

BUFx10_ASAP7_75t_L g974 ( 
.A(n_550),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_113),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_892),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_367),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_902),
.Y(n_978)
);

CKINVDCx16_ASAP7_75t_R g979 ( 
.A(n_606),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_918),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_919),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_827),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_939),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_884),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_258),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_208),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_682),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_125),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_87),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_902),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_374),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_837),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_85),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_94),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_393),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_847),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_482),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_890),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_750),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_231),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_501),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_931),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_512),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_271),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_474),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_220),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_655),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_341),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_614),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_44),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_589),
.Y(n_1011)
);

BUFx10_ASAP7_75t_L g1012 ( 
.A(n_546),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_26),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_392),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_946),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_408),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_424),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_867),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_627),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_60),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_823),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_822),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_810),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_666),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_904),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_925),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_208),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_525),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_857),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_389),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_836),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_516),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_656),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_599),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_740),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_882),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_820),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_399),
.Y(n_1038)
);

BUFx10_ASAP7_75t_L g1039 ( 
.A(n_99),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_417),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_241),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_816),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_917),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_524),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_51),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_518),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_587),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_844),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_937),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_109),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_928),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_428),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_933),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_829),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_858),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_701),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_253),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_358),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_493),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_371),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_839),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_511),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_850),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_412),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_403),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_940),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_929),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_394),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_49),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_211),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_601),
.Y(n_1071)
);

CKINVDCx16_ASAP7_75t_R g1072 ( 
.A(n_16),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_354),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_174),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_109),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_333),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_698),
.Y(n_1077)
);

BUFx5_ASAP7_75t_L g1078 ( 
.A(n_672),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_501),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_428),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_306),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_866),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_811),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_775),
.Y(n_1084)
);

CKINVDCx16_ASAP7_75t_R g1085 ( 
.A(n_910),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_851),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_821),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_923),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_947),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_741),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_160),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_417),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_880),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_951),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_226),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_785),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_246),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_751),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_834),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_102),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_617),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_667),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_908),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_451),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_144),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_931),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_451),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_321),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_784),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_602),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_352),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_69),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_434),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_912),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_763),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_291),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_433),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_652),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_869),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_310),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_876),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_617),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_320),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_447),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_209),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_753),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_494),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_747),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_366),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_915),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_804),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_523),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_896),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_820),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_342),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_508),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_377),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_227),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_171),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_95),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_52),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_883),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_257),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_596),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_675),
.Y(n_1145)
);

CKINVDCx14_ASAP7_75t_R g1146 ( 
.A(n_167),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_647),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_544),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_257),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_723),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_842),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_768),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_141),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_864),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_770),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_168),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_470),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_97),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_89),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_835),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_241),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_327),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_771),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_816),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_879),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_700),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_596),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_24),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_385),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_620),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_118),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_118),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_674),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_843),
.Y(n_1174)
);

BUFx10_ASAP7_75t_L g1175 ( 
.A(n_954),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_930),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_286),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_427),
.Y(n_1178)
);

CKINVDCx14_ASAP7_75t_R g1179 ( 
.A(n_741),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_746),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_846),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_386),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_916),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_403),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_749),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_133),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_944),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_20),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_848),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_815),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_585),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_65),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_926),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_236),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_887),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_699),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_956),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_814),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_824),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_873),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_844),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_42),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_907),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_945),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_856),
.Y(n_1205)
);

CKINVDCx16_ASAP7_75t_R g1206 ( 
.A(n_942),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_469),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_798),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_876),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_861),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_720),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_819),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_195),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_874),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_174),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_118),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_48),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_767),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_498),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_261),
.Y(n_1220)
);

BUFx5_ASAP7_75t_L g1221 ( 
.A(n_925),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_154),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_158),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_207),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_828),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_356),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_857),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_883),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_364),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_448),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_389),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_870),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_137),
.Y(n_1233)
);

CKINVDCx14_ASAP7_75t_R g1234 ( 
.A(n_922),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_329),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_598),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_367),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_817),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_522),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_185),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_19),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_691),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_895),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_851),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_585),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_885),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_886),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_214),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_831),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_949),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_522),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_841),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_59),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_439),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_748),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_336),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_900),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_141),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_911),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_186),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_286),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_185),
.Y(n_1262)
);

BUFx8_ASAP7_75t_SL g1263 ( 
.A(n_821),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_299),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_849),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_377),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_452),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_27),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_873),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_272),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_878),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_792),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_732),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_955),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_863),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_411),
.Y(n_1276)
);

BUFx10_ASAP7_75t_L g1277 ( 
.A(n_934),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_492),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_897),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_927),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_231),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_702),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_85),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_840),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_339),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_639),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_749),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_941),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_920),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_932),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_379),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_325),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_517),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_662),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_901),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_656),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_798),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_541),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_801),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_39),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_800),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_276),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_384),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_578),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_456),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_6),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_331),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_877),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_833),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_185),
.Y(n_1310)
);

CKINVDCx14_ASAP7_75t_R g1311 ( 
.A(n_830),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_364),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_151),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_708),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_871),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_36),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_650),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_885),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_875),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_826),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_530),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_12),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_726),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_73),
.Y(n_1324)
);

BUFx10_ASAP7_75t_L g1325 ( 
.A(n_674),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_554),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_603),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_502),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_832),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_721),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_335),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_952),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_107),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_148),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_734),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_32),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_160),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_523),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_899),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_77),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_721),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_269),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_865),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_597),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_98),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_888),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_942),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_854),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_940),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_249),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_435),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_98),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_914),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_55),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_709),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_490),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_492),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_761),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_794),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_743),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_66),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_19),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_4),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_805),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_860),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_358),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_686),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_543),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_540),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_745),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_924),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_326),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_317),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_4),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_958),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_34),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_587),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_831),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_255),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_593),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_946),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_728),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_32),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_750),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_369),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_50),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_866),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_95),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_92),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_631),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_865),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_250),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_825),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_74),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_732),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_835),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_731),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_303),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_738),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_453),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_353),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_658),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_41),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_153),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_950),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_954),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_45),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_330),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_957),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_943),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_532),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_457),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_936),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_328),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_897),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_26),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_852),
.Y(n_1417)
);

BUFx10_ASAP7_75t_L g1418 ( 
.A(n_549),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_548),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_235),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_838),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_921),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_56),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_127),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_175),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_640),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_475),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_609),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_135),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_153),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_779),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_742),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_291),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_855),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_818),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_144),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_780),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_243),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_894),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_868),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_881),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_129),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_864),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_909),
.Y(n_1444)
);

BUFx5_ASAP7_75t_L g1445 ( 
.A(n_573),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_348),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_384),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_331),
.Y(n_1448)
);

BUFx10_ASAP7_75t_L g1449 ( 
.A(n_913),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_923),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_903),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_370),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_532),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_359),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_624),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_132),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_698),
.Y(n_1457)
);

CKINVDCx16_ASAP7_75t_R g1458 ( 
.A(n_133),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_516),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_450),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_276),
.Y(n_1461)
);

CKINVDCx16_ASAP7_75t_R g1462 ( 
.A(n_569),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_444),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_292),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_173),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_638),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_552),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_855),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_567),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_862),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_117),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_692),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_726),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_579),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_859),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_427),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_235),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_641),
.Y(n_1478)
);

CKINVDCx16_ASAP7_75t_R g1479 ( 
.A(n_427),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_938),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_894),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_806),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_853),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_353),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_653),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_904),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_903),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_129),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_282),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_278),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_643),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_813),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_492),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_385),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_805),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_861),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_150),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_906),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_271),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_409),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_767),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_189),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_79),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_705),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_144),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_417),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_520),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_322),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_310),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_948),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_489),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_187),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_710),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_302),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_302),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_214),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_575),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_407),
.Y(n_1518)
);

CKINVDCx14_ASAP7_75t_R g1519 ( 
.A(n_16),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_874),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_61),
.Y(n_1521)
);

CKINVDCx16_ASAP7_75t_R g1522 ( 
.A(n_908),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_893),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_112),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_257),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_8),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_152),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_872),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_150),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_463),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_932),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_368),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_680),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_89),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_562),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_852),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_905),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_891),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_608),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_778),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_785),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_530),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_182),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_341),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_444),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_461),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_487),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_941),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_364),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_889),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_953),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_848),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_271),
.Y(n_1553)
);

BUFx10_ASAP7_75t_L g1554 ( 
.A(n_853),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_575),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_898),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_272),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_2),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_870),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1019),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1146),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1019),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1068),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1146),
.Y(n_1564)
);

CKINVDCx20_ASAP7_75t_R g1565 ( 
.A(n_1519),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1519),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1129),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1420),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1179),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1079),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1179),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1234),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1234),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_990),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1442),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1169),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1311),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1169),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1296),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1452),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1132),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1215),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1354),
.B(n_1),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1311),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1263),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1008),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1263),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1072),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1067),
.B(n_0),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1484),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_975),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1078),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1095),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1008),
.Y(n_1594)
);

INVxp67_ASAP7_75t_SL g1595 ( 
.A(n_1058),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1270),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1458),
.B(n_0),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1078),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_985),
.Y(n_1599)
);

CKINVDCx16_ASAP7_75t_R g1600 ( 
.A(n_1479),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1078),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_993),
.Y(n_1602)
);

INVxp33_ASAP7_75t_SL g1603 ( 
.A(n_980),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_962),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_967),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1000),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1001),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1005),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1058),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1010),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_968),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_977),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1038),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1069),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1207),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1207),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1075),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1258),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1076),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1091),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1092),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1104),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1107),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1108),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_986),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1123),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1136),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_988),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1265),
.B(n_0),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1143),
.Y(n_1630)
);

INVxp33_ASAP7_75t_SL g1631 ( 
.A(n_1126),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_989),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1153),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1162),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1124),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1238),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1258),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1171),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1172),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1186),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1188),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1216),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1219),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1262),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_991),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1124),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1296),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_994),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1078),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1222),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_995),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1346),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1223),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1262),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_997),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1231),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1233),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1237),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1003),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1441),
.B(n_1),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1006),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1013),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1533),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1240),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1078),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1016),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1248),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1508),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1254),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1266),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1276),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1017),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1283),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1138),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1285),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1303),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1338),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1300),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1020),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1352),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1027),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1300),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1366),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1374),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1376),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1385),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1386),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1340),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_963),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1078),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1682),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1579),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1570),
.B(n_963),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1609),
.B(n_1028),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1579),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1600),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1579),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1594),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1647),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1609),
.B(n_1030),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1592),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1598),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1601),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1647),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1582),
.B(n_963),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1574),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1563),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1678),
.B(n_1032),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1604),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1678),
.B(n_1040),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1586),
.B(n_1041),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1668),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1594),
.B(n_1044),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1589),
.B(n_1046),
.C(n_1045),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1576),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1605),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1649),
.A2(n_1112),
.B(n_1111),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1560),
.Y(n_1718)
);

OA21x2_ASAP7_75t_L g1719 ( 
.A1(n_1665),
.A2(n_1112),
.B(n_1111),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1647),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1595),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1562),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1690),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1567),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1595),
.Y(n_1725)
);

BUFx8_ASAP7_75t_L g1726 ( 
.A(n_1652),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1635),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1635),
.Y(n_1728)
);

INVx5_ASAP7_75t_L g1729 ( 
.A(n_1646),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1646),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1689),
.B(n_1052),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1568),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1575),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1611),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1580),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1612),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1591),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1663),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1599),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1561),
.B(n_1057),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1625),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1636),
.B(n_1039),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1564),
.B(n_1059),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1581),
.B(n_1042),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1602),
.B(n_1060),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1606),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1607),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1608),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1610),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1613),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1628),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1590),
.B(n_1583),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1614),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1617),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1632),
.B(n_1039),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1619),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1620),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1621),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1622),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1623),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1624),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1578),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1626),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1627),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1645),
.B(n_1039),
.Y(n_1765)
);

XNOR2xp5_ASAP7_75t_L g1766 ( 
.A(n_1615),
.B(n_1342),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1630),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1648),
.B(n_979),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1633),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1634),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1638),
.Y(n_1771)
);

AND2x2_ASAP7_75t_SL g1772 ( 
.A(n_1597),
.B(n_1085),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1639),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1569),
.B(n_1093),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1640),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1641),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1642),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1643),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1650),
.Y(n_1779)
);

AND3x1_ASAP7_75t_L g1780 ( 
.A(n_1629),
.B(n_1145),
.C(n_1130),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1653),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1656),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1657),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1658),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1664),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1667),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1660),
.B(n_1148),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1669),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1651),
.B(n_1206),
.Y(n_1789)
);

OA21x2_ASAP7_75t_L g1790 ( 
.A1(n_1670),
.A2(n_1137),
.B(n_1120),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1671),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1673),
.B(n_1257),
.Y(n_1792)
);

AND2x6_ASAP7_75t_L g1793 ( 
.A(n_1675),
.B(n_1350),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1676),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1677),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1680),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1683),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1684),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1655),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1685),
.B(n_1064),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1686),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1659),
.B(n_1462),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1687),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1661),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1571),
.B(n_1065),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1662),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1572),
.B(n_1359),
.Y(n_1807)
);

BUFx3_ASAP7_75t_L g1808 ( 
.A(n_1666),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1672),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1573),
.B(n_1393),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1679),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1616),
.A2(n_1408),
.B1(n_1459),
.B2(n_1379),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1681),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1577),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1584),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1588),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1593),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1603),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1631),
.A2(n_1137),
.B(n_1120),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1596),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1565),
.B(n_1522),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1566),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1585),
.Y(n_1823)
);

AOI22x1_ASAP7_75t_L g1824 ( 
.A1(n_1587),
.A2(n_1333),
.B1(n_1351),
.B2(n_1239),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1618),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1674),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1637),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1644),
.B(n_1550),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1654),
.B(n_1070),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1688),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1574),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1592),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1592),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1581),
.B(n_990),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1581),
.B(n_1043),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1570),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1574),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1574),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1574),
.Y(n_1839)
);

BUFx8_ASAP7_75t_L g1840 ( 
.A(n_1652),
.Y(n_1840)
);

BUFx6f_ASAP7_75t_L g1841 ( 
.A(n_1579),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1574),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1592),
.Y(n_1843)
);

AND3x2_ASAP7_75t_L g1844 ( 
.A(n_1570),
.B(n_1278),
.C(n_1239),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1563),
.B(n_1073),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1570),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1592),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1563),
.B(n_1074),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1574),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1682),
.B(n_1081),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1682),
.B(n_1097),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1574),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1574),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1574),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1574),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1592),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1574),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1592),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1574),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1682),
.B(n_1105),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1570),
.B(n_1350),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1579),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1581),
.B(n_1043),
.Y(n_1863)
);

XNOR2x2_ASAP7_75t_R g1864 ( 
.A(n_1576),
.B(n_1),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1563),
.B(n_1113),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1574),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1563),
.B(n_1116),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1570),
.Y(n_1868)
);

CKINVDCx11_ASAP7_75t_R g1869 ( 
.A(n_1576),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1570),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1570),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1574),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1592),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1592),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1592),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1594),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1594),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1574),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1570),
.B(n_1407),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1574),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1594),
.Y(n_1881)
);

CKINVDCx11_ASAP7_75t_R g1882 ( 
.A(n_1576),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1574),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1570),
.B(n_1407),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1563),
.B(n_1117),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1574),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1574),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1570),
.B(n_1448),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1570),
.B(n_1448),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1574),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1594),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1574),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1574),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1579),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1594),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1682),
.B(n_1125),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1574),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1574),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1563),
.B(n_1127),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1579),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1594),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1594),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1594),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1574),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1729),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1724),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1739),
.B(n_1135),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1846),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1869),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1729),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1729),
.Y(n_1911)
);

BUFx3_ASAP7_75t_L g1912 ( 
.A(n_1709),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1761),
.B(n_1139),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1752),
.A2(n_1141),
.B1(n_1149),
.B2(n_1140),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1774),
.B(n_1156),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1717),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1790),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1781),
.B(n_1157),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1732),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1733),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1790),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1735),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1819),
.Y(n_1923)
);

BUFx3_ASAP7_75t_L g1924 ( 
.A(n_1709),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1788),
.B(n_1158),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1719),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1752),
.A2(n_1161),
.B1(n_1168),
.B2(n_1159),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1791),
.B(n_1178),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1707),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1724),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1718),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1734),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1698),
.A2(n_1400),
.B1(n_1416),
.B2(n_1394),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1722),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1721),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1836),
.B(n_974),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1725),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1719),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1727),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1831),
.Y(n_1940)
);

AND2x6_ASAP7_75t_L g1941 ( 
.A(n_1755),
.B(n_1333),
.Y(n_1941)
);

AND2x6_ASAP7_75t_L g1942 ( 
.A(n_1765),
.B(n_1351),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1728),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1749),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1730),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1838),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1749),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1868),
.Y(n_1948)
);

OR2x6_ASAP7_75t_L g1949 ( 
.A(n_1734),
.B(n_1490),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1750),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1870),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1826),
.B(n_996),
.Y(n_1952)
);

OR2x6_ASAP7_75t_L g1953 ( 
.A(n_1830),
.B(n_996),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1876),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1787),
.B(n_1373),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1882),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1859),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1750),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1787),
.B(n_1373),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1694),
.B(n_1182),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1877),
.Y(n_1961)
);

INVx4_ASAP7_75t_L g1962 ( 
.A(n_1793),
.Y(n_1962)
);

NAND2xp33_ASAP7_75t_L g1963 ( 
.A(n_1793),
.B(n_1078),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1741),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1778),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1778),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1801),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1693),
.B(n_1433),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1801),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1881),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1871),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1706),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1837),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1731),
.B(n_1433),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1712),
.B(n_974),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1891),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1839),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1793),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1895),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1901),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1842),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1849),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1902),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1691),
.B(n_1184),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1738),
.Y(n_1985)
);

NAND3xp33_ASAP7_75t_L g1986 ( 
.A(n_1824),
.B(n_1194),
.C(n_1192),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1903),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1700),
.B(n_1202),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1792),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1792),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1740),
.B(n_1454),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1743),
.B(n_1454),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1852),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1853),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1742),
.A2(n_1217),
.B1(n_1220),
.B2(n_1213),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1854),
.Y(n_1996)
);

OAI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1716),
.A2(n_999),
.B1(n_1180),
.B2(n_1002),
.Y(n_1997)
);

INVx4_ASAP7_75t_L g1998 ( 
.A(n_1866),
.Y(n_1998)
);

INVx3_ASAP7_75t_L g1999 ( 
.A(n_1855),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1747),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_1713),
.A2(n_1438),
.B1(n_1447),
.B2(n_1423),
.Y(n_2001)
);

BUFx2_ASAP7_75t_L g2002 ( 
.A(n_1726),
.Y(n_2002)
);

INVx3_ASAP7_75t_L g2003 ( 
.A(n_1857),
.Y(n_2003)
);

BUFx10_ASAP7_75t_L g2004 ( 
.A(n_1696),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1748),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1754),
.Y(n_2006)
);

BUFx2_ASAP7_75t_L g2007 ( 
.A(n_1726),
.Y(n_2007)
);

INVx1_ASAP7_75t_SL g2008 ( 
.A(n_1861),
.Y(n_2008)
);

INVx4_ASAP7_75t_L g2009 ( 
.A(n_1890),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1872),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1805),
.B(n_1224),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1708),
.B(n_1226),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1878),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1880),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1883),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1705),
.B(n_1229),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1879),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1757),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1884),
.B(n_974),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1824),
.A2(n_1460),
.B1(n_1461),
.B2(n_1456),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1759),
.A2(n_1477),
.B1(n_1488),
.B2(n_1476),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1710),
.B(n_1230),
.Y(n_2022)
);

AOI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1760),
.A2(n_1511),
.B1(n_1516),
.B2(n_1506),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1773),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1711),
.B(n_1235),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1775),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1829),
.B(n_1888),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1776),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1808),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1889),
.B(n_1012),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1886),
.Y(n_2031)
);

INVx5_ASAP7_75t_L g2032 ( 
.A(n_1723),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1714),
.B(n_1241),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1806),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1887),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1745),
.B(n_1800),
.Y(n_2036)
);

AOI21x1_ASAP7_75t_L g2037 ( 
.A1(n_1701),
.A2(n_1526),
.B(n_1518),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1744),
.B(n_1251),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1813),
.B(n_1253),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1807),
.B(n_1256),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1777),
.A2(n_1534),
.B1(n_1545),
.B2(n_1529),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_1818),
.B(n_1062),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_1736),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1737),
.B(n_1260),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1807),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1810),
.B(n_1261),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_1892),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1893),
.Y(n_2048)
);

OR2x6_ASAP7_75t_L g2049 ( 
.A(n_1828),
.B(n_1806),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1746),
.B(n_1753),
.Y(n_2050)
);

AND3x2_ASAP7_75t_L g2051 ( 
.A(n_1864),
.B(n_1002),
.C(n_999),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_SL g2052 ( 
.A(n_1751),
.B(n_1180),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1897),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1810),
.B(n_1264),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1779),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1782),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_SL g2057 ( 
.A(n_1799),
.B(n_1267),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1898),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1784),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1794),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1840),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1744),
.B(n_1268),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1772),
.B(n_1012),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_L g2064 ( 
.A(n_1812),
.B(n_1100),
.C(n_1080),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1795),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1904),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_1756),
.A2(n_1558),
.B1(n_1553),
.B2(n_1014),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1758),
.B(n_1543),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1723),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1763),
.B(n_1544),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1764),
.B(n_1546),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_SL g2072 ( 
.A(n_1828),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_1767),
.A2(n_1014),
.B1(n_1050),
.B2(n_1004),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1769),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1770),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1771),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1783),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1785),
.B(n_1547),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1786),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1796),
.B(n_1549),
.Y(n_2080)
);

BUFx8_ASAP7_75t_SL g2081 ( 
.A(n_1715),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1797),
.B(n_1557),
.Y(n_2082)
);

INVx5_ASAP7_75t_L g2083 ( 
.A(n_1692),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1798),
.B(n_1281),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1900),
.Y(n_2085)
);

INVxp67_ASAP7_75t_SL g2086 ( 
.A(n_1850),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1803),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1701),
.Y(n_2088)
);

NAND3xp33_ASAP7_75t_L g2089 ( 
.A(n_1851),
.B(n_1292),
.C(n_1291),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1860),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1692),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1702),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1896),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1834),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1768),
.B(n_1012),
.Y(n_2095)
);

AND3x2_ASAP7_75t_L g2096 ( 
.A(n_1821),
.B(n_1214),
.C(n_1187),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1834),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1835),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1702),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1815),
.B(n_1293),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1789),
.B(n_1175),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1840),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1804),
.B(n_1305),
.Y(n_2103)
);

INVxp33_ASAP7_75t_L g2104 ( 
.A(n_1766),
.Y(n_2104)
);

OR2x6_ASAP7_75t_L g2105 ( 
.A(n_1823),
.B(n_1187),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_1802),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1845),
.B(n_1848),
.Y(n_2107)
);

OAI22xp33_ASAP7_75t_SL g2108 ( 
.A1(n_1827),
.A2(n_1307),
.B1(n_1310),
.B2(n_1306),
.Y(n_2108)
);

AND2x6_ASAP7_75t_L g2109 ( 
.A(n_1809),
.B(n_1004),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_1811),
.B(n_1816),
.Y(n_2110)
);

AOI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_1865),
.A2(n_1313),
.B1(n_1316),
.B2(n_1312),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1835),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1863),
.Y(n_2113)
);

BUFx10_ASAP7_75t_L g2114 ( 
.A(n_1823),
.Y(n_2114)
);

NAND2xp33_ASAP7_75t_L g2115 ( 
.A(n_1814),
.B(n_1221),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1863),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1900),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1703),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1703),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_1820),
.Y(n_2120)
);

OR2x6_ASAP7_75t_L g2121 ( 
.A(n_1822),
.B(n_1214),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_1817),
.B(n_1322),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_1780),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1832),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1867),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1885),
.B(n_1324),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1762),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1832),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_1844),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1899),
.Y(n_2130)
);

INVxp67_ASAP7_75t_SL g2131 ( 
.A(n_1833),
.Y(n_2131)
);

OAI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_1827),
.A2(n_1250),
.B1(n_1339),
.B2(n_1243),
.Y(n_2132)
);

NAND2xp33_ASAP7_75t_L g2133 ( 
.A(n_1833),
.B(n_1221),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_1766),
.Y(n_2134)
);

INVx4_ASAP7_75t_L g2135 ( 
.A(n_1843),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_1825),
.B(n_1392),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1843),
.B(n_1328),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_1847),
.B(n_1331),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1847),
.B(n_1856),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1856),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_1858),
.B(n_1414),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_1858),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1873),
.Y(n_2143)
);

OAI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1873),
.A2(n_1061),
.B(n_965),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1874),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1874),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1875),
.Y(n_2147)
);

BUFx8_ASAP7_75t_SL g2148 ( 
.A(n_1695),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1875),
.B(n_1334),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_1695),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_1697),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_1697),
.Y(n_2152)
);

AOI22xp33_ASAP7_75t_L g2153 ( 
.A1(n_1699),
.A2(n_1014),
.B1(n_1050),
.B2(n_1004),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1699),
.Y(n_2154)
);

NAND2x1p5_ASAP7_75t_L g2155 ( 
.A(n_1704),
.B(n_1464),
.Y(n_2155)
);

OR2x6_ASAP7_75t_L g2156 ( 
.A(n_1704),
.B(n_1243),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1720),
.B(n_1336),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_1720),
.B(n_1337),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_1841),
.A2(n_1014),
.B1(n_1050),
.B2(n_1004),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1841),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1862),
.B(n_1345),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1862),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1894),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1894),
.B(n_1356),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1729),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1729),
.Y(n_2166)
);

INVx3_ASAP7_75t_L g2167 ( 
.A(n_1724),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1717),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_1724),
.Y(n_2169)
);

INVx3_ASAP7_75t_L g2170 ( 
.A(n_1724),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_SL g2171 ( 
.A(n_1826),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1787),
.B(n_1357),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_1709),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1774),
.B(n_1361),
.Y(n_2174)
);

BUFx3_ASAP7_75t_L g2175 ( 
.A(n_1709),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1729),
.Y(n_2176)
);

INVxp67_ASAP7_75t_SL g2177 ( 
.A(n_1836),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1739),
.B(n_1363),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1717),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1787),
.B(n_1372),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1729),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1709),
.Y(n_2182)
);

XNOR2xp5_ASAP7_75t_L g2183 ( 
.A(n_1766),
.B(n_1250),
.Y(n_2183)
);

INVx4_ASAP7_75t_L g2184 ( 
.A(n_1793),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1739),
.B(n_1383),
.Y(n_2185)
);

AOI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_1698),
.A2(n_1177),
.B1(n_1302),
.B2(n_1050),
.Y(n_2186)
);

OR2x6_ASAP7_75t_L g2187 ( 
.A(n_1709),
.B(n_1339),
.Y(n_2187)
);

NOR2x1p5_ASAP7_75t_L g2188 ( 
.A(n_1696),
.B(n_1388),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1774),
.B(n_1389),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1717),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1729),
.Y(n_2191)
);

INVx3_ASAP7_75t_L g2192 ( 
.A(n_1724),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_1752),
.A2(n_1401),
.B1(n_1403),
.B2(n_1398),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1729),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1717),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1729),
.Y(n_2196)
);

NAND2xp33_ASAP7_75t_SL g2197 ( 
.A(n_1709),
.B(n_1404),
.Y(n_2197)
);

INVx2_ASAP7_75t_SL g2198 ( 
.A(n_1846),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_1698),
.A2(n_1177),
.B1(n_1362),
.B2(n_1302),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1729),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1729),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1717),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_1698),
.A2(n_1177),
.B1(n_1362),
.B2(n_1302),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_1971),
.B(n_1515),
.Y(n_2204)
);

AND2x4_ASAP7_75t_SL g2205 ( 
.A(n_2114),
.B(n_1175),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1951),
.B(n_1412),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2086),
.B(n_1424),
.Y(n_2207)
);

INVx2_ASAP7_75t_SL g2208 ( 
.A(n_1912),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2141),
.B(n_1425),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2135),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2135),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2036),
.B(n_1427),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1935),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_2198),
.B(n_1497),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2177),
.A2(n_1430),
.B1(n_1436),
.B2(n_1429),
.Y(n_2215)
);

OR2x6_ASAP7_75t_L g2216 ( 
.A(n_1949),
.B(n_965),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_L g2217 ( 
.A(n_1978),
.Y(n_2217)
);

INVx2_ASAP7_75t_SL g2218 ( 
.A(n_1924),
.Y(n_2218)
);

AOI22xp33_ASAP7_75t_L g2219 ( 
.A1(n_2125),
.A2(n_1190),
.B1(n_1197),
.B2(n_1176),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_1985),
.B(n_1446),
.Y(n_2220)
);

NAND3xp33_ASAP7_75t_L g2221 ( 
.A(n_1915),
.B(n_1465),
.C(n_1463),
.Y(n_2221)
);

INVx3_ASAP7_75t_L g2222 ( 
.A(n_1932),
.Y(n_2222)
);

NOR3xp33_ASAP7_75t_L g2223 ( 
.A(n_1997),
.B(n_1244),
.C(n_1181),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1937),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1939),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2090),
.B(n_1471),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1978),
.Y(n_2227)
);

NOR2xp67_ASAP7_75t_L g2228 ( 
.A(n_2123),
.B(n_2),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2145),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_SL g2230 ( 
.A(n_2043),
.B(n_969),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_1948),
.B(n_1175),
.Y(n_2231)
);

NOR3xp33_ASAP7_75t_L g2232 ( 
.A(n_2132),
.B(n_1539),
.C(n_1411),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1943),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2093),
.B(n_1489),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1945),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1978),
.B(n_1962),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2130),
.B(n_1493),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2142),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_1962),
.B(n_1505),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2025),
.B(n_1494),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2142),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2184),
.B(n_1908),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2131),
.B(n_1499),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_2173),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2138),
.B(n_1500),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2088),
.Y(n_2246)
);

NOR2xp67_ASAP7_75t_L g2247 ( 
.A(n_2123),
.B(n_2),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2050),
.B(n_1502),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_2184),
.B(n_1514),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_2175),
.B(n_1530),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1954),
.B(n_1503),
.Y(n_2251)
);

CKINVDCx20_ASAP7_75t_R g2252 ( 
.A(n_2081),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1961),
.B(n_1532),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1970),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1976),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1979),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2092),
.Y(n_2257)
);

OAI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_2027),
.A2(n_1037),
.B1(n_1082),
.B2(n_1034),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1980),
.B(n_1507),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1983),
.B(n_1509),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_2192),
.Y(n_2261)
);

INVx5_ASAP7_75t_L g2262 ( 
.A(n_2148),
.Y(n_2262)
);

BUFx4f_ASAP7_75t_L g2263 ( 
.A(n_2002),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1987),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1989),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2182),
.B(n_1277),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2099),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2044),
.B(n_1512),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1990),
.Y(n_2269)
);

INVx2_ASAP7_75t_SL g2270 ( 
.A(n_1964),
.Y(n_2270)
);

INVx2_ASAP7_75t_SL g2271 ( 
.A(n_2114),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2068),
.B(n_1521),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2197),
.B(n_1524),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2057),
.B(n_1525),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2070),
.B(n_1527),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2078),
.B(n_970),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2008),
.B(n_1277),
.Y(n_2277)
);

NOR3xp33_ASAP7_75t_L g2278 ( 
.A(n_2108),
.B(n_2064),
.C(n_2106),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2029),
.B(n_972),
.Y(n_2279)
);

OAI22xp33_ASAP7_75t_L g2280 ( 
.A1(n_2052),
.A2(n_1369),
.B1(n_1397),
.B2(n_1114),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_1984),
.B(n_973),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2139),
.A2(n_1528),
.B1(n_1439),
.B2(n_966),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2001),
.A2(n_971),
.B1(n_978),
.B2(n_964),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_2110),
.B(n_976),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_1949),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2118),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2019),
.B(n_1277),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2030),
.B(n_1325),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2074),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2080),
.B(n_981),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2075),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2082),
.B(n_983),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1960),
.B(n_984),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2077),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_1914),
.B(n_1325),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2095),
.B(n_992),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_1988),
.B(n_1007),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2012),
.B(n_1011),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2079),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2101),
.B(n_1021),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2119),
.Y(n_2301)
);

INVx3_ASAP7_75t_L g2302 ( 
.A(n_2192),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_2061),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2076),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_1927),
.B(n_1325),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_2022),
.B(n_1022),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2087),
.B(n_1026),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2193),
.B(n_1418),
.Y(n_2308)
);

AOI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_1995),
.A2(n_1035),
.B1(n_1036),
.B2(n_1033),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_2102),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2042),
.B(n_1418),
.Y(n_2311)
);

INVx4_ASAP7_75t_L g2312 ( 
.A(n_2049),
.Y(n_2312)
);

NOR3xp33_ASAP7_75t_L g2313 ( 
.A(n_2134),
.B(n_1327),
.C(n_1048),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2124),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_2172),
.B(n_1047),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2089),
.B(n_1053),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_1907),
.B(n_1054),
.Y(n_2317)
);

INVx2_ASAP7_75t_SL g2318 ( 
.A(n_2049),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2045),
.B(n_982),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_1913),
.B(n_1918),
.Y(n_2320)
);

AOI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2180),
.A2(n_1071),
.B1(n_1077),
.B2(n_1055),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2097),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2149),
.B(n_1083),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2016),
.B(n_1086),
.Y(n_2324)
);

INVx2_ASAP7_75t_SL g2325 ( 
.A(n_2156),
.Y(n_2325)
);

BUFx12f_ASAP7_75t_L g2326 ( 
.A(n_1909),
.Y(n_2326)
);

INVxp33_ASAP7_75t_L g2327 ( 
.A(n_2136),
.Y(n_2327)
);

HB1xp67_ASAP7_75t_L g2328 ( 
.A(n_2156),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2098),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2017),
.B(n_1418),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_1925),
.B(n_1087),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2128),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1919),
.B(n_1089),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2140),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1920),
.B(n_1090),
.Y(n_2335)
);

NOR2x1_ASAP7_75t_L g2336 ( 
.A(n_2188),
.B(n_1176),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1928),
.B(n_2178),
.Y(n_2337)
);

AOI22xp33_ASAP7_75t_L g2338 ( 
.A1(n_1941),
.A2(n_1190),
.B1(n_1320),
.B2(n_1197),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1922),
.B(n_1094),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_1956),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2185),
.B(n_1098),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2174),
.B(n_1101),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2143),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_2107),
.B(n_1102),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_2187),
.Y(n_2345)
);

AOI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_1916),
.A2(n_998),
.B(n_987),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2189),
.B(n_1106),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2063),
.B(n_1449),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1955),
.B(n_1959),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2112),
.Y(n_2350)
);

NAND3xp33_ASAP7_75t_L g2351 ( 
.A(n_2103),
.B(n_1118),
.C(n_1115),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2113),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2116),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_2040),
.B(n_2046),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2147),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2054),
.B(n_1936),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2168),
.A2(n_1015),
.B(n_1009),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2000),
.B(n_1119),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2094),
.Y(n_2359)
);

NOR3x1_ASAP7_75t_L g2360 ( 
.A(n_2007),
.B(n_1023),
.C(n_1018),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2094),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2005),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2006),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2018),
.B(n_1128),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_SL g2365 ( 
.A(n_2004),
.B(n_1449),
.Y(n_2365)
);

AOI22xp5_ASAP7_75t_L g2366 ( 
.A1(n_1975),
.A2(n_1133),
.B1(n_1144),
.B2(n_1131),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2024),
.B(n_1151),
.Y(n_2367)
);

NAND3xp33_ASAP7_75t_L g2368 ( 
.A(n_2100),
.B(n_1163),
.C(n_1160),
.Y(n_2368)
);

AND2x4_ASAP7_75t_SL g2369 ( 
.A(n_2004),
.B(n_1449),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2187),
.B(n_1554),
.Y(n_2370)
);

NOR2xp67_ASAP7_75t_SL g2371 ( 
.A(n_2032),
.B(n_1164),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1917),
.Y(n_2372)
);

AND2x2_ASAP7_75t_SL g2373 ( 
.A(n_2051),
.B(n_1061),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2026),
.B(n_1166),
.Y(n_2374)
);

BUFx6f_ASAP7_75t_L g2375 ( 
.A(n_1921),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2028),
.B(n_1167),
.Y(n_2376)
);

NOR2xp33_ASAP7_75t_L g2377 ( 
.A(n_1968),
.B(n_1170),
.Y(n_2377)
);

AOI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_1941),
.A2(n_1326),
.B1(n_1344),
.B2(n_1320),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2055),
.B(n_1173),
.Y(n_2379)
);

INVxp67_ASAP7_75t_SL g2380 ( 
.A(n_1926),
.Y(n_2380)
);

NAND3xp33_ASAP7_75t_L g2381 ( 
.A(n_2038),
.B(n_1185),
.C(n_1174),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1938),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2146),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_1905),
.B(n_1193),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2056),
.B(n_1196),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_1910),
.B(n_1199),
.Y(n_2386)
);

INVx3_ASAP7_75t_L g2387 ( 
.A(n_1911),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2059),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2060),
.B(n_1200),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2065),
.B(n_1203),
.Y(n_2390)
);

INVx2_ASAP7_75t_SL g2391 ( 
.A(n_2034),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2111),
.B(n_1208),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_2165),
.B(n_1209),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2166),
.B(n_1212),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_2176),
.B(n_1218),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_1941),
.B(n_1232),
.Y(n_2396)
);

BUFx6f_ASAP7_75t_L g2397 ( 
.A(n_2085),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2181),
.B(n_1236),
.Y(n_2398)
);

OR2x6_ASAP7_75t_L g2399 ( 
.A(n_1952),
.B(n_1110),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_1941),
.B(n_1942),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_1931),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2191),
.B(n_1242),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1934),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_2194),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2196),
.B(n_1247),
.Y(n_2405)
);

INVx2_ASAP7_75t_SL g2406 ( 
.A(n_2155),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1929),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_1942),
.B(n_1249),
.Y(n_2408)
);

NOR3xp33_ASAP7_75t_L g2409 ( 
.A(n_2129),
.B(n_2127),
.C(n_2011),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1923),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_1972),
.Y(n_2411)
);

NOR2xp33_ASAP7_75t_L g2412 ( 
.A(n_2062),
.B(n_1259),
.Y(n_2412)
);

INVx5_ASAP7_75t_L g2413 ( 
.A(n_2109),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2120),
.B(n_1269),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2200),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2201),
.B(n_1272),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_1973),
.Y(n_2417)
);

AND2x6_ASAP7_75t_L g2418 ( 
.A(n_2179),
.B(n_1177),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2105),
.B(n_1554),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_2122),
.B(n_1273),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2126),
.B(n_1275),
.Y(n_2421)
);

INVxp67_ASAP7_75t_L g2422 ( 
.A(n_2105),
.Y(n_2422)
);

INVx2_ASAP7_75t_SL g2423 ( 
.A(n_1998),
.Y(n_2423)
);

AO22x2_ASAP7_75t_L g2424 ( 
.A1(n_2183),
.A2(n_1025),
.B1(n_1029),
.B2(n_1024),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_1942),
.B(n_1279),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_1953),
.B(n_1554),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_1942),
.B(n_1280),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_1933),
.B(n_1282),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1977),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2039),
.B(n_1284),
.Y(n_2430)
);

INVxp33_ASAP7_75t_SL g2431 ( 
.A(n_2072),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_1953),
.B(n_1286),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2071),
.B(n_1031),
.Y(n_2433)
);

INVx4_ASAP7_75t_L g2434 ( 
.A(n_2032),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_1974),
.B(n_1287),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_2032),
.B(n_1289),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_1986),
.B(n_1998),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2021),
.B(n_2023),
.Y(n_2438)
);

AOI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2084),
.A2(n_1299),
.B1(n_1301),
.B2(n_1295),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2009),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2041),
.B(n_1308),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_SL g2442 ( 
.A(n_2009),
.B(n_1309),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_1940),
.B(n_1314),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1991),
.B(n_1315),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2020),
.B(n_1317),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1982),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_1993),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_1946),
.B(n_1318),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_1992),
.B(n_1321),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2033),
.B(n_1323),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_1994),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_1957),
.B(n_1329),
.Y(n_2452)
);

BUFx6f_ASAP7_75t_L g2453 ( 
.A(n_2085),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_1996),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2013),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2015),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2031),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2137),
.B(n_1330),
.Y(n_2458)
);

AOI22xp33_ASAP7_75t_L g2459 ( 
.A1(n_2067),
.A2(n_2144),
.B1(n_2048),
.B2(n_2058),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_1952),
.B(n_2121),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2121),
.B(n_1335),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2164),
.B(n_1341),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2035),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_1981),
.B(n_1347),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1981),
.B(n_1348),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2066),
.Y(n_2466)
);

OAI21xp5_ASAP7_75t_L g2467 ( 
.A1(n_2190),
.A2(n_1051),
.B(n_1049),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1999),
.B(n_1349),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1999),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2195),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_1906),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2003),
.Y(n_2472)
);

INVx2_ASAP7_75t_SL g2473 ( 
.A(n_2167),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2003),
.B(n_1358),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2010),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2010),
.B(n_1360),
.Y(n_2476)
);

O2A1O1Ixp5_ASAP7_75t_L g2477 ( 
.A1(n_2157),
.A2(n_2202),
.B(n_2037),
.C(n_2161),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_1930),
.B(n_2158),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2096),
.B(n_1364),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2014),
.B(n_1365),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2014),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2047),
.B(n_2053),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2053),
.B(n_2169),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2170),
.B(n_1367),
.Y(n_2484)
);

AOI22xp5_ASAP7_75t_L g2485 ( 
.A1(n_1963),
.A2(n_1370),
.B1(n_1381),
.B2(n_1368),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_1944),
.B(n_1382),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2104),
.B(n_1387),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2115),
.B(n_1390),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2037),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_1947),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2171),
.B(n_1391),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_1950),
.B(n_1395),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2109),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_1958),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_1965),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_1966),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_1967),
.B(n_1405),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_1969),
.B(n_1406),
.Y(n_2498)
);

INVx2_ASAP7_75t_SL g2499 ( 
.A(n_2109),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2186),
.B(n_1399),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2203),
.B(n_1410),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2199),
.B(n_1413),
.Y(n_2502)
);

AND2x4_ASAP7_75t_L g2503 ( 
.A(n_2151),
.B(n_1056),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2133),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2109),
.B(n_1415),
.Y(n_2505)
);

INVx2_ASAP7_75t_SL g2506 ( 
.A(n_2150),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2151),
.B(n_1421),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2069),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2073),
.B(n_1428),
.Y(n_2509)
);

BUFx6f_ASAP7_75t_L g2510 ( 
.A(n_2085),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2152),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2083),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2160),
.B(n_1432),
.Y(n_2513)
);

AOI22xp33_ASAP7_75t_L g2514 ( 
.A1(n_2154),
.A2(n_1326),
.B1(n_1422),
.B2(n_1344),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2083),
.Y(n_2515)
);

OR2x2_ASAP7_75t_L g2516 ( 
.A(n_2163),
.B(n_1434),
.Y(n_2516)
);

INVx2_ASAP7_75t_SL g2517 ( 
.A(n_2083),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_2091),
.B(n_2117),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2091),
.B(n_1435),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_SL g2520 ( 
.A(n_2091),
.B(n_1443),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2117),
.B(n_1444),
.Y(n_2521)
);

INVxp67_ASAP7_75t_L g2522 ( 
.A(n_2117),
.Y(n_2522)
);

CKINVDCx5p33_ASAP7_75t_R g2523 ( 
.A(n_2162),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2153),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2159),
.B(n_1451),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2135),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2086),
.B(n_1453),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2135),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_1951),
.B(n_1457),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_1971),
.B(n_1455),
.Y(n_2530)
);

NAND2xp33_ASAP7_75t_L g2531 ( 
.A(n_1978),
.B(n_1221),
.Y(n_2531)
);

INVx2_ASAP7_75t_SL g2532 ( 
.A(n_1912),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2086),
.B(n_1466),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_1935),
.Y(n_2534)
);

BUFx6f_ASAP7_75t_L g2535 ( 
.A(n_1978),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2086),
.B(n_1467),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_1971),
.B(n_1468),
.Y(n_2537)
);

INVx2_ASAP7_75t_SL g2538 ( 
.A(n_1912),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2086),
.B(n_1469),
.Y(n_2539)
);

OAI221xp5_ASAP7_75t_L g2540 ( 
.A1(n_2008),
.A2(n_1480),
.B1(n_1481),
.B2(n_1474),
.C(n_1473),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2086),
.B(n_1482),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2135),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2086),
.B(n_1485),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_1951),
.B(n_1486),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_L g2545 ( 
.A(n_1951),
.B(n_1491),
.Y(n_2545)
);

INVxp67_ASAP7_75t_L g2546 ( 
.A(n_1948),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_1971),
.B(n_1495),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_1971),
.B(n_1496),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_1951),
.B(n_1498),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_1951),
.B(n_1513),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_1951),
.B(n_1523),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2086),
.B(n_1538),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2086),
.B(n_1540),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_1935),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_1971),
.B(n_1542),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_1935),
.Y(n_2556)
);

INVx4_ASAP7_75t_L g2557 ( 
.A(n_1978),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2086),
.B(n_1548),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_1951),
.B(n_1551),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2135),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_1951),
.B(n_1552),
.Y(n_2561)
);

INVxp33_ASAP7_75t_L g2562 ( 
.A(n_1908),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_1935),
.Y(n_2563)
);

AO22x1_ASAP7_75t_L g2564 ( 
.A1(n_2061),
.A2(n_1559),
.B1(n_1556),
.B2(n_1450),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2086),
.B(n_1063),
.Y(n_2565)
);

AND2x4_ASAP7_75t_L g2566 ( 
.A(n_2086),
.B(n_1066),
.Y(n_2566)
);

OR2x6_ASAP7_75t_L g2567 ( 
.A(n_1949),
.B(n_1110),
.Y(n_2567)
);

INVxp33_ASAP7_75t_L g2568 ( 
.A(n_1908),
.Y(n_2568)
);

A2O1A1Ixp33_ASAP7_75t_L g2569 ( 
.A1(n_2036),
.A2(n_1450),
.B(n_1483),
.C(n_1422),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2086),
.B(n_1084),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_1951),
.B(n_1302),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2135),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_1951),
.B(n_1537),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2135),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2086),
.B(n_1088),
.Y(n_2575)
);

OAI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2036),
.A2(n_1099),
.B(n_1096),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_1951),
.B(n_1362),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2086),
.B(n_1103),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_1951),
.B(n_1362),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2086),
.B(n_1109),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2372),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2546),
.B(n_1531),
.Y(n_2582)
);

AOI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_2380),
.A2(n_1134),
.B(n_1121),
.Y(n_2583)
);

BUFx6f_ASAP7_75t_L g2584 ( 
.A(n_2397),
.Y(n_2584)
);

NAND2xp33_ASAP7_75t_L g2585 ( 
.A(n_2397),
.B(n_2453),
.Y(n_2585)
);

AOI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2320),
.A2(n_1147),
.B(n_1142),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2327),
.B(n_1510),
.Y(n_2587)
);

AOI21xp5_ASAP7_75t_L g2588 ( 
.A1(n_2337),
.A2(n_1155),
.B(n_1150),
.Y(n_2588)
);

INVx3_ASAP7_75t_L g2589 ( 
.A(n_2557),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2213),
.Y(n_2590)
);

AOI21xp5_ASAP7_75t_L g2591 ( 
.A1(n_2470),
.A2(n_1183),
.B(n_1165),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2557),
.Y(n_2592)
);

OAI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2212),
.A2(n_1531),
.B1(n_1483),
.B2(n_1191),
.Y(n_2593)
);

AOI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2230),
.A2(n_1195),
.B1(n_1198),
.B2(n_1189),
.Y(n_2594)
);

INVxp67_ASAP7_75t_L g2595 ( 
.A(n_2204),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2289),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_2410),
.A2(n_1204),
.B(n_1201),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_L g2598 ( 
.A(n_2562),
.B(n_1478),
.Y(n_2598)
);

AOI21xp5_ASAP7_75t_L g2599 ( 
.A1(n_2382),
.A2(n_1210),
.B(n_1205),
.Y(n_2599)
);

BUFx3_ASAP7_75t_L g2600 ( 
.A(n_2252),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2224),
.Y(n_2601)
);

AOI21xp5_ASAP7_75t_L g2602 ( 
.A1(n_2489),
.A2(n_1225),
.B(n_1211),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_SL g2603 ( 
.A(n_2365),
.B(n_1221),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2438),
.B(n_1517),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2397),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2291),
.Y(n_2606)
);

OAI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2477),
.A2(n_1228),
.B(n_1227),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2576),
.B(n_1541),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2294),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2566),
.B(n_1555),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2311),
.B(n_1245),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2299),
.B(n_1246),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2434),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2566),
.B(n_1426),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2248),
.B(n_1431),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2225),
.Y(n_2616)
);

AOI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2268),
.A2(n_1255),
.B(n_1252),
.Y(n_2617)
);

OAI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2346),
.A2(n_1274),
.B(n_1271),
.Y(n_2618)
);

NOR2x1_ASAP7_75t_L g2619 ( 
.A(n_2216),
.B(n_1288),
.Y(n_2619)
);

AND2x4_ASAP7_75t_L g2620 ( 
.A(n_2233),
.B(n_2235),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2530),
.B(n_1475),
.Y(n_2621)
);

AO21x1_ASAP7_75t_L g2622 ( 
.A1(n_2467),
.A2(n_1297),
.B(n_1290),
.Y(n_2622)
);

AOI21x1_ASAP7_75t_L g2623 ( 
.A1(n_2518),
.A2(n_1152),
.B(n_1122),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2254),
.B(n_1501),
.Y(n_2624)
);

A2O1A1Ixp33_ASAP7_75t_L g2625 ( 
.A1(n_2357),
.A2(n_1304),
.B(n_1319),
.C(n_1298),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2255),
.B(n_1332),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2256),
.B(n_1353),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2272),
.A2(n_1371),
.B(n_1355),
.Y(n_2628)
);

CKINVDCx10_ASAP7_75t_R g2629 ( 
.A(n_2216),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2264),
.B(n_2534),
.Y(n_2630)
);

AOI21x1_ASAP7_75t_L g2631 ( 
.A1(n_2437),
.A2(n_1152),
.B(n_1122),
.Y(n_2631)
);

AOI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2275),
.A2(n_1378),
.B(n_1375),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2554),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_2556),
.B(n_1380),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2568),
.B(n_1221),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2563),
.B(n_1470),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2304),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2383),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2207),
.B(n_1472),
.Y(n_2639)
);

AOI21xp5_ASAP7_75t_L g2640 ( 
.A1(n_2240),
.A2(n_1402),
.B(n_1396),
.Y(n_2640)
);

OAI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_2569),
.A2(n_1417),
.B(n_1409),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2208),
.B(n_1221),
.Y(n_2642)
);

OR2x6_ASAP7_75t_L g2643 ( 
.A(n_2567),
.B(n_1154),
.Y(n_2643)
);

O2A1O1Ixp5_ASAP7_75t_L g2644 ( 
.A1(n_2400),
.A2(n_1294),
.B(n_1377),
.C(n_1154),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2537),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2209),
.B(n_1419),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2548),
.B(n_1437),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2565),
.B(n_2570),
.Y(n_2648)
);

AOI21xp33_ASAP7_75t_L g2649 ( 
.A1(n_2529),
.A2(n_1487),
.B(n_1440),
.Y(n_2649)
);

AOI21xp5_ASAP7_75t_L g2650 ( 
.A1(n_2251),
.A2(n_1504),
.B(n_1492),
.Y(n_2650)
);

AO21x1_ASAP7_75t_L g2651 ( 
.A1(n_2504),
.A2(n_1535),
.B(n_1520),
.Y(n_2651)
);

AO21x2_ASAP7_75t_L g2652 ( 
.A1(n_2228),
.A2(n_1377),
.B(n_1294),
.Y(n_2652)
);

AOI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2282),
.A2(n_1445),
.B1(n_1221),
.B2(n_1384),
.Y(n_2653)
);

AOI21xp5_ASAP7_75t_L g2654 ( 
.A1(n_2253),
.A2(n_1384),
.B(n_1343),
.Y(n_2654)
);

AOI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2259),
.A2(n_1343),
.B(n_1296),
.Y(n_2655)
);

AOI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2260),
.A2(n_1343),
.B(n_1296),
.Y(n_2656)
);

AOI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2323),
.A2(n_1536),
.B(n_1343),
.Y(n_2657)
);

AOI21xp5_ASAP7_75t_L g2658 ( 
.A1(n_2276),
.A2(n_1536),
.B(n_1445),
.Y(n_2658)
);

AOI21xp5_ASAP7_75t_L g2659 ( 
.A1(n_2290),
.A2(n_1536),
.B(n_1445),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2218),
.B(n_1445),
.Y(n_2660)
);

AOI21xp5_ASAP7_75t_L g2661 ( 
.A1(n_2292),
.A2(n_1536),
.B(n_1445),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2453),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2297),
.A2(n_1445),
.B(n_3),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2575),
.B(n_1445),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2532),
.B(n_4),
.Y(n_2665)
);

NOR2xp67_ASAP7_75t_L g2666 ( 
.A(n_2413),
.B(n_3),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2578),
.B(n_3),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2580),
.B(n_5),
.Y(n_2668)
);

AOI22xp33_ASAP7_75t_L g2669 ( 
.A1(n_2223),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2669)
);

O2A1O1Ixp33_ASAP7_75t_L g2670 ( 
.A1(n_2237),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2243),
.B(n_2220),
.Y(n_2671)
);

AOI21xp5_ASAP7_75t_L g2672 ( 
.A1(n_2306),
.A2(n_7),
.B(n_8),
.Y(n_2672)
);

AOI21xp5_ASAP7_75t_L g2673 ( 
.A1(n_2293),
.A2(n_8),
.B(n_9),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2244),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2287),
.B(n_9),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2246),
.Y(n_2676)
);

OAI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2459),
.A2(n_9),
.B(n_10),
.Y(n_2677)
);

O2A1O1Ixp5_ASAP7_75t_L g2678 ( 
.A1(n_2316),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2288),
.B(n_10),
.Y(n_2679)
);

AOI21xp33_ASAP7_75t_L g2680 ( 
.A1(n_2544),
.A2(n_11),
.B(n_12),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_2345),
.B(n_11),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2285),
.B(n_2348),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2362),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2363),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2265),
.B(n_13),
.Y(n_2685)
);

NAND2x1_ASAP7_75t_L g2686 ( 
.A(n_2453),
.B(n_13),
.Y(n_2686)
);

AND2x6_ASAP7_75t_L g2687 ( 
.A(n_2217),
.B(n_13),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2269),
.B(n_14),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2555),
.B(n_14),
.Y(n_2689)
);

O2A1O1Ixp33_ASAP7_75t_L g2690 ( 
.A1(n_2232),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_2690)
);

O2A1O1Ixp33_ASAP7_75t_L g2691 ( 
.A1(n_2245),
.A2(n_18),
.B(n_15),
.C(n_17),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2424),
.B(n_2277),
.Y(n_2692)
);

OAI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_2257),
.A2(n_15),
.B(n_17),
.Y(n_2693)
);

INVx3_ASAP7_75t_L g2694 ( 
.A(n_2434),
.Y(n_2694)
);

A2O1A1Ixp33_ASAP7_75t_L g2695 ( 
.A1(n_2573),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2356),
.B(n_18),
.Y(n_2696)
);

NOR2x2_ASAP7_75t_L g2697 ( 
.A(n_2567),
.B(n_20),
.Y(n_2697)
);

INVx11_ASAP7_75t_L g2698 ( 
.A(n_2326),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2388),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2527),
.B(n_20),
.Y(n_2700)
);

A2O1A1Ixp33_ASAP7_75t_L g2701 ( 
.A1(n_2247),
.A2(n_2221),
.B(n_2286),
.C(n_2267),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2538),
.Y(n_2702)
);

AOI21xp33_ASAP7_75t_L g2703 ( 
.A1(n_2545),
.A2(n_21),
.B(n_22),
.Y(n_2703)
);

AOI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2298),
.A2(n_21),
.B(n_22),
.Y(n_2704)
);

OAI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2301),
.A2(n_21),
.B(n_22),
.Y(n_2705)
);

AO21x1_ASAP7_75t_L g2706 ( 
.A1(n_2278),
.A2(n_527),
.B(n_526),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2314),
.Y(n_2707)
);

OAI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2332),
.A2(n_23),
.B(n_24),
.Y(n_2708)
);

AOI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2510),
.A2(n_23),
.B(n_24),
.Y(n_2709)
);

AO21x1_ASAP7_75t_L g2710 ( 
.A1(n_2524),
.A2(n_527),
.B(n_526),
.Y(n_2710)
);

AOI21xp5_ASAP7_75t_L g2711 ( 
.A1(n_2510),
.A2(n_23),
.B(n_25),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2401),
.Y(n_2712)
);

A2O1A1Ixp33_ASAP7_75t_L g2713 ( 
.A1(n_2334),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2510),
.A2(n_25),
.B(n_27),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2533),
.B(n_2536),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2539),
.B(n_28),
.Y(n_2716)
);

A2O1A1Ixp33_ASAP7_75t_L g2717 ( 
.A1(n_2343),
.A2(n_2355),
.B(n_2412),
.C(n_2403),
.Y(n_2717)
);

NOR2xp33_ASAP7_75t_L g2718 ( 
.A(n_2422),
.B(n_28),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_L g2719 ( 
.A(n_2325),
.B(n_28),
.Y(n_2719)
);

A2O1A1Ixp33_ASAP7_75t_L g2720 ( 
.A1(n_2238),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_SL g2721 ( 
.A(n_2340),
.B(n_29),
.Y(n_2721)
);

INVx4_ASAP7_75t_L g2722 ( 
.A(n_2262),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2541),
.B(n_29),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2424),
.B(n_30),
.Y(n_2724)
);

AOI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2375),
.A2(n_30),
.B(n_31),
.Y(n_2725)
);

OAI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2241),
.A2(n_31),
.B(n_32),
.Y(n_2726)
);

AOI21xp5_ASAP7_75t_L g2727 ( 
.A1(n_2375),
.A2(n_33),
.B(n_34),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2543),
.B(n_33),
.Y(n_2728)
);

NOR2xp33_ASAP7_75t_L g2729 ( 
.A(n_2487),
.B(n_33),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2322),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_2303),
.Y(n_2731)
);

AOI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2375),
.A2(n_34),
.B(n_35),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2329),
.Y(n_2733)
);

O2A1O1Ixp33_ASAP7_75t_L g2734 ( 
.A1(n_2283),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2552),
.B(n_2553),
.Y(n_2735)
);

NOR2x1_ASAP7_75t_R g2736 ( 
.A(n_2262),
.B(n_35),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2258),
.B(n_36),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2421),
.A2(n_37),
.B(n_38),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2350),
.Y(n_2739)
);

AOI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2558),
.A2(n_37),
.B(n_38),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_L g2741 ( 
.A(n_2328),
.B(n_2206),
.Y(n_2741)
);

AOI21xp5_ASAP7_75t_L g2742 ( 
.A1(n_2284),
.A2(n_38),
.B(n_39),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2214),
.B(n_39),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2231),
.B(n_40),
.Y(n_2744)
);

AOI22x1_ASAP7_75t_L g2745 ( 
.A1(n_2493),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2215),
.B(n_40),
.Y(n_2746)
);

OAI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2415),
.A2(n_2211),
.B(n_2210),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2352),
.B(n_41),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2353),
.Y(n_2749)
);

AO21x1_ASAP7_75t_L g2750 ( 
.A1(n_2478),
.A2(n_529),
.B(n_528),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2344),
.A2(n_2281),
.B(n_2317),
.Y(n_2751)
);

OAI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2526),
.A2(n_42),
.B(n_43),
.Y(n_2752)
);

NAND3xp33_ASAP7_75t_L g2753 ( 
.A(n_2313),
.B(n_43),
.C(n_44),
.Y(n_2753)
);

OAI21xp5_ASAP7_75t_L g2754 ( 
.A1(n_2528),
.A2(n_43),
.B(n_44),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2295),
.B(n_45),
.Y(n_2755)
);

OAI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2542),
.A2(n_45),
.B(n_46),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2433),
.B(n_46),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2280),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2758)
);

AND2x4_ASAP7_75t_SL g2759 ( 
.A(n_2312),
.B(n_47),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2520),
.B(n_48),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2349),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2305),
.B(n_47),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2433),
.B(n_49),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2308),
.B(n_49),
.Y(n_2764)
);

INVx3_ASAP7_75t_L g2765 ( 
.A(n_2217),
.Y(n_2765)
);

BUFx6f_ASAP7_75t_L g2766 ( 
.A(n_2217),
.Y(n_2766)
);

BUFx4f_ASAP7_75t_L g2767 ( 
.A(n_2399),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2227),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2331),
.A2(n_50),
.B(n_51),
.Y(n_2769)
);

A2O1A1Ixp33_ASAP7_75t_L g2770 ( 
.A1(n_2296),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2226),
.B(n_52),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2227),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2341),
.A2(n_53),
.B(n_54),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_SL g2774 ( 
.A(n_2547),
.B(n_54),
.Y(n_2774)
);

NAND2x1p5_ASAP7_75t_L g2775 ( 
.A(n_2263),
.B(n_53),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2234),
.B(n_53),
.Y(n_2776)
);

OAI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2560),
.A2(n_54),
.B(n_55),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2420),
.A2(n_55),
.B(n_56),
.Y(n_2778)
);

INVx1_ASAP7_75t_SL g2779 ( 
.A(n_2222),
.Y(n_2779)
);

O2A1O1Ixp33_ASAP7_75t_L g2780 ( 
.A1(n_2428),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_2780)
);

AOI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2333),
.A2(n_57),
.B(n_58),
.Y(n_2781)
);

AOI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2335),
.A2(n_57),
.B(n_58),
.Y(n_2782)
);

AOI21x1_ASAP7_75t_L g2783 ( 
.A1(n_2579),
.A2(n_59),
.B(n_60),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2300),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2354),
.B(n_2319),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2319),
.Y(n_2786)
);

AOI21xp5_ASAP7_75t_L g2787 ( 
.A1(n_2339),
.A2(n_61),
.B(n_62),
.Y(n_2787)
);

INVx4_ASAP7_75t_L g2788 ( 
.A(n_2262),
.Y(n_2788)
);

AO21x1_ASAP7_75t_L g2789 ( 
.A1(n_2531),
.A2(n_529),
.B(n_528),
.Y(n_2789)
);

AOI21xp5_ASAP7_75t_L g2790 ( 
.A1(n_2358),
.A2(n_62),
.B(n_63),
.Y(n_2790)
);

NOR3xp33_ASAP7_75t_L g2791 ( 
.A(n_2564),
.B(n_64),
.C(n_63),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2559),
.B(n_63),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2364),
.A2(n_62),
.B(n_64),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2367),
.A2(n_64),
.B(n_65),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2407),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2342),
.B(n_65),
.Y(n_2796)
);

NOR2x2_ASAP7_75t_L g2797 ( 
.A(n_2399),
.B(n_66),
.Y(n_2797)
);

AOI21xp5_ASAP7_75t_L g2798 ( 
.A1(n_2374),
.A2(n_66),
.B(n_67),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2572),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_L g2800 ( 
.A(n_2312),
.B(n_67),
.Y(n_2800)
);

OAI21xp5_ASAP7_75t_L g2801 ( 
.A1(n_2574),
.A2(n_68),
.B(n_69),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_SL g2802 ( 
.A(n_2561),
.B(n_69),
.Y(n_2802)
);

A2O1A1Ixp33_ASAP7_75t_L g2803 ( 
.A1(n_2347),
.A2(n_71),
.B(n_68),
.C(n_70),
.Y(n_2803)
);

AOI222xp33_ASAP7_75t_L g2804 ( 
.A1(n_2460),
.A2(n_71),
.B1(n_73),
.B2(n_68),
.C1(n_70),
.C2(n_72),
.Y(n_2804)
);

O2A1O1Ixp33_ASAP7_75t_L g2805 ( 
.A1(n_2445),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2429),
.Y(n_2806)
);

NAND2x1p5_ASAP7_75t_L g2807 ( 
.A(n_2271),
.B(n_72),
.Y(n_2807)
);

INVx4_ASAP7_75t_L g2808 ( 
.A(n_2227),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2406),
.B(n_74),
.Y(n_2809)
);

BUFx6f_ASAP7_75t_L g2810 ( 
.A(n_2535),
.Y(n_2810)
);

AOI21xp5_ASAP7_75t_L g2811 ( 
.A1(n_2376),
.A2(n_73),
.B(n_74),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2441),
.B(n_75),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2446),
.Y(n_2813)
);

A2O1A1Ixp33_ASAP7_75t_L g2814 ( 
.A1(n_2338),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_2814)
);

NOR2xp67_ASAP7_75t_L g2815 ( 
.A(n_2413),
.B(n_75),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2379),
.A2(n_76),
.B(n_77),
.Y(n_2816)
);

A2O1A1Ixp33_ASAP7_75t_L g2817 ( 
.A1(n_2378),
.A2(n_79),
.B(n_76),
.C(n_78),
.Y(n_2817)
);

BUFx6f_ASAP7_75t_L g2818 ( 
.A(n_2535),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2330),
.B(n_78),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2229),
.B(n_2307),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2411),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2250),
.B(n_78),
.Y(n_2822)
);

INVxp67_ASAP7_75t_L g2823 ( 
.A(n_2266),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2385),
.A2(n_79),
.B(n_80),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2389),
.A2(n_80),
.B(n_81),
.Y(n_2825)
);

AOI21xp5_ASAP7_75t_L g2826 ( 
.A1(n_2390),
.A2(n_80),
.B(n_81),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2270),
.B(n_2535),
.Y(n_2827)
);

BUFx6f_ASAP7_75t_L g2828 ( 
.A(n_2418),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2392),
.B(n_81),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2423),
.B(n_83),
.Y(n_2830)
);

A2O1A1Ixp33_ASAP7_75t_L g2831 ( 
.A1(n_2451),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2488),
.A2(n_82),
.B(n_83),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2366),
.B(n_82),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2418),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2359),
.B(n_84),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2494),
.A2(n_2495),
.B(n_2249),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2239),
.A2(n_2447),
.B(n_2417),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2370),
.B(n_84),
.Y(n_2838)
);

CKINVDCx16_ASAP7_75t_R g2839 ( 
.A(n_2432),
.Y(n_2839)
);

BUFx6f_ASAP7_75t_L g2840 ( 
.A(n_2418),
.Y(n_2840)
);

AOI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2454),
.A2(n_85),
.B(n_86),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_SL g2842 ( 
.A(n_2440),
.B(n_87),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2310),
.Y(n_2843)
);

AOI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_2455),
.A2(n_86),
.B(n_87),
.Y(n_2844)
);

NOR2x1_ASAP7_75t_L g2845 ( 
.A(n_2336),
.B(n_86),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2549),
.B(n_88),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2318),
.Y(n_2847)
);

OAI21xp5_ASAP7_75t_L g2848 ( 
.A1(n_2456),
.A2(n_88),
.B(n_89),
.Y(n_2848)
);

CKINVDCx11_ASAP7_75t_R g2849 ( 
.A(n_2431),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2361),
.B(n_2315),
.Y(n_2850)
);

BUFx12f_ASAP7_75t_L g2851 ( 
.A(n_2373),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2461),
.B(n_88),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2457),
.A2(n_90),
.B(n_91),
.Y(n_2853)
);

AOI21xp33_ASAP7_75t_L g2854 ( 
.A1(n_2414),
.A2(n_90),
.B(n_91),
.Y(n_2854)
);

BUFx4f_ASAP7_75t_L g2855 ( 
.A(n_2369),
.Y(n_2855)
);

AOI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2463),
.A2(n_2466),
.B(n_2490),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2396),
.B(n_91),
.Y(n_2857)
);

AOI21xp33_ASAP7_75t_L g2858 ( 
.A1(n_2324),
.A2(n_90),
.B(n_92),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2426),
.A2(n_2419),
.B1(n_2540),
.B2(n_2309),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2360),
.B(n_92),
.Y(n_2860)
);

OAI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2408),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_2861)
);

OAI21xp33_ASAP7_75t_L g2862 ( 
.A1(n_2443),
.A2(n_93),
.B(n_94),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2550),
.B(n_93),
.Y(n_2863)
);

O2A1O1Ixp33_ASAP7_75t_L g2864 ( 
.A1(n_2273),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2205),
.B(n_96),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2507),
.B(n_96),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2387),
.Y(n_2867)
);

AOI21x1_ASAP7_75t_L g2868 ( 
.A1(n_2577),
.A2(n_97),
.B(n_99),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2425),
.B(n_100),
.Y(n_2869)
);

AOI21xp5_ASAP7_75t_L g2870 ( 
.A1(n_2496),
.A2(n_99),
.B(n_100),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2508),
.A2(n_100),
.B(n_101),
.Y(n_2871)
);

INVx4_ASAP7_75t_L g2872 ( 
.A(n_2413),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2444),
.A2(n_101),
.B(n_102),
.Y(n_2873)
);

INVx3_ASAP7_75t_L g2874 ( 
.A(n_2387),
.Y(n_2874)
);

OAI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2351),
.A2(n_101),
.B(n_102),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2404),
.Y(n_2876)
);

CKINVDCx8_ASAP7_75t_R g2877 ( 
.A(n_2491),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2404),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2449),
.A2(n_103),
.B(n_104),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2503),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2430),
.B(n_103),
.Y(n_2881)
);

AOI21xp5_ASAP7_75t_L g2882 ( 
.A1(n_2464),
.A2(n_2468),
.B(n_2465),
.Y(n_2882)
);

AOI21x1_ASAP7_75t_L g2883 ( 
.A1(n_2571),
.A2(n_103),
.B(n_104),
.Y(n_2883)
);

O2A1O1Ixp33_ASAP7_75t_L g2884 ( 
.A1(n_2274),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2503),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2516),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2391),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2377),
.B(n_105),
.Y(n_2888)
);

NOR2x1_ASAP7_75t_L g2889 ( 
.A(n_2381),
.B(n_105),
.Y(n_2889)
);

INVx2_ASAP7_75t_SL g2890 ( 
.A(n_2506),
.Y(n_2890)
);

O2A1O1Ixp5_ASAP7_75t_L g2891 ( 
.A1(n_2236),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2891)
);

O2A1O1Ixp33_ASAP7_75t_L g2892 ( 
.A1(n_2462),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2500),
.B(n_108),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_SL g2894 ( 
.A(n_2427),
.B(n_110),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_L g2895 ( 
.A(n_2551),
.B(n_109),
.Y(n_2895)
);

AND2x2_ASAP7_75t_SL g2896 ( 
.A(n_2479),
.B(n_110),
.Y(n_2896)
);

OAI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2368),
.A2(n_2509),
.B(n_2502),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2261),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2474),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2219),
.B(n_110),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2469),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2476),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2321),
.B(n_111),
.Y(n_2903)
);

HB1xp67_ASAP7_75t_L g2904 ( 
.A(n_2519),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2480),
.A2(n_2435),
.B(n_2442),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2472),
.A2(n_111),
.B(n_112),
.Y(n_2906)
);

OAI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2501),
.A2(n_111),
.B(n_113),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2475),
.Y(n_2908)
);

OAI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2481),
.A2(n_2450),
.B(n_2458),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2261),
.Y(n_2910)
);

HB1xp67_ASAP7_75t_L g2911 ( 
.A(n_2521),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2409),
.B(n_113),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2483),
.A2(n_114),
.B(n_115),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2523),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2522),
.A2(n_114),
.B(n_115),
.Y(n_2915)
);

O2A1O1Ixp5_ASAP7_75t_L g2916 ( 
.A1(n_2436),
.A2(n_119),
.B(n_116),
.C(n_117),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2482),
.A2(n_116),
.B(n_117),
.Y(n_2917)
);

NOR2xp67_ASAP7_75t_L g2918 ( 
.A(n_2499),
.B(n_119),
.Y(n_2918)
);

AOI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2242),
.A2(n_119),
.B(n_120),
.Y(n_2919)
);

AOI21x1_ASAP7_75t_L g2920 ( 
.A1(n_2505),
.A2(n_120),
.B(n_121),
.Y(n_2920)
);

AOI21xp33_ASAP7_75t_L g2921 ( 
.A1(n_2448),
.A2(n_120),
.B(n_121),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2439),
.B(n_121),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2452),
.B(n_122),
.Y(n_2923)
);

AOI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2485),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2513),
.B(n_122),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2384),
.B(n_123),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2386),
.B(n_123),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2302),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_SL g2929 ( 
.A(n_2484),
.B(n_125),
.Y(n_2929)
);

OAI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2492),
.A2(n_124),
.B(n_125),
.Y(n_2930)
);

AO21x2_ASAP7_75t_L g2931 ( 
.A1(n_2418),
.A2(n_2486),
.B(n_2394),
.Y(n_2931)
);

NOR3xp33_ASAP7_75t_L g2932 ( 
.A(n_2279),
.B(n_127),
.C(n_126),
.Y(n_2932)
);

OAI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2497),
.A2(n_124),
.B(n_126),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2498),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_2934)
);

AO22x1_ASAP7_75t_L g2935 ( 
.A1(n_2517),
.A2(n_130),
.B1(n_131),
.B2(n_129),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2393),
.B(n_128),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2525),
.B(n_130),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2395),
.A2(n_128),
.B(n_130),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2371),
.Y(n_2939)
);

AND2x4_ASAP7_75t_L g2940 ( 
.A(n_2398),
.B(n_131),
.Y(n_2940)
);

AND2x4_ASAP7_75t_L g2941 ( 
.A(n_2402),
.B(n_131),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_SL g2942 ( 
.A(n_2515),
.B(n_132),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2405),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2416),
.B(n_132),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2473),
.B(n_2511),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2471),
.B(n_133),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2302),
.A2(n_134),
.B(n_135),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2471),
.B(n_134),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2512),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2514),
.B(n_134),
.Y(n_2950)
);

INVx4_ASAP7_75t_L g2951 ( 
.A(n_2262),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2372),
.Y(n_2952)
);

NOR3xp33_ASAP7_75t_L g2953 ( 
.A(n_2280),
.B(n_137),
.C(n_136),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2289),
.Y(n_2954)
);

OAI321xp33_ASAP7_75t_L g2955 ( 
.A1(n_2280),
.A2(n_137),
.A3(n_139),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2380),
.A2(n_136),
.B(n_138),
.Y(n_2956)
);

OAI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2477),
.A2(n_138),
.B(n_139),
.Y(n_2957)
);

A2O1A1Ixp33_ASAP7_75t_L g2958 ( 
.A1(n_2346),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_2958)
);

AOI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2380),
.A2(n_140),
.B(n_142),
.Y(n_2959)
);

AOI21x1_ASAP7_75t_L g2960 ( 
.A1(n_2489),
.A2(n_140),
.B(n_142),
.Y(n_2960)
);

AOI21x1_ASAP7_75t_L g2961 ( 
.A1(n_2489),
.A2(n_142),
.B(n_143),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_2397),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2289),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2372),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2230),
.A2(n_146),
.B1(n_143),
.B2(n_145),
.Y(n_2965)
);

A2O1A1Ixp33_ASAP7_75t_L g2966 ( 
.A1(n_2346),
.A2(n_146),
.B(n_143),
.C(n_145),
.Y(n_2966)
);

INVx2_ASAP7_75t_SL g2967 ( 
.A(n_2263),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2372),
.Y(n_2968)
);

AOI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2230),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_2969)
);

AOI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2380),
.A2(n_147),
.B(n_148),
.Y(n_2970)
);

BUFx6f_ASAP7_75t_L g2971 ( 
.A(n_2397),
.Y(n_2971)
);

INVx2_ASAP7_75t_SL g2972 ( 
.A(n_2263),
.Y(n_2972)
);

OAI21xp33_ASAP7_75t_L g2973 ( 
.A1(n_2327),
.A2(n_147),
.B(n_148),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2327),
.B(n_149),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2212),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_2975)
);

AOI21xp5_ASAP7_75t_L g2976 ( 
.A1(n_2380),
.A2(n_149),
.B(n_151),
.Y(n_2976)
);

BUFx6f_ASAP7_75t_L g2977 ( 
.A(n_2397),
.Y(n_2977)
);

O2A1O1Ixp5_ASAP7_75t_L g2978 ( 
.A1(n_2569),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2212),
.B(n_152),
.Y(n_2979)
);

AOI22xp5_ASAP7_75t_L g2980 ( 
.A1(n_2230),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2980)
);

AOI22xp33_ASAP7_75t_L g2981 ( 
.A1(n_2223),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_2981)
);

NOR3xp33_ASAP7_75t_L g2982 ( 
.A(n_2280),
.B(n_157),
.C(n_156),
.Y(n_2982)
);

O2A1O1Ixp33_ASAP7_75t_L g2983 ( 
.A1(n_2569),
.A2(n_158),
.B(n_155),
.C(n_157),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_L g2984 ( 
.A(n_2327),
.B(n_158),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2212),
.B(n_159),
.Y(n_2985)
);

AOI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2380),
.A2(n_159),
.B(n_160),
.Y(n_2986)
);

AOI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2380),
.A2(n_159),
.B(n_161),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_L g2988 ( 
.A(n_2327),
.B(n_161),
.Y(n_2988)
);

HB1xp67_ASAP7_75t_L g2989 ( 
.A(n_2546),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_SL g2990 ( 
.A(n_2546),
.B(n_162),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_L g2991 ( 
.A(n_2327),
.B(n_161),
.Y(n_2991)
);

AOI21xp5_ASAP7_75t_L g2992 ( 
.A1(n_2380),
.A2(n_162),
.B(n_163),
.Y(n_2992)
);

NOR2xp33_ASAP7_75t_L g2993 ( 
.A(n_2327),
.B(n_162),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_SL g2994 ( 
.A(n_2546),
.B(n_164),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2372),
.Y(n_2995)
);

OAI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2477),
.A2(n_163),
.B(n_164),
.Y(n_2996)
);

AOI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2380),
.A2(n_163),
.B(n_164),
.Y(n_2997)
);

AOI21xp5_ASAP7_75t_L g2998 ( 
.A1(n_2380),
.A2(n_165),
.B(n_166),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2204),
.B(n_165),
.Y(n_2999)
);

AOI21xp5_ASAP7_75t_L g3000 ( 
.A1(n_2380),
.A2(n_165),
.B(n_166),
.Y(n_3000)
);

AOI21x1_ASAP7_75t_L g3001 ( 
.A1(n_2489),
.A2(n_166),
.B(n_167),
.Y(n_3001)
);

HB1xp67_ASAP7_75t_L g3002 ( 
.A(n_2546),
.Y(n_3002)
);

INVx2_ASAP7_75t_SL g3003 ( 
.A(n_2263),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2546),
.B(n_168),
.Y(n_3004)
);

NOR3xp33_ASAP7_75t_L g3005 ( 
.A(n_2280),
.B(n_170),
.C(n_169),
.Y(n_3005)
);

BUFx3_ASAP7_75t_L g3006 ( 
.A(n_2252),
.Y(n_3006)
);

AOI22xp5_ASAP7_75t_L g3007 ( 
.A1(n_2230),
.A2(n_170),
.B1(n_167),
.B2(n_169),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2289),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2372),
.Y(n_3009)
);

O2A1O1Ixp5_ASAP7_75t_L g3010 ( 
.A1(n_2569),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_3010)
);

AOI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2380),
.A2(n_171),
.B(n_172),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2289),
.B(n_172),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2326),
.Y(n_3013)
);

BUFx6f_ASAP7_75t_L g3014 ( 
.A(n_2397),
.Y(n_3014)
);

OAI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2477),
.A2(n_172),
.B(n_173),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2372),
.Y(n_3016)
);

O2A1O1Ixp33_ASAP7_75t_L g3017 ( 
.A1(n_2569),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2212),
.B(n_175),
.Y(n_3018)
);

OAI21xp5_ASAP7_75t_L g3019 ( 
.A1(n_2477),
.A2(n_176),
.B(n_177),
.Y(n_3019)
);

AOI21x1_ASAP7_75t_L g3020 ( 
.A1(n_2489),
.A2(n_176),
.B(n_177),
.Y(n_3020)
);

OAI321xp33_ASAP7_75t_L g3021 ( 
.A1(n_2280),
.A2(n_178),
.A3(n_180),
.B1(n_176),
.B2(n_177),
.C(n_179),
.Y(n_3021)
);

INVx3_ASAP7_75t_L g3022 ( 
.A(n_2557),
.Y(n_3022)
);

BUFx6f_ASAP7_75t_L g3023 ( 
.A(n_2397),
.Y(n_3023)
);

AOI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2380),
.A2(n_178),
.B(n_179),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2212),
.B(n_178),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2372),
.Y(n_3026)
);

NOR2xp33_ASAP7_75t_SL g3027 ( 
.A(n_2230),
.B(n_179),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2212),
.B(n_180),
.Y(n_3028)
);

O2A1O1Ixp33_ASAP7_75t_L g3029 ( 
.A1(n_2569),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2212),
.B(n_181),
.Y(n_3030)
);

AOI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2380),
.A2(n_181),
.B(n_182),
.Y(n_3031)
);

AOI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2380),
.A2(n_183),
.B(n_184),
.Y(n_3032)
);

AOI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2230),
.A2(n_186),
.B1(n_183),
.B2(n_184),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2372),
.Y(n_3034)
);

AOI21xp5_ASAP7_75t_L g3035 ( 
.A1(n_2380),
.A2(n_183),
.B(n_184),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2372),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2212),
.B(n_186),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2212),
.B(n_187),
.Y(n_3038)
);

OR2x6_ASAP7_75t_L g3039 ( 
.A(n_2216),
.B(n_187),
.Y(n_3039)
);

INVx3_ASAP7_75t_L g3040 ( 
.A(n_2557),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_2546),
.B(n_189),
.Y(n_3041)
);

A2O1A1Ixp33_ASAP7_75t_L g3042 ( 
.A1(n_2346),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2212),
.B(n_188),
.Y(n_3043)
);

OAI21xp33_ASAP7_75t_L g3044 ( 
.A1(n_2327),
.A2(n_188),
.B(n_190),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2212),
.B(n_190),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2289),
.Y(n_3046)
);

OAI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2477),
.A2(n_191),
.B(n_192),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2212),
.B(n_191),
.Y(n_3048)
);

AOI21xp33_ASAP7_75t_L g3049 ( 
.A1(n_2327),
.A2(n_191),
.B(n_192),
.Y(n_3049)
);

AOI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2380),
.A2(n_192),
.B(n_193),
.Y(n_3050)
);

BUFx6f_ASAP7_75t_L g3051 ( 
.A(n_2397),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2212),
.B(n_193),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2546),
.B(n_194),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2327),
.B(n_193),
.Y(n_3054)
);

AO21x1_ASAP7_75t_L g3055 ( 
.A1(n_2489),
.A2(n_533),
.B(n_531),
.Y(n_3055)
);

NOR3xp33_ASAP7_75t_L g3056 ( 
.A(n_2280),
.B(n_196),
.C(n_195),
.Y(n_3056)
);

INVx3_ASAP7_75t_L g3057 ( 
.A(n_2557),
.Y(n_3057)
);

NOR2xp67_ASAP7_75t_L g3058 ( 
.A(n_2413),
.B(n_194),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2212),
.B(n_194),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2212),
.B(n_195),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_L g3061 ( 
.A(n_2327),
.B(n_196),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2289),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2380),
.A2(n_196),
.B(n_197),
.Y(n_3063)
);

AOI21x1_ASAP7_75t_L g3064 ( 
.A1(n_2489),
.A2(n_197),
.B(n_198),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2212),
.B(n_197),
.Y(n_3065)
);

BUFx6f_ASAP7_75t_SL g3066 ( 
.A(n_2216),
.Y(n_3066)
);

HB1xp67_ASAP7_75t_L g3067 ( 
.A(n_2546),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2289),
.Y(n_3068)
);

OAI21xp33_ASAP7_75t_L g3069 ( 
.A1(n_2327),
.A2(n_198),
.B(n_199),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_L g3070 ( 
.A(n_2327),
.B(n_198),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2289),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2289),
.Y(n_3072)
);

AOI21xp5_ASAP7_75t_L g3073 ( 
.A1(n_2380),
.A2(n_199),
.B(n_200),
.Y(n_3073)
);

BUFx4f_ASAP7_75t_L g3074 ( 
.A(n_2326),
.Y(n_3074)
);

OA21x2_ASAP7_75t_L g3075 ( 
.A1(n_2489),
.A2(n_199),
.B(n_200),
.Y(n_3075)
);

OAI21xp33_ASAP7_75t_L g3076 ( 
.A1(n_2327),
.A2(n_200),
.B(n_201),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2327),
.B(n_201),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2212),
.B(n_201),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2212),
.B(n_202),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2212),
.B(n_202),
.Y(n_3080)
);

O2A1O1Ixp33_ASAP7_75t_L g3081 ( 
.A1(n_2569),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2212),
.B(n_203),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2212),
.B(n_203),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2212),
.B(n_204),
.Y(n_3084)
);

A2O1A1Ixp33_ASAP7_75t_L g3085 ( 
.A1(n_2346),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_3085)
);

AOI21xp5_ASAP7_75t_L g3086 ( 
.A1(n_2380),
.A2(n_205),
.B(n_206),
.Y(n_3086)
);

HB1xp67_ASAP7_75t_L g3087 ( 
.A(n_2546),
.Y(n_3087)
);

OAI21xp33_ASAP7_75t_L g3088 ( 
.A1(n_2327),
.A2(n_205),
.B(n_206),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2372),
.Y(n_3089)
);

BUFx4f_ASAP7_75t_L g3090 ( 
.A(n_2326),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2212),
.B(n_207),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2380),
.A2(n_207),
.B(n_208),
.Y(n_3092)
);

INVxp67_ASAP7_75t_L g3093 ( 
.A(n_2230),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2212),
.B(n_209),
.Y(n_3094)
);

BUFx6f_ASAP7_75t_L g3095 ( 
.A(n_2397),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2327),
.B(n_209),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2289),
.Y(n_3097)
);

AOI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_2380),
.A2(n_210),
.B(n_211),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2289),
.Y(n_3099)
);

NOR2xp33_ASAP7_75t_L g3100 ( 
.A(n_2327),
.B(n_210),
.Y(n_3100)
);

NAND2x1p5_ASAP7_75t_L g3101 ( 
.A(n_2263),
.B(n_210),
.Y(n_3101)
);

AOI33xp33_ASAP7_75t_L g3102 ( 
.A1(n_2311),
.A2(n_213),
.A3(n_215),
.B1(n_211),
.B2(n_212),
.B3(n_214),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2212),
.B(n_212),
.Y(n_3103)
);

INVxp67_ASAP7_75t_L g3104 ( 
.A(n_2230),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2380),
.A2(n_212),
.B(n_213),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2380),
.A2(n_213),
.B(n_215),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2212),
.B(n_215),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2380),
.A2(n_216),
.B(n_217),
.Y(n_3108)
);

AOI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2380),
.A2(n_216),
.B(n_217),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2380),
.A2(n_216),
.B(n_217),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2212),
.B(n_218),
.Y(n_3111)
);

BUFx12f_ASAP7_75t_L g3112 ( 
.A(n_2326),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2372),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2212),
.B(n_218),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2380),
.A2(n_218),
.B(n_219),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2212),
.B(n_219),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2546),
.B(n_220),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2380),
.A2(n_219),
.B(n_220),
.Y(n_3118)
);

NAND3xp33_ASAP7_75t_L g3119 ( 
.A(n_2412),
.B(n_221),
.C(n_222),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2289),
.Y(n_3120)
);

NAND2x1_ASAP7_75t_L g3121 ( 
.A(n_2397),
.B(n_221),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2289),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2546),
.B(n_222),
.Y(n_3123)
);

HB1xp67_ASAP7_75t_L g3124 ( 
.A(n_2546),
.Y(n_3124)
);

OAI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_2477),
.A2(n_221),
.B(n_222),
.Y(n_3125)
);

AOI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2380),
.A2(n_223),
.B(n_224),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2380),
.A2(n_223),
.B(n_224),
.Y(n_3127)
);

O2A1O1Ixp5_ASAP7_75t_L g3128 ( 
.A1(n_2569),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2212),
.B(n_225),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2212),
.B(n_225),
.Y(n_3130)
);

AO21x1_ASAP7_75t_L g3131 ( 
.A1(n_2489),
.A2(n_533),
.B(n_531),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2212),
.B(n_226),
.Y(n_3132)
);

AOI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_2380),
.A2(n_226),
.B(n_227),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2372),
.Y(n_3134)
);

CKINVDCx10_ASAP7_75t_R g3135 ( 
.A(n_2216),
.Y(n_3135)
);

AOI21x1_ASAP7_75t_L g3136 ( 
.A1(n_2489),
.A2(n_227),
.B(n_228),
.Y(n_3136)
);

OAI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_2477),
.A2(n_228),
.B(n_229),
.Y(n_3137)
);

NOR2xp33_ASAP7_75t_L g3138 ( 
.A(n_2327),
.B(n_228),
.Y(n_3138)
);

NOR2xp67_ASAP7_75t_L g3139 ( 
.A(n_2413),
.B(n_229),
.Y(n_3139)
);

AOI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_2380),
.A2(n_229),
.B(n_230),
.Y(n_3140)
);

OAI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2477),
.A2(n_230),
.B(n_231),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_SL g3142 ( 
.A(n_2546),
.B(n_232),
.Y(n_3142)
);

INVxp67_ASAP7_75t_L g3143 ( 
.A(n_2230),
.Y(n_3143)
);

AOI21xp5_ASAP7_75t_L g3144 ( 
.A1(n_2380),
.A2(n_230),
.B(n_232),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2372),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2289),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2557),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2212),
.B(n_232),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_2327),
.B(n_233),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2372),
.Y(n_3150)
);

OAI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_2212),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2372),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_2380),
.A2(n_233),
.B(n_234),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_2204),
.B(n_234),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2212),
.B(n_236),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_2380),
.A2(n_236),
.B(n_237),
.Y(n_3156)
);

OR2x2_ASAP7_75t_L g3157 ( 
.A(n_2258),
.B(n_237),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2380),
.A2(n_237),
.B(n_238),
.Y(n_3158)
);

OAI22xp5_ASAP7_75t_L g3159 ( 
.A1(n_2212),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_3159)
);

INVx3_ASAP7_75t_L g3160 ( 
.A(n_2557),
.Y(n_3160)
);

OAI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_2212),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_3161)
);

NOR2xp33_ASAP7_75t_L g3162 ( 
.A(n_2327),
.B(n_239),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2380),
.A2(n_240),
.B(n_241),
.Y(n_3163)
);

AOI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_2380),
.A2(n_242),
.B(n_243),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2212),
.B(n_242),
.Y(n_3165)
);

NOR2x1_ASAP7_75t_L g3166 ( 
.A(n_2252),
.B(n_242),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2212),
.B(n_243),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2380),
.A2(n_244),
.B(n_245),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_SL g3169 ( 
.A(n_2546),
.B(n_245),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2212),
.B(n_244),
.Y(n_3170)
);

AOI21xp33_ASAP7_75t_L g3171 ( 
.A1(n_2327),
.A2(n_244),
.B(n_245),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2546),
.B(n_247),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2289),
.Y(n_3173)
);

OAI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_2212),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_3174)
);

OAI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_2477),
.A2(n_246),
.B(n_247),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2212),
.B(n_248),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2289),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2380),
.A2(n_248),
.B(n_249),
.Y(n_3178)
);

BUFx6f_ASAP7_75t_L g3179 ( 
.A(n_2397),
.Y(n_3179)
);

OAI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2477),
.A2(n_249),
.B(n_250),
.Y(n_3180)
);

HB1xp67_ASAP7_75t_L g3181 ( 
.A(n_2546),
.Y(n_3181)
);

OAI21xp5_ASAP7_75t_L g3182 ( 
.A1(n_2477),
.A2(n_250),
.B(n_251),
.Y(n_3182)
);

A2O1A1Ixp33_ASAP7_75t_L g3183 ( 
.A1(n_2346),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2380),
.A2(n_251),
.B(n_252),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2380),
.A2(n_252),
.B(n_253),
.Y(n_3185)
);

AO21x1_ASAP7_75t_L g3186 ( 
.A1(n_2489),
.A2(n_535),
.B(n_534),
.Y(n_3186)
);

NOR2x1_ASAP7_75t_R g3187 ( 
.A(n_2262),
.B(n_254),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2212),
.B(n_254),
.Y(n_3188)
);

O2A1O1Ixp33_ASAP7_75t_L g3189 ( 
.A1(n_2569),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2212),
.B(n_255),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_2204),
.B(n_256),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2212),
.B(n_256),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2212),
.B(n_258),
.Y(n_3193)
);

NOR2xp33_ASAP7_75t_SL g3194 ( 
.A(n_2230),
.B(n_258),
.Y(n_3194)
);

BUFx2_ASAP7_75t_L g3195 ( 
.A(n_2546),
.Y(n_3195)
);

OAI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_2477),
.A2(n_259),
.B(n_260),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2372),
.Y(n_3197)
);

O2A1O1Ixp33_ASAP7_75t_L g3198 ( 
.A1(n_2569),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_3198)
);

INVx3_ASAP7_75t_L g3199 ( 
.A(n_2557),
.Y(n_3199)
);

OAI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_2477),
.A2(n_259),
.B(n_260),
.Y(n_3200)
);

A2O1A1Ixp33_ASAP7_75t_L g3201 ( 
.A1(n_2346),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2289),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2212),
.B(n_262),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2289),
.Y(n_3204)
);

OAI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_2477),
.A2(n_262),
.B(n_263),
.Y(n_3205)
);

OR2x2_ASAP7_75t_L g3206 ( 
.A(n_2258),
.B(n_263),
.Y(n_3206)
);

OAI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_2212),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_3207)
);

AOI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_2380),
.A2(n_264),
.B(n_265),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2212),
.B(n_264),
.Y(n_3209)
);

INVx2_ASAP7_75t_L g3210 ( 
.A(n_2372),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2372),
.Y(n_3211)
);

A2O1A1Ixp33_ASAP7_75t_L g3212 ( 
.A1(n_2346),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_3212)
);

OR2x6_ASAP7_75t_L g3213 ( 
.A(n_2216),
.B(n_266),
.Y(n_3213)
);

AOI21xp5_ASAP7_75t_L g3214 ( 
.A1(n_2380),
.A2(n_267),
.B(n_268),
.Y(n_3214)
);

AOI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2380),
.A2(n_267),
.B(n_268),
.Y(n_3215)
);

A2O1A1Ixp33_ASAP7_75t_L g3216 ( 
.A1(n_2346),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_3216)
);

INVxp67_ASAP7_75t_L g3217 ( 
.A(n_2230),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2327),
.B(n_269),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2289),
.Y(n_3219)
);

BUFx3_ASAP7_75t_L g3220 ( 
.A(n_3074),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2859),
.B(n_270),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_SL g3222 ( 
.A(n_2855),
.B(n_270),
.Y(n_3222)
);

AOI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_2595),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_3223)
);

AOI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_2645),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_2767),
.B(n_534),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_L g3226 ( 
.A(n_2584),
.Y(n_3226)
);

CKINVDCx5p33_ASAP7_75t_R g3227 ( 
.A(n_2849),
.Y(n_3227)
);

OAI21xp33_ASAP7_75t_L g3228 ( 
.A1(n_3027),
.A2(n_273),
.B(n_274),
.Y(n_3228)
);

CKINVDCx5p33_ASAP7_75t_R g3229 ( 
.A(n_2629),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2648),
.B(n_275),
.Y(n_3230)
);

O2A1O1Ixp33_ASAP7_75t_L g3231 ( 
.A1(n_2671),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2620),
.B(n_277),
.Y(n_3232)
);

OR2x6_ASAP7_75t_SL g3233 ( 
.A(n_2731),
.B(n_277),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2590),
.Y(n_3234)
);

INVxp67_ASAP7_75t_SL g3235 ( 
.A(n_2989),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_SL g3236 ( 
.A(n_2767),
.B(n_535),
.Y(n_3236)
);

INVx2_ASAP7_75t_SL g3237 ( 
.A(n_2855),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2601),
.Y(n_3238)
);

O2A1O1Ixp33_ASAP7_75t_L g3239 ( 
.A1(n_2715),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_SL g3240 ( 
.A(n_3194),
.B(n_536),
.Y(n_3240)
);

CKINVDCx5p33_ASAP7_75t_R g3241 ( 
.A(n_3135),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2616),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2596),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_L g3244 ( 
.A(n_2692),
.B(n_278),
.Y(n_3244)
);

CKINVDCx11_ASAP7_75t_R g3245 ( 
.A(n_3112),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2620),
.B(n_279),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2581),
.Y(n_3247)
);

O2A1O1Ixp33_ASAP7_75t_L g3248 ( 
.A1(n_2735),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2886),
.B(n_280),
.Y(n_3249)
);

BUFx4f_ASAP7_75t_SL g3250 ( 
.A(n_2600),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2606),
.B(n_281),
.Y(n_3251)
);

OAI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_3039),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3252)
);

HB1xp67_ASAP7_75t_L g3253 ( 
.A(n_3195),
.Y(n_3253)
);

BUFx3_ASAP7_75t_L g3254 ( 
.A(n_3074),
.Y(n_3254)
);

BUFx3_ASAP7_75t_L g3255 ( 
.A(n_3090),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2839),
.B(n_282),
.Y(n_3256)
);

O2A1O1Ixp5_ASAP7_75t_L g3257 ( 
.A1(n_2957),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_3257)
);

INVx2_ASAP7_75t_SL g3258 ( 
.A(n_3090),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2609),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_L g3260 ( 
.A(n_2584),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_3093),
.B(n_536),
.Y(n_3261)
);

NOR3xp33_ASAP7_75t_SL g3262 ( 
.A(n_3013),
.B(n_2843),
.C(n_2955),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2633),
.Y(n_3263)
);

AOI21xp33_ASAP7_75t_L g3264 ( 
.A1(n_2923),
.A2(n_283),
.B(n_284),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2952),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_2584),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2954),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2963),
.B(n_284),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_L g3269 ( 
.A(n_2823),
.B(n_285),
.Y(n_3269)
);

CKINVDCx8_ASAP7_75t_R g3270 ( 
.A(n_3039),
.Y(n_3270)
);

BUFx2_ASAP7_75t_L g3271 ( 
.A(n_3039),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2964),
.Y(n_3272)
);

INVx6_ASAP7_75t_L g3273 ( 
.A(n_2722),
.Y(n_3273)
);

INVx3_ASAP7_75t_L g3274 ( 
.A(n_2872),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3008),
.Y(n_3275)
);

INVx3_ASAP7_75t_L g3276 ( 
.A(n_2872),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_2896),
.B(n_285),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3046),
.Y(n_3278)
);

AOI22xp33_ASAP7_75t_L g3279 ( 
.A1(n_3213),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_2882),
.A2(n_287),
.B(n_288),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3062),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_2658),
.A2(n_287),
.B(n_288),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2682),
.B(n_289),
.Y(n_3283)
);

O2A1O1Ixp5_ASAP7_75t_L g3284 ( 
.A1(n_2996),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_3284)
);

NOR2xp33_ASAP7_75t_SL g3285 ( 
.A(n_2736),
.B(n_3187),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_3104),
.B(n_537),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_2724),
.B(n_289),
.Y(n_3287)
);

INVx3_ASAP7_75t_L g3288 ( 
.A(n_2613),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_3143),
.B(n_537),
.Y(n_3289)
);

O2A1O1Ixp33_ASAP7_75t_L g3290 ( 
.A1(n_2649),
.A2(n_293),
.B(n_290),
.C(n_292),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_L g3291 ( 
.A1(n_3213),
.A2(n_293),
.B1(n_290),
.B2(n_292),
.Y(n_3291)
);

INVx4_ASAP7_75t_L g3292 ( 
.A(n_3213),
.Y(n_3292)
);

NOR2xp33_ASAP7_75t_L g3293 ( 
.A(n_2785),
.B(n_293),
.Y(n_3293)
);

A2O1A1Ixp33_ASAP7_75t_L g3294 ( 
.A1(n_2983),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3068),
.B(n_294),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_2659),
.A2(n_294),
.B(n_295),
.Y(n_3296)
);

AO21x2_ASAP7_75t_L g3297 ( 
.A1(n_2607),
.A2(n_295),
.B(n_296),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3071),
.B(n_296),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_2968),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3072),
.B(n_297),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3097),
.Y(n_3301)
);

INVx3_ASAP7_75t_L g3302 ( 
.A(n_2613),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3099),
.B(n_297),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_3217),
.B(n_538),
.Y(n_3304)
);

INVx2_ASAP7_75t_SL g3305 ( 
.A(n_2698),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2995),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3120),
.B(n_297),
.Y(n_3307)
);

AOI21x1_ASAP7_75t_L g3308 ( 
.A1(n_3015),
.A2(n_298),
.B(n_299),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_3002),
.B(n_3067),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3122),
.B(n_298),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3146),
.Y(n_3311)
);

A2O1A1Ixp33_ASAP7_75t_L g3312 ( 
.A1(n_3017),
.A2(n_300),
.B(n_298),
.C(n_299),
.Y(n_3312)
);

AND2x4_ASAP7_75t_L g3313 ( 
.A(n_2899),
.B(n_300),
.Y(n_3313)
);

INVxp67_ASAP7_75t_SL g3314 ( 
.A(n_3087),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_2942),
.B(n_538),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3173),
.B(n_3177),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3202),
.B(n_300),
.Y(n_3317)
);

OAI21xp33_ASAP7_75t_L g3318 ( 
.A1(n_2862),
.A2(n_301),
.B(n_302),
.Y(n_3318)
);

INVx3_ASAP7_75t_L g3319 ( 
.A(n_2694),
.Y(n_3319)
);

A2O1A1Ixp33_ASAP7_75t_L g3320 ( 
.A1(n_3029),
.A2(n_304),
.B(n_301),
.C(n_303),
.Y(n_3320)
);

O2A1O1Ixp33_ASAP7_75t_L g3321 ( 
.A1(n_2770),
.A2(n_304),
.B(n_301),
.C(n_303),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3009),
.Y(n_3322)
);

NOR3xp33_ASAP7_75t_L g3323 ( 
.A(n_2736),
.B(n_304),
.C(n_305),
.Y(n_3323)
);

NOR2xp67_ASAP7_75t_SL g3324 ( 
.A(n_2851),
.B(n_305),
.Y(n_3324)
);

BUFx6f_ASAP7_75t_L g3325 ( 
.A(n_2605),
.Y(n_3325)
);

OAI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_2617),
.A2(n_305),
.B(n_306),
.Y(n_3326)
);

O2A1O1Ixp33_ASAP7_75t_L g3327 ( 
.A1(n_2784),
.A2(n_308),
.B(n_306),
.C(n_307),
.Y(n_3327)
);

NOR2x1_ASAP7_75t_R g3328 ( 
.A(n_3006),
.B(n_307),
.Y(n_3328)
);

OAI22x1_ASAP7_75t_L g3329 ( 
.A1(n_2775),
.A2(n_3101),
.B1(n_2807),
.B2(n_2969),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_L g3330 ( 
.A(n_3124),
.B(n_307),
.Y(n_3330)
);

BUFx12f_ASAP7_75t_L g3331 ( 
.A(n_2722),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_SL g3332 ( 
.A(n_2721),
.B(n_539),
.Y(n_3332)
);

OAI22x1_ASAP7_75t_L g3333 ( 
.A1(n_2965),
.A2(n_310),
.B1(n_308),
.B2(n_309),
.Y(n_3333)
);

NOR3xp33_ASAP7_75t_SL g3334 ( 
.A(n_3021),
.B(n_308),
.C(n_309),
.Y(n_3334)
);

OA21x2_ASAP7_75t_L g3335 ( 
.A1(n_3019),
.A2(n_309),
.B(n_311),
.Y(n_3335)
);

OAI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_2643),
.A2(n_3012),
.B1(n_2630),
.B2(n_2717),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3016),
.Y(n_3337)
);

HB1xp67_ASAP7_75t_L g3338 ( 
.A(n_3181),
.Y(n_3338)
);

A2O1A1Ixp33_ASAP7_75t_L g3339 ( 
.A1(n_3081),
.A2(n_313),
.B(n_311),
.C(n_312),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3204),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_2661),
.A2(n_311),
.B(n_312),
.Y(n_3341)
);

BUFx3_ASAP7_75t_L g3342 ( 
.A(n_2967),
.Y(n_3342)
);

CKINVDCx5p33_ASAP7_75t_R g3343 ( 
.A(n_3066),
.Y(n_3343)
);

A2O1A1Ixp33_ASAP7_75t_L g3344 ( 
.A1(n_3189),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_3344)
);

INVx1_ASAP7_75t_SL g3345 ( 
.A(n_2779),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_SL g3346 ( 
.A(n_2619),
.B(n_539),
.Y(n_3346)
);

AOI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_2838),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_2701),
.A2(n_314),
.B(n_315),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3219),
.B(n_315),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2683),
.Y(n_3350)
);

AOI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_2905),
.A2(n_316),
.B(n_317),
.Y(n_3351)
);

OAI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_2643),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_2664),
.A2(n_316),
.B(n_318),
.Y(n_3353)
);

AOI21xp5_ASAP7_75t_L g3354 ( 
.A1(n_2604),
.A2(n_318),
.B(n_319),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2755),
.B(n_319),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2684),
.Y(n_3356)
);

INVx2_ASAP7_75t_L g3357 ( 
.A(n_3026),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_2699),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_2762),
.B(n_2621),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_2647),
.B(n_319),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2611),
.B(n_320),
.Y(n_3361)
);

AOI21xp33_ASAP7_75t_L g3362 ( 
.A1(n_2979),
.A2(n_320),
.B(n_321),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_3012),
.B(n_540),
.Y(n_3363)
);

OAI22xp5_ASAP7_75t_L g3364 ( 
.A1(n_2643),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3034),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_3036),
.Y(n_3366)
);

OAI21xp33_ASAP7_75t_SL g3367 ( 
.A1(n_2848),
.A2(n_322),
.B(n_323),
.Y(n_3367)
);

HB1xp67_ASAP7_75t_L g3368 ( 
.A(n_2674),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_2741),
.B(n_323),
.Y(n_3369)
);

BUFx2_ASAP7_75t_L g3370 ( 
.A(n_2687),
.Y(n_3370)
);

NOR2xp67_ASAP7_75t_L g3371 ( 
.A(n_2972),
.B(n_324),
.Y(n_3371)
);

OR2x6_ASAP7_75t_L g3372 ( 
.A(n_3003),
.B(n_324),
.Y(n_3372)
);

AND2x4_ASAP7_75t_L g3373 ( 
.A(n_2902),
.B(n_324),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_2837),
.A2(n_325),
.B(n_326),
.Y(n_3374)
);

HB1xp67_ASAP7_75t_L g3375 ( 
.A(n_2702),
.Y(n_3375)
);

A2O1A1Ixp33_ASAP7_75t_L g3376 ( 
.A1(n_3198),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_2712),
.B(n_2694),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2730),
.B(n_327),
.Y(n_3378)
);

INVx1_ASAP7_75t_SL g3379 ( 
.A(n_2759),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_L g3380 ( 
.A(n_2764),
.B(n_328),
.Y(n_3380)
);

BUFx6f_ASAP7_75t_L g3381 ( 
.A(n_2605),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2637),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_2733),
.B(n_328),
.Y(n_3383)
);

NOR3xp33_ASAP7_75t_L g3384 ( 
.A(n_3187),
.B(n_329),
.C(n_330),
.Y(n_3384)
);

O2A1O1Ixp33_ASAP7_75t_L g3385 ( 
.A1(n_2792),
.A2(n_331),
.B(n_329),
.C(n_330),
.Y(n_3385)
);

HB1xp67_ASAP7_75t_L g3386 ( 
.A(n_3066),
.Y(n_3386)
);

CKINVDCx5p33_ASAP7_75t_R g3387 ( 
.A(n_2788),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_2657),
.A2(n_332),
.B(n_333),
.Y(n_3388)
);

NOR2x1_ASAP7_75t_R g3389 ( 
.A(n_2788),
.B(n_332),
.Y(n_3389)
);

O2A1O1Ixp5_ASAP7_75t_L g3390 ( 
.A1(n_3047),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_2796),
.A2(n_334),
.B(n_335),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_2655),
.A2(n_334),
.B(n_335),
.Y(n_3392)
);

A2O1A1Ixp33_ASAP7_75t_L g3393 ( 
.A1(n_2673),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_3393)
);

OR2x6_ASAP7_75t_L g3394 ( 
.A(n_2951),
.B(n_336),
.Y(n_3394)
);

NOR3xp33_ASAP7_75t_SL g3395 ( 
.A(n_2753),
.B(n_337),
.C(n_338),
.Y(n_3395)
);

NOR2xp33_ASAP7_75t_L g3396 ( 
.A(n_2786),
.B(n_337),
.Y(n_3396)
);

OAI21x1_ASAP7_75t_L g3397 ( 
.A1(n_2623),
.A2(n_338),
.B(n_339),
.Y(n_3397)
);

O2A1O1Ixp33_ASAP7_75t_SL g3398 ( 
.A1(n_2814),
.A2(n_341),
.B(n_339),
.C(n_340),
.Y(n_3398)
);

AOI21x1_ASAP7_75t_L g3399 ( 
.A1(n_3125),
.A2(n_340),
.B(n_342),
.Y(n_3399)
);

INVxp67_ASAP7_75t_L g3400 ( 
.A(n_2800),
.Y(n_3400)
);

AOI221xp5_ASAP7_75t_L g3401 ( 
.A1(n_2587),
.A2(n_343),
.B1(n_340),
.B2(n_342),
.C(n_344),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_2656),
.A2(n_343),
.B(n_344),
.Y(n_3402)
);

O2A1O1Ixp33_ASAP7_75t_L g3403 ( 
.A1(n_2802),
.A2(n_2690),
.B(n_2774),
.C(n_2703),
.Y(n_3403)
);

NAND2x1p5_ASAP7_75t_L g3404 ( 
.A(n_2951),
.B(n_343),
.Y(n_3404)
);

A2O1A1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_2704),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_2880),
.B(n_345),
.Y(n_3406)
);

HB1xp67_ASAP7_75t_L g3407 ( 
.A(n_2638),
.Y(n_3407)
);

A2O1A1Ixp33_ASAP7_75t_L g3408 ( 
.A1(n_2677),
.A2(n_347),
.B(n_345),
.C(n_346),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_L g3409 ( 
.A1(n_2953),
.A2(n_2982),
.B1(n_3056),
.B2(n_3005),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_2885),
.B(n_2729),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_2654),
.A2(n_346),
.B(n_347),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2806),
.Y(n_3412)
);

NOR3xp33_ASAP7_75t_SL g3413 ( 
.A(n_2990),
.B(n_347),
.C(n_348),
.Y(n_3413)
);

INVxp67_ASAP7_75t_L g3414 ( 
.A(n_2999),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3089),
.Y(n_3415)
);

O2A1O1Ixp33_ASAP7_75t_L g3416 ( 
.A1(n_2680),
.A2(n_350),
.B(n_348),
.C(n_349),
.Y(n_3416)
);

O2A1O1Ixp5_ASAP7_75t_L g3417 ( 
.A1(n_3137),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2813),
.Y(n_3418)
);

NAND3xp33_ASAP7_75t_L g3419 ( 
.A(n_2791),
.B(n_349),
.C(n_350),
.Y(n_3419)
);

NOR2xp33_ASAP7_75t_L g3420 ( 
.A(n_2744),
.B(n_351),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_L g3421 ( 
.A(n_2850),
.B(n_351),
.Y(n_3421)
);

NOR2xp33_ASAP7_75t_SL g3422 ( 
.A(n_2687),
.B(n_352),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_2739),
.B(n_352),
.Y(n_3423)
);

A2O1A1Ixp33_ASAP7_75t_SL g3424 ( 
.A1(n_3141),
.A2(n_355),
.B(n_353),
.C(n_354),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2749),
.B(n_354),
.Y(n_3425)
);

BUFx6f_ASAP7_75t_L g3426 ( 
.A(n_2605),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_2828),
.B(n_2834),
.Y(n_3427)
);

NOR2x1_ASAP7_75t_L g3428 ( 
.A(n_2845),
.B(n_355),
.Y(n_3428)
);

NOR2xp33_ASAP7_75t_L g3429 ( 
.A(n_2904),
.B(n_355),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_2985),
.A2(n_3209),
.B(n_3025),
.Y(n_3430)
);

OAI22xp5_ASAP7_75t_L g3431 ( 
.A1(n_2667),
.A2(n_2668),
.B1(n_2893),
.B2(n_2653),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3113),
.Y(n_3432)
);

O2A1O1Ixp33_ASAP7_75t_L g3433 ( 
.A1(n_2695),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_3433)
);

CKINVDCx5p33_ASAP7_75t_R g3434 ( 
.A(n_2877),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3154),
.B(n_356),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3191),
.B(n_357),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_2852),
.A2(n_360),
.B1(n_357),
.B2(n_359),
.Y(n_3437)
);

INVx1_ASAP7_75t_SL g3438 ( 
.A(n_2865),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_L g3439 ( 
.A(n_2911),
.B(n_359),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_2828),
.B(n_541),
.Y(n_3440)
);

BUFx3_ASAP7_75t_L g3441 ( 
.A(n_2847),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_2828),
.B(n_542),
.Y(n_3442)
);

CKINVDCx5p33_ASAP7_75t_R g3443 ( 
.A(n_2860),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_2834),
.B(n_542),
.Y(n_3444)
);

AOI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_2974),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_3445)
);

OAI22xp5_ASAP7_75t_L g3446 ( 
.A1(n_2758),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_2808),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_2795),
.B(n_361),
.Y(n_3448)
);

HB1xp67_ASAP7_75t_L g3449 ( 
.A(n_2940),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_2737),
.B(n_362),
.Y(n_3450)
);

AOI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_2984),
.A2(n_366),
.B1(n_363),
.B2(n_365),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_2761),
.B(n_363),
.Y(n_3452)
);

NAND2xp33_ASAP7_75t_L g3453 ( 
.A(n_2687),
.B(n_2834),
.Y(n_3453)
);

OAI21x1_ASAP7_75t_L g3454 ( 
.A1(n_3175),
.A2(n_363),
.B(n_365),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_3018),
.A2(n_365),
.B(n_366),
.Y(n_3455)
);

INVx3_ASAP7_75t_L g3456 ( 
.A(n_2808),
.Y(n_3456)
);

OR2x2_ASAP7_75t_L g3457 ( 
.A(n_3157),
.B(n_367),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_2612),
.B(n_368),
.Y(n_3458)
);

O2A1O1Ixp33_ASAP7_75t_L g3459 ( 
.A1(n_2854),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_3459)
);

BUFx8_ASAP7_75t_L g3460 ( 
.A(n_2687),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3028),
.A2(n_369),
.B(n_370),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2612),
.B(n_371),
.Y(n_3462)
);

BUFx6f_ASAP7_75t_L g3463 ( 
.A(n_2662),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_SL g3464 ( 
.A(n_2840),
.B(n_543),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_2840),
.B(n_544),
.Y(n_3465)
);

HB1xp67_ASAP7_75t_L g3466 ( 
.A(n_2940),
.Y(n_3466)
);

OR2x2_ASAP7_75t_L g3467 ( 
.A(n_3206),
.B(n_371),
.Y(n_3467)
);

AOI21x1_ASAP7_75t_L g3468 ( 
.A1(n_3180),
.A2(n_372),
.B(n_373),
.Y(n_3468)
);

A2O1A1Ixp33_ASAP7_75t_SL g3469 ( 
.A1(n_3182),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_3469)
);

INVx2_ASAP7_75t_SL g3470 ( 
.A(n_2887),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_2634),
.B(n_2608),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3030),
.A2(n_372),
.B(n_373),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_2634),
.B(n_374),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_2685),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_2646),
.B(n_375),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3134),
.Y(n_3476)
);

BUFx2_ASAP7_75t_L g3477 ( 
.A(n_2697),
.Y(n_3477)
);

A2O1A1Ixp33_ASAP7_75t_L g3478 ( 
.A1(n_2930),
.A2(n_377),
.B(n_375),
.C(n_376),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_2804),
.B(n_375),
.Y(n_3479)
);

NOR2xp33_ASAP7_75t_L g3480 ( 
.A(n_2689),
.B(n_376),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3145),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2610),
.B(n_376),
.Y(n_3482)
);

BUFx3_ASAP7_75t_L g3483 ( 
.A(n_2890),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_2688),
.Y(n_3484)
);

BUFx3_ASAP7_75t_L g3485 ( 
.A(n_2945),
.Y(n_3485)
);

AOI21x1_ASAP7_75t_L g3486 ( 
.A1(n_3196),
.A2(n_378),
.B(n_379),
.Y(n_3486)
);

OR2x2_ASAP7_75t_L g3487 ( 
.A(n_2757),
.B(n_2763),
.Y(n_3487)
);

A2O1A1Ixp33_ASAP7_75t_L g3488 ( 
.A1(n_2933),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_3488)
);

CKINVDCx5p33_ASAP7_75t_R g3489 ( 
.A(n_2594),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_2988),
.B(n_378),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_2748),
.Y(n_3491)
);

BUFx3_ASAP7_75t_L g3492 ( 
.A(n_2949),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_2614),
.B(n_380),
.Y(n_3493)
);

INVx1_ASAP7_75t_SL g3494 ( 
.A(n_2797),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3102),
.Y(n_3495)
);

INVx3_ASAP7_75t_L g3496 ( 
.A(n_2589),
.Y(n_3496)
);

NOR3xp33_ASAP7_75t_SL g3497 ( 
.A(n_2994),
.B(n_380),
.C(n_381),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3037),
.A2(n_381),
.B(n_382),
.Y(n_3498)
);

INVx1_ASAP7_75t_SL g3499 ( 
.A(n_2941),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_2615),
.B(n_381),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_2835),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_2676),
.Y(n_3502)
);

AND2x4_ASAP7_75t_L g3503 ( 
.A(n_2820),
.B(n_2943),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3150),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_2840),
.B(n_545),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3038),
.A2(n_382),
.B(n_383),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_2707),
.Y(n_3507)
);

NOR3xp33_ASAP7_75t_L g3508 ( 
.A(n_3119),
.B(n_2921),
.C(n_2912),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_2918),
.B(n_545),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2946),
.Y(n_3510)
);

A2O1A1Ixp33_ASAP7_75t_L g3511 ( 
.A1(n_2691),
.A2(n_385),
.B(n_382),
.C(n_383),
.Y(n_3511)
);

NOR3xp33_ASAP7_75t_L g3512 ( 
.A(n_2973),
.B(n_383),
.C(n_386),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_2639),
.B(n_386),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_R g3514 ( 
.A(n_2589),
.B(n_387),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3152),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_2675),
.B(n_387),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3043),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_3517)
);

O2A1O1Ixp33_ASAP7_75t_L g3518 ( 
.A1(n_2881),
.A2(n_391),
.B(n_388),
.C(n_390),
.Y(n_3518)
);

A2O1A1Ixp33_ASAP7_75t_L g3519 ( 
.A1(n_2670),
.A2(n_391),
.B(n_388),
.C(n_390),
.Y(n_3519)
);

HB1xp67_ASAP7_75t_L g3520 ( 
.A(n_2941),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_2948),
.Y(n_3521)
);

CKINVDCx20_ASAP7_75t_R g3522 ( 
.A(n_2980),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3197),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_2640),
.B(n_390),
.Y(n_3524)
);

NAND3xp33_ASAP7_75t_SL g3525 ( 
.A(n_2706),
.B(n_391),
.C(n_392),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_2821),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3045),
.A2(n_392),
.B(n_393),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_2628),
.B(n_393),
.Y(n_3528)
);

INVxp67_ASAP7_75t_L g3529 ( 
.A(n_2991),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3210),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_2632),
.B(n_394),
.Y(n_3531)
);

INVx3_ASAP7_75t_L g3532 ( 
.A(n_2592),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3048),
.A2(n_3193),
.B(n_3192),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_2650),
.B(n_394),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_2918),
.Y(n_3535)
);

BUFx3_ASAP7_75t_L g3536 ( 
.A(n_2592),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_2666),
.B(n_546),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_2662),
.Y(n_3538)
);

AOI22xp5_ASAP7_75t_L g3539 ( 
.A1(n_2993),
.A2(n_3054),
.B1(n_3070),
.B2(n_3061),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3211),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_2679),
.B(n_395),
.Y(n_3541)
);

NOR2xp33_ASAP7_75t_L g3542 ( 
.A(n_2819),
.B(n_395),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3077),
.B(n_395),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3096),
.B(n_396),
.Y(n_3544)
);

CKINVDCx5p33_ASAP7_75t_R g3545 ( 
.A(n_3007),
.Y(n_3545)
);

AOI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_3052),
.A2(n_396),
.B(n_397),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3100),
.B(n_396),
.Y(n_3547)
);

NOR2xp33_ASAP7_75t_SL g3548 ( 
.A(n_2745),
.B(n_397),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_L g3549 ( 
.A1(n_3138),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2866),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_2666),
.B(n_547),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_3059),
.A2(n_3065),
.B(n_3060),
.Y(n_3552)
);

INVx1_ASAP7_75t_SL g3553 ( 
.A(n_2939),
.Y(n_3553)
);

A2O1A1Ixp33_ASAP7_75t_L g3554 ( 
.A1(n_2740),
.A2(n_400),
.B(n_398),
.C(n_399),
.Y(n_3554)
);

INVx3_ASAP7_75t_L g3555 ( 
.A(n_3022),
.Y(n_3555)
);

NOR2xp33_ASAP7_75t_L g3556 ( 
.A(n_3149),
.B(n_398),
.Y(n_3556)
);

AOI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_3162),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_3557)
);

OAI21x1_ASAP7_75t_L g3558 ( 
.A1(n_3200),
.A2(n_400),
.B(n_401),
.Y(n_3558)
);

BUFx8_ASAP7_75t_L g3559 ( 
.A(n_2950),
.Y(n_3559)
);

INVxp67_ASAP7_75t_L g3560 ( 
.A(n_3218),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3078),
.A2(n_401),
.B(n_402),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3079),
.A2(n_402),
.B(n_403),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_2975),
.Y(n_3563)
);

A2O1A1Ixp33_ASAP7_75t_SL g3564 ( 
.A1(n_3205),
.A2(n_406),
.B(n_404),
.C(n_405),
.Y(n_3564)
);

AOI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_2932),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_3565)
);

NOR3xp33_ASAP7_75t_SL g3566 ( 
.A(n_3004),
.B(n_404),
.C(n_405),
.Y(n_3566)
);

O2A1O1Ixp33_ASAP7_75t_L g3567 ( 
.A1(n_2803),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_3080),
.A2(n_407),
.B(n_408),
.Y(n_3568)
);

INVx2_ASAP7_75t_SL g3569 ( 
.A(n_3022),
.Y(n_3569)
);

O2A1O1Ixp33_ASAP7_75t_L g3570 ( 
.A1(n_3041),
.A2(n_411),
.B(n_409),
.C(n_410),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_3033),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_2582),
.B(n_409),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_3082),
.A2(n_410),
.B(n_411),
.Y(n_3573)
);

A2O1A1Ixp33_ASAP7_75t_L g3574 ( 
.A1(n_2892),
.A2(n_413),
.B(n_410),
.C(n_412),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3151),
.Y(n_3575)
);

AOI21x1_ASAP7_75t_L g3576 ( 
.A1(n_2631),
.A2(n_412),
.B(n_413),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3083),
.A2(n_413),
.B(n_414),
.Y(n_3577)
);

BUFx6f_ASAP7_75t_L g3578 ( 
.A(n_2662),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_2815),
.B(n_547),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_2920),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_2962),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3159),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_3084),
.A2(n_414),
.B(n_415),
.Y(n_3583)
);

BUFx6f_ASAP7_75t_L g3584 ( 
.A(n_2962),
.Y(n_3584)
);

NOR2xp33_ASAP7_75t_L g3585 ( 
.A(n_2598),
.B(n_414),
.Y(n_3585)
);

O2A1O1Ixp5_ASAP7_75t_L g3586 ( 
.A1(n_2622),
.A2(n_418),
.B(n_415),
.C(n_416),
.Y(n_3586)
);

BUFx6f_ASAP7_75t_L g3587 ( 
.A(n_2962),
.Y(n_3587)
);

CKINVDCx16_ASAP7_75t_R g3588 ( 
.A(n_3166),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3091),
.A2(n_415),
.B(n_416),
.Y(n_3589)
);

OAI21xp33_ASAP7_75t_SL g3590 ( 
.A1(n_2752),
.A2(n_416),
.B(n_418),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_SL g3591 ( 
.A(n_2815),
.B(n_548),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_SL g3592 ( 
.A(n_3058),
.B(n_3139),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3161),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3174),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3053),
.B(n_418),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3207),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3094),
.A2(n_419),
.B(n_420),
.Y(n_3597)
);

AOI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_2743),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_2833),
.B(n_419),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_2669),
.B(n_420),
.Y(n_3600)
);

AO21x1_ASAP7_75t_L g3601 ( 
.A1(n_2693),
.A2(n_550),
.B(n_549),
.Y(n_3601)
);

HB1xp67_ASAP7_75t_L g3602 ( 
.A(n_2830),
.Y(n_3602)
);

OAI22x1_ASAP7_75t_L g3603 ( 
.A1(n_2934),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3058),
.B(n_551),
.Y(n_3604)
);

O2A1O1Ixp5_ASAP7_75t_L g3605 ( 
.A1(n_2641),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_2799),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_2901),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3103),
.B(n_422),
.Y(n_3608)
);

CKINVDCx6p67_ASAP7_75t_R g3609 ( 
.A(n_2760),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3139),
.B(n_2971),
.Y(n_3610)
);

OAI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3107),
.A2(n_3114),
.B1(n_3116),
.B2(n_3111),
.Y(n_3611)
);

INVxp67_ASAP7_75t_SL g3612 ( 
.A(n_2971),
.Y(n_3612)
);

CKINVDCx5p33_ASAP7_75t_R g3613 ( 
.A(n_2681),
.Y(n_3613)
);

AND2x4_ASAP7_75t_L g3614 ( 
.A(n_2874),
.B(n_423),
.Y(n_3614)
);

AND2x2_ASAP7_75t_L g3615 ( 
.A(n_2981),
.B(n_2718),
.Y(n_3615)
);

O2A1O1Ixp33_ASAP7_75t_L g3616 ( 
.A1(n_3117),
.A2(n_426),
.B(n_424),
.C(n_425),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_2971),
.B(n_551),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_3129),
.A2(n_424),
.B(n_425),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_2624),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3130),
.A2(n_3148),
.B(n_3132),
.Y(n_3620)
);

OAI21xp33_ASAP7_75t_L g3621 ( 
.A1(n_3044),
.A2(n_425),
.B(n_426),
.Y(n_3621)
);

HB1xp67_ASAP7_75t_L g3622 ( 
.A(n_2842),
.Y(n_3622)
);

A2O1A1Ixp33_ASAP7_75t_L g3623 ( 
.A1(n_2781),
.A2(n_429),
.B(n_426),
.C(n_428),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3155),
.B(n_429),
.Y(n_3624)
);

A2O1A1Ixp33_ASAP7_75t_L g3625 ( 
.A1(n_2782),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_3625)
);

HB1xp67_ASAP7_75t_L g3626 ( 
.A(n_2665),
.Y(n_3626)
);

OAI22xp5_ASAP7_75t_L g3627 ( 
.A1(n_3165),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_3627)
);

NAND3xp33_ASAP7_75t_SL g3628 ( 
.A(n_2651),
.B(n_430),
.C(n_431),
.Y(n_3628)
);

AOI22xp33_ASAP7_75t_L g3629 ( 
.A1(n_2846),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_3629)
);

O2A1O1Ixp33_ASAP7_75t_L g3630 ( 
.A1(n_3123),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3167),
.B(n_435),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_SL g3632 ( 
.A(n_3069),
.B(n_435),
.Y(n_3632)
);

OAI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_2644),
.A2(n_436),
.B(n_437),
.Y(n_3633)
);

OR2x6_ASAP7_75t_SL g3634 ( 
.A(n_2914),
.B(n_436),
.Y(n_3634)
);

BUFx3_ASAP7_75t_L g3635 ( 
.A(n_3040),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_L g3636 ( 
.A(n_3142),
.B(n_436),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3170),
.A2(n_437),
.B(n_438),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3176),
.B(n_437),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_L g3639 ( 
.A(n_3169),
.B(n_438),
.Y(n_3639)
);

BUFx6f_ASAP7_75t_L g3640 ( 
.A(n_2977),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3188),
.B(n_438),
.Y(n_3641)
);

AOI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_3190),
.A2(n_439),
.B(n_440),
.Y(n_3642)
);

AOI21xp33_ASAP7_75t_L g3643 ( 
.A1(n_3203),
.A2(n_439),
.B(n_440),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_2863),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_3644)
);

INVxp67_ASAP7_75t_L g3645 ( 
.A(n_2895),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3172),
.B(n_441),
.Y(n_3646)
);

O2A1O1Ixp33_ASAP7_75t_L g3647 ( 
.A1(n_2858),
.A2(n_443),
.B(n_441),
.C(n_442),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_2908),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_2626),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_2960),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_2627),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_2746),
.B(n_442),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_2636),
.Y(n_3653)
);

OR2x6_ASAP7_75t_L g3654 ( 
.A(n_2935),
.B(n_443),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_2961),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_2888),
.B(n_443),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_2977),
.B(n_552),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_2719),
.B(n_444),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_2927),
.Y(n_3659)
);

AOI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_2856),
.A2(n_445),
.B(n_446),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_2597),
.B(n_445),
.Y(n_3661)
);

BUFx6f_ASAP7_75t_L g3662 ( 
.A(n_2977),
.Y(n_3662)
);

BUFx6f_ASAP7_75t_L g3663 ( 
.A(n_3014),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_2936),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_2696),
.B(n_445),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_2771),
.B(n_446),
.Y(n_3666)
);

NOR3xp33_ASAP7_75t_L g3667 ( 
.A(n_3076),
.B(n_446),
.C(n_447),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_SL g3668 ( 
.A(n_3014),
.B(n_553),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_2776),
.B(n_447),
.Y(n_3669)
);

AOI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_2836),
.A2(n_448),
.B(n_449),
.Y(n_3670)
);

HB1xp67_ASAP7_75t_L g3671 ( 
.A(n_2809),
.Y(n_3671)
);

INVx2_ASAP7_75t_L g3672 ( 
.A(n_3001),
.Y(n_3672)
);

CKINVDCx5p33_ASAP7_75t_R g3673 ( 
.A(n_2822),
.Y(n_3673)
);

HB1xp67_ASAP7_75t_L g3674 ( 
.A(n_2925),
.Y(n_3674)
);

A2O1A1Ixp33_ASAP7_75t_L g3675 ( 
.A1(n_2787),
.A2(n_450),
.B(n_448),
.C(n_449),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_2700),
.B(n_449),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_2903),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_SL g3678 ( 
.A(n_3088),
.B(n_3014),
.Y(n_3678)
);

BUFx6f_ASAP7_75t_L g3679 ( 
.A(n_3023),
.Y(n_3679)
);

BUFx2_ASAP7_75t_L g3680 ( 
.A(n_3040),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_2861),
.Y(n_3681)
);

INVx1_ASAP7_75t_SL g3682 ( 
.A(n_3057),
.Y(n_3682)
);

O2A1O1Ixp33_ASAP7_75t_L g3683 ( 
.A1(n_2625),
.A2(n_2929),
.B(n_2593),
.C(n_3049),
.Y(n_3683)
);

INVx2_ASAP7_75t_SL g3684 ( 
.A(n_3057),
.Y(n_3684)
);

O2A1O1Ixp33_ASAP7_75t_L g3685 ( 
.A1(n_3171),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_3685)
);

BUFx2_ASAP7_75t_L g3686 ( 
.A(n_3147),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_SL g3687 ( 
.A(n_3023),
.B(n_553),
.Y(n_3687)
);

NOR2xp33_ASAP7_75t_L g3688 ( 
.A(n_2716),
.B(n_2723),
.Y(n_3688)
);

INVx1_ASAP7_75t_SL g3689 ( 
.A(n_3147),
.Y(n_3689)
);

BUFx3_ASAP7_75t_L g3690 ( 
.A(n_3160),
.Y(n_3690)
);

AO32x1_ASAP7_75t_L g3691 ( 
.A1(n_3055),
.A2(n_3131),
.A3(n_3186),
.B1(n_2710),
.B2(n_2750),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3020),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_2812),
.Y(n_3693)
);

AOI22x1_ASAP7_75t_SL g3694 ( 
.A1(n_3160),
.A2(n_454),
.B1(n_455),
.B2(n_453),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_2728),
.B(n_452),
.Y(n_3695)
);

BUFx6f_ASAP7_75t_L g3696 ( 
.A(n_3023),
.Y(n_3696)
);

BUFx3_ASAP7_75t_L g3697 ( 
.A(n_3199),
.Y(n_3697)
);

NAND2x1p5_ASAP7_75t_L g3698 ( 
.A(n_3199),
.B(n_453),
.Y(n_3698)
);

CKINVDCx5p33_ASAP7_75t_R g3699 ( 
.A(n_2926),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_L g3700 ( 
.A(n_2751),
.B(n_454),
.Y(n_3700)
);

OAI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_2924),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_3701)
);

O2A1O1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_2829),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_3702)
);

O2A1O1Ixp33_ASAP7_75t_L g3703 ( 
.A1(n_2734),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3064),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3136),
.Y(n_3705)
);

OAI21xp33_ASAP7_75t_L g3706 ( 
.A1(n_2875),
.A2(n_458),
.B(n_459),
.Y(n_3706)
);

NAND3xp33_ASAP7_75t_SL g3707 ( 
.A(n_2780),
.B(n_458),
.C(n_459),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_R g3708 ( 
.A(n_2783),
.B(n_460),
.Y(n_3708)
);

BUFx2_ASAP7_75t_L g3709 ( 
.A(n_2874),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_L g3710 ( 
.A(n_2909),
.B(n_460),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_2586),
.B(n_460),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_2922),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_2944),
.B(n_461),
.Y(n_3713)
);

BUFx8_ASAP7_75t_L g3714 ( 
.A(n_2910),
.Y(n_3714)
);

BUFx2_ASAP7_75t_L g3715 ( 
.A(n_2747),
.Y(n_3715)
);

INVx2_ASAP7_75t_SL g3716 ( 
.A(n_2898),
.Y(n_3716)
);

BUFx3_ASAP7_75t_L g3717 ( 
.A(n_3051),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_2585),
.A2(n_461),
.B(n_462),
.Y(n_3718)
);

NAND3xp33_ASAP7_75t_L g3719 ( 
.A(n_2978),
.B(n_462),
.C(n_463),
.Y(n_3719)
);

INVx3_ASAP7_75t_L g3720 ( 
.A(n_3051),
.Y(n_3720)
);

OAI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_2583),
.A2(n_462),
.B(n_463),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_2588),
.B(n_464),
.Y(n_3722)
);

OAI21xp33_ASAP7_75t_SL g3723 ( 
.A1(n_2754),
.A2(n_464),
.B(n_465),
.Y(n_3723)
);

OA22x2_ASAP7_75t_L g3724 ( 
.A1(n_2756),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.Y(n_3724)
);

NOR2xp67_ASAP7_75t_L g3725 ( 
.A(n_2738),
.B(n_2672),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_2958),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_3051),
.B(n_3095),
.Y(n_3727)
);

INVx6_ASAP7_75t_L g3728 ( 
.A(n_2766),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3075),
.Y(n_3729)
);

CKINVDCx5p33_ASAP7_75t_R g3730 ( 
.A(n_2769),
.Y(n_3730)
);

INVx2_ASAP7_75t_SL g3731 ( 
.A(n_2898),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_2618),
.B(n_465),
.Y(n_3732)
);

OAI21x1_ASAP7_75t_L g3733 ( 
.A1(n_2765),
.A2(n_466),
.B(n_467),
.Y(n_3733)
);

OAI22xp5_ASAP7_75t_L g3734 ( 
.A1(n_2900),
.A2(n_2817),
.B1(n_2777),
.B2(n_2801),
.Y(n_3734)
);

BUFx6f_ASAP7_75t_L g3735 ( 
.A(n_3095),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_2599),
.B(n_466),
.Y(n_3736)
);

BUFx6f_ASAP7_75t_L g3737 ( 
.A(n_3095),
.Y(n_3737)
);

NOR2xp33_ASAP7_75t_L g3738 ( 
.A(n_2857),
.B(n_467),
.Y(n_3738)
);

AND2x4_ASAP7_75t_L g3739 ( 
.A(n_2867),
.B(n_467),
.Y(n_3739)
);

NOR2xp33_ASAP7_75t_L g3740 ( 
.A(n_2869),
.B(n_468),
.Y(n_3740)
);

NOR3xp33_ASAP7_75t_SL g3741 ( 
.A(n_2773),
.B(n_468),
.C(n_469),
.Y(n_3741)
);

INVx1_ASAP7_75t_SL g3742 ( 
.A(n_2827),
.Y(n_3742)
);

NOR2xp33_ASAP7_75t_L g3743 ( 
.A(n_2894),
.B(n_468),
.Y(n_3743)
);

NOR2xp33_ASAP7_75t_L g3744 ( 
.A(n_2635),
.B(n_469),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_2966),
.Y(n_3745)
);

A2O1A1Ixp33_ASAP7_75t_L g3746 ( 
.A1(n_2790),
.A2(n_472),
.B(n_470),
.C(n_471),
.Y(n_3746)
);

AOI21x1_ASAP7_75t_L g3747 ( 
.A1(n_2686),
.A2(n_470),
.B(n_471),
.Y(n_3747)
);

A2O1A1Ixp33_ASAP7_75t_L g3748 ( 
.A1(n_2793),
.A2(n_473),
.B(n_471),
.C(n_472),
.Y(n_3748)
);

OAI21x1_ASAP7_75t_L g3749 ( 
.A1(n_2765),
.A2(n_472),
.B(n_473),
.Y(n_3749)
);

O2A1O1Ixp33_ASAP7_75t_L g3750 ( 
.A1(n_3042),
.A2(n_3183),
.B(n_3201),
.C(n_3085),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3075),
.Y(n_3751)
);

CKINVDCx5p33_ASAP7_75t_R g3752 ( 
.A(n_2938),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_SL g3753 ( 
.A(n_3179),
.B(n_554),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_2591),
.B(n_473),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3430),
.A2(n_3179),
.B(n_2768),
.Y(n_3755)
);

OAI22xp5_ASAP7_75t_L g3756 ( 
.A1(n_3270),
.A2(n_2708),
.B1(n_2705),
.B2(n_2726),
.Y(n_3756)
);

BUFx2_ASAP7_75t_L g3757 ( 
.A(n_3714),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3495),
.B(n_2794),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3533),
.A2(n_3179),
.B(n_2768),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_3552),
.A2(n_3620),
.B(n_3336),
.Y(n_3760)
);

OAI21x1_ASAP7_75t_L g3761 ( 
.A1(n_3650),
.A2(n_3121),
.B(n_2883),
.Y(n_3761)
);

AND2x4_ASAP7_75t_L g3762 ( 
.A(n_3237),
.B(n_2876),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3655),
.A2(n_2868),
.B(n_2727),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3243),
.Y(n_3764)
);

OAI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3403),
.A2(n_2891),
.B(n_2916),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_3489),
.B(n_2889),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3359),
.B(n_2798),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_SL g3768 ( 
.A1(n_3292),
.A2(n_2713),
.B(n_2831),
.Y(n_3768)
);

O2A1O1Ixp33_ASAP7_75t_L g3769 ( 
.A1(n_3611),
.A2(n_3216),
.B(n_3212),
.C(n_2720),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3422),
.A2(n_3734),
.B(n_3431),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3453),
.A2(n_2768),
.B(n_2766),
.Y(n_3771)
);

O2A1O1Ixp33_ASAP7_75t_SL g3772 ( 
.A1(n_3408),
.A2(n_2603),
.B(n_2907),
.C(n_2937),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3259),
.Y(n_3773)
);

OAI21x1_ASAP7_75t_L g3774 ( 
.A1(n_3672),
.A2(n_2732),
.B(n_2725),
.Y(n_3774)
);

AOI21x1_ASAP7_75t_L g3775 ( 
.A1(n_3692),
.A2(n_2660),
.B(n_2642),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3704),
.A2(n_3128),
.B(n_3010),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3619),
.B(n_2811),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3649),
.B(n_2816),
.Y(n_3778)
);

O2A1O1Ixp5_ASAP7_75t_L g3779 ( 
.A1(n_3592),
.A2(n_2789),
.B(n_2678),
.C(n_2956),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3705),
.A2(n_2711),
.B(n_2709),
.Y(n_3780)
);

AOI221x1_ASAP7_75t_L g3781 ( 
.A1(n_3525),
.A2(n_2714),
.B1(n_2917),
.B2(n_2841),
.C(n_2959),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3727),
.A2(n_2772),
.B(n_2766),
.Y(n_3782)
);

NOR2xp33_ASAP7_75t_L g3783 ( 
.A(n_3292),
.B(n_2778),
.Y(n_3783)
);

INVx4_ASAP7_75t_L g3784 ( 
.A(n_3220),
.Y(n_3784)
);

A2O1A1Ixp33_ASAP7_75t_L g3785 ( 
.A1(n_3590),
.A2(n_2884),
.B(n_2864),
.C(n_2805),
.Y(n_3785)
);

BUFx2_ASAP7_75t_L g3786 ( 
.A(n_3714),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_SL g3787 ( 
.A(n_3370),
.B(n_2772),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3234),
.Y(n_3788)
);

BUFx2_ASAP7_75t_L g3789 ( 
.A(n_3460),
.Y(n_3789)
);

INVx3_ASAP7_75t_SL g3790 ( 
.A(n_3229),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3263),
.Y(n_3791)
);

INVxp67_ASAP7_75t_L g3792 ( 
.A(n_3309),
.Y(n_3792)
);

AO21x2_ASAP7_75t_L g3793 ( 
.A1(n_3580),
.A2(n_2652),
.B(n_2970),
.Y(n_3793)
);

AOI21x1_ASAP7_75t_L g3794 ( 
.A1(n_3729),
.A2(n_3751),
.B(n_3610),
.Y(n_3794)
);

AO32x2_ASAP7_75t_L g3795 ( 
.A1(n_3252),
.A2(n_2652),
.A3(n_2913),
.B1(n_2879),
.B2(n_2873),
.Y(n_3795)
);

OA21x2_ASAP7_75t_L g3796 ( 
.A1(n_3454),
.A2(n_2871),
.B(n_2870),
.Y(n_3796)
);

OAI21xp5_ASAP7_75t_L g3797 ( 
.A1(n_3257),
.A2(n_2663),
.B(n_2742),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3651),
.B(n_2824),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3653),
.B(n_3221),
.Y(n_3799)
);

BUFx3_ASAP7_75t_L g3800 ( 
.A(n_3331),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3479),
.B(n_2825),
.Y(n_3801)
);

OAI221xp5_ASAP7_75t_L g3802 ( 
.A1(n_3539),
.A2(n_2826),
.B1(n_2897),
.B2(n_2832),
.C(n_2853),
.Y(n_3802)
);

AO32x2_ASAP7_75t_L g3803 ( 
.A1(n_3352),
.A2(n_2844),
.A3(n_2986),
.B1(n_2987),
.B2(n_2976),
.Y(n_3803)
);

NOR2xp33_ASAP7_75t_SL g3804 ( 
.A(n_3285),
.B(n_2772),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3691),
.A2(n_2818),
.B(n_2810),
.Y(n_3805)
);

INVx3_ASAP7_75t_SL g3806 ( 
.A(n_3241),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3267),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3275),
.Y(n_3808)
);

INVx1_ASAP7_75t_SL g3809 ( 
.A(n_3379),
.Y(n_3809)
);

A2O1A1Ixp33_ASAP7_75t_L g3810 ( 
.A1(n_3723),
.A2(n_2992),
.B(n_2998),
.C(n_2997),
.Y(n_3810)
);

OAI21x1_ASAP7_75t_L g3811 ( 
.A1(n_3397),
.A2(n_3011),
.B(n_3000),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3634),
.A2(n_3024),
.B1(n_3032),
.B2(n_3031),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3278),
.Y(n_3813)
);

OAI21x1_ASAP7_75t_L g3814 ( 
.A1(n_3576),
.A2(n_3050),
.B(n_3035),
.Y(n_3814)
);

BUFx3_ASAP7_75t_L g3815 ( 
.A(n_3254),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3691),
.A2(n_2818),
.B(n_2810),
.Y(n_3816)
);

NAND3xp33_ASAP7_75t_L g3817 ( 
.A(n_3323),
.B(n_3384),
.C(n_3508),
.Y(n_3817)
);

AOI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_3522),
.A2(n_2919),
.B1(n_2906),
.B2(n_2915),
.Y(n_3818)
);

INVxp67_ASAP7_75t_SL g3819 ( 
.A(n_3460),
.Y(n_3819)
);

O2A1O1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_3400),
.A2(n_2947),
.B(n_3073),
.C(n_3063),
.Y(n_3820)
);

HB1xp67_ASAP7_75t_L g3821 ( 
.A(n_3338),
.Y(n_3821)
);

AOI211x1_ASAP7_75t_L g3822 ( 
.A1(n_3277),
.A2(n_3324),
.B(n_3363),
.C(n_3236),
.Y(n_3822)
);

OAI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3284),
.A2(n_3092),
.B(n_3086),
.Y(n_3823)
);

AO31x2_ASAP7_75t_L g3824 ( 
.A1(n_3601),
.A2(n_3098),
.A3(n_3106),
.B(n_3105),
.Y(n_3824)
);

OAI21x1_ASAP7_75t_L g3825 ( 
.A1(n_3720),
.A2(n_3109),
.B(n_3108),
.Y(n_3825)
);

OAI21x1_ASAP7_75t_L g3826 ( 
.A1(n_3720),
.A2(n_3115),
.B(n_3110),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3545),
.B(n_3571),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3691),
.A2(n_2818),
.B(n_2810),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3281),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3301),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3293),
.B(n_3140),
.Y(n_3831)
);

AOI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3308),
.A2(n_3126),
.B(n_3118),
.Y(n_3832)
);

NOR3xp33_ASAP7_75t_L g3833 ( 
.A(n_3389),
.B(n_3133),
.C(n_3127),
.Y(n_3833)
);

O2A1O1Ixp33_ASAP7_75t_L g3834 ( 
.A1(n_3645),
.A2(n_3144),
.B(n_3156),
.C(n_3153),
.Y(n_3834)
);

O2A1O1Ixp33_ASAP7_75t_L g3835 ( 
.A1(n_3688),
.A2(n_3158),
.B(n_3164),
.C(n_3163),
.Y(n_3835)
);

NAND3xp33_ASAP7_75t_L g3836 ( 
.A(n_3413),
.B(n_3178),
.C(n_3168),
.Y(n_3836)
);

AOI21xp5_ASAP7_75t_L g3837 ( 
.A1(n_3548),
.A2(n_2602),
.B(n_2931),
.Y(n_3837)
);

BUFx8_ASAP7_75t_L g3838 ( 
.A(n_3305),
.Y(n_3838)
);

O2A1O1Ixp33_ASAP7_75t_SL g3839 ( 
.A1(n_3478),
.A2(n_3184),
.B(n_3208),
.C(n_3185),
.Y(n_3839)
);

NAND3x1_ASAP7_75t_L g3840 ( 
.A(n_3256),
.B(n_3215),
.C(n_3214),
.Y(n_3840)
);

AO31x2_ASAP7_75t_L g3841 ( 
.A1(n_3715),
.A2(n_2878),
.A3(n_2928),
.B(n_2931),
.Y(n_3841)
);

OAI21x1_ASAP7_75t_L g3842 ( 
.A1(n_3558),
.A2(n_476),
.B(n_475),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3238),
.Y(n_3843)
);

A2O1A1Ixp33_ASAP7_75t_L g3844 ( 
.A1(n_3703),
.A2(n_476),
.B(n_474),
.C(n_475),
.Y(n_3844)
);

INVx3_ASAP7_75t_L g3845 ( 
.A(n_3255),
.Y(n_3845)
);

OR2x2_ASAP7_75t_L g3846 ( 
.A(n_3235),
.B(n_3314),
.Y(n_3846)
);

AOI21xp5_ASAP7_75t_L g3847 ( 
.A1(n_3725),
.A2(n_3726),
.B(n_3745),
.Y(n_3847)
);

O2A1O1Ixp33_ASAP7_75t_L g3848 ( 
.A1(n_3511),
.A2(n_477),
.B(n_474),
.C(n_476),
.Y(n_3848)
);

OAI21x1_ASAP7_75t_L g3849 ( 
.A1(n_3399),
.A2(n_479),
.B(n_478),
.Y(n_3849)
);

OAI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3390),
.A2(n_477),
.B(n_478),
.Y(n_3850)
);

A2O1A1Ixp33_ASAP7_75t_L g3851 ( 
.A1(n_3367),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3311),
.B(n_479),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3340),
.B(n_3350),
.Y(n_3853)
);

OR2x2_ASAP7_75t_L g3854 ( 
.A(n_3457),
.B(n_3467),
.Y(n_3854)
);

BUFx6f_ASAP7_75t_L g3855 ( 
.A(n_3245),
.Y(n_3855)
);

OA22x2_ASAP7_75t_L g3856 ( 
.A1(n_3494),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3750),
.A2(n_480),
.B(n_481),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3615),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_3858)
);

OAI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_3417),
.A2(n_483),
.B(n_484),
.Y(n_3859)
);

OAI21xp5_ASAP7_75t_L g3860 ( 
.A1(n_3683),
.A2(n_3409),
.B(n_3719),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_3424),
.A2(n_483),
.B(n_484),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_SL g3862 ( 
.A1(n_3654),
.A2(n_483),
.B(n_484),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3356),
.B(n_485),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3358),
.B(n_485),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3382),
.Y(n_3865)
);

OAI21x1_ASAP7_75t_L g3866 ( 
.A1(n_3468),
.A2(n_487),
.B(n_486),
.Y(n_3866)
);

OAI21x1_ASAP7_75t_L g3867 ( 
.A1(n_3486),
.A2(n_487),
.B(n_486),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3242),
.Y(n_3868)
);

A2O1A1Ixp33_ASAP7_75t_L g3869 ( 
.A1(n_3321),
.A2(n_3327),
.B(n_3433),
.C(n_3567),
.Y(n_3869)
);

A2O1A1Ixp33_ASAP7_75t_L g3870 ( 
.A1(n_3239),
.A2(n_488),
.B(n_485),
.C(n_486),
.Y(n_3870)
);

AND2x2_ASAP7_75t_L g3871 ( 
.A(n_3287),
.B(n_488),
.Y(n_3871)
);

OAI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3271),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_3872)
);

NOR2x1_ASAP7_75t_R g3873 ( 
.A(n_3227),
.B(n_489),
.Y(n_3873)
);

INVx8_ASAP7_75t_L g3874 ( 
.A(n_3394),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3471),
.B(n_490),
.Y(n_3875)
);

AO22x2_ASAP7_75t_L g3876 ( 
.A1(n_3694),
.A2(n_494),
.B1(n_491),
.B2(n_493),
.Y(n_3876)
);

O2A1O1Ixp33_ASAP7_75t_L g3877 ( 
.A1(n_3519),
.A2(n_494),
.B(n_491),
.C(n_493),
.Y(n_3877)
);

O2A1O1Ixp33_ASAP7_75t_SL g3878 ( 
.A1(n_3488),
.A2(n_496),
.B(n_491),
.C(n_495),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3469),
.A2(n_3564),
.B(n_3633),
.Y(n_3879)
);

A2O1A1Ixp33_ASAP7_75t_L g3880 ( 
.A1(n_3248),
.A2(n_497),
.B(n_495),
.C(n_496),
.Y(n_3880)
);

OAI21x1_ASAP7_75t_L g3881 ( 
.A1(n_3427),
.A2(n_497),
.B(n_496),
.Y(n_3881)
);

INVxp67_ASAP7_75t_SL g3882 ( 
.A(n_3407),
.Y(n_3882)
);

OAI21x1_ASAP7_75t_L g3883 ( 
.A1(n_3733),
.A2(n_498),
.B(n_497),
.Y(n_3883)
);

AO21x1_ASAP7_75t_L g3884 ( 
.A1(n_3632),
.A2(n_495),
.B(n_498),
.Y(n_3884)
);

INVxp67_ASAP7_75t_L g3885 ( 
.A(n_3253),
.Y(n_3885)
);

AO31x2_ASAP7_75t_L g3886 ( 
.A1(n_3348),
.A2(n_501),
.A3(n_499),
.B(n_500),
.Y(n_3886)
);

AO31x2_ASAP7_75t_L g3887 ( 
.A1(n_3710),
.A2(n_502),
.A3(n_499),
.B(n_500),
.Y(n_3887)
);

O2A1O1Ixp33_ASAP7_75t_L g3888 ( 
.A1(n_3529),
.A2(n_502),
.B(n_499),
.C(n_500),
.Y(n_3888)
);

BUFx10_ASAP7_75t_L g3889 ( 
.A(n_3258),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3421),
.B(n_503),
.Y(n_3890)
);

CKINVDCx20_ASAP7_75t_R g3891 ( 
.A(n_3250),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3412),
.Y(n_3892)
);

NOR2xp33_ASAP7_75t_L g3893 ( 
.A(n_3443),
.B(n_503),
.Y(n_3893)
);

OR2x2_ASAP7_75t_L g3894 ( 
.A(n_3368),
.B(n_503),
.Y(n_3894)
);

OAI21x1_ASAP7_75t_L g3895 ( 
.A1(n_3749),
.A2(n_506),
.B(n_505),
.Y(n_3895)
);

AOI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3693),
.A2(n_504),
.B(n_505),
.Y(n_3896)
);

OAI21x1_ASAP7_75t_L g3897 ( 
.A1(n_3747),
.A2(n_506),
.B(n_505),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3607),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_3563),
.A2(n_504),
.B(n_506),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3418),
.Y(n_3900)
);

A2O1A1Ixp33_ASAP7_75t_L g3901 ( 
.A1(n_3706),
.A2(n_508),
.B(n_504),
.C(n_507),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3648),
.Y(n_3902)
);

INVx3_ASAP7_75t_L g3903 ( 
.A(n_3387),
.Y(n_3903)
);

CKINVDCx6p67_ASAP7_75t_R g3904 ( 
.A(n_3233),
.Y(n_3904)
);

INVx3_ASAP7_75t_L g3905 ( 
.A(n_3273),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3316),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3575),
.A2(n_507),
.B(n_508),
.Y(n_3907)
);

AOI21x1_ASAP7_75t_L g3908 ( 
.A1(n_3535),
.A2(n_556),
.B(n_555),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3582),
.A2(n_507),
.B(n_509),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3313),
.B(n_509),
.Y(n_3910)
);

OR2x2_ASAP7_75t_L g3911 ( 
.A(n_3313),
.B(n_509),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3283),
.B(n_3677),
.Y(n_3912)
);

OAI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3280),
.A2(n_3605),
.B(n_3695),
.Y(n_3913)
);

O2A1O1Ixp33_ASAP7_75t_SL g3914 ( 
.A1(n_3315),
.A2(n_512),
.B(n_510),
.C(n_511),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3502),
.Y(n_3915)
);

O2A1O1Ixp33_ASAP7_75t_L g3916 ( 
.A1(n_3560),
.A2(n_512),
.B(n_510),
.C(n_511),
.Y(n_3916)
);

O2A1O1Ixp33_ASAP7_75t_SL g3917 ( 
.A1(n_3240),
.A2(n_514),
.B(n_510),
.C(n_513),
.Y(n_3917)
);

AO31x2_ASAP7_75t_L g3918 ( 
.A1(n_3294),
.A2(n_515),
.A3(n_513),
.B(n_514),
.Y(n_3918)
);

OAI21x1_ASAP7_75t_L g3919 ( 
.A1(n_3612),
.A2(n_515),
.B(n_514),
.Y(n_3919)
);

BUFx3_ASAP7_75t_L g3920 ( 
.A(n_3441),
.Y(n_3920)
);

BUFx3_ASAP7_75t_L g3921 ( 
.A(n_3483),
.Y(n_3921)
);

O2A1O1Ixp33_ASAP7_75t_SL g3922 ( 
.A1(n_3332),
.A2(n_516),
.B(n_513),
.C(n_515),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_SL g3923 ( 
.A(n_3222),
.B(n_517),
.Y(n_3923)
);

O2A1O1Ixp33_ASAP7_75t_SL g3924 ( 
.A1(n_3537),
.A2(n_519),
.B(n_517),
.C(n_518),
.Y(n_3924)
);

A2O1A1Ixp33_ASAP7_75t_L g3925 ( 
.A1(n_3721),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_3925)
);

INVx3_ASAP7_75t_R g3926 ( 
.A(n_3477),
.Y(n_3926)
);

AOI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3593),
.A2(n_519),
.B(n_520),
.Y(n_3927)
);

INVx3_ASAP7_75t_L g3928 ( 
.A(n_3273),
.Y(n_3928)
);

AOI22xp5_ASAP7_75t_L g3929 ( 
.A1(n_3613),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_3929)
);

OAI21x1_ASAP7_75t_L g3930 ( 
.A1(n_3447),
.A2(n_525),
.B(n_524),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3712),
.B(n_521),
.Y(n_3931)
);

INVx5_ASAP7_75t_L g3932 ( 
.A(n_3394),
.Y(n_3932)
);

HB1xp67_ASAP7_75t_L g3933 ( 
.A(n_3485),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3230),
.B(n_521),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3507),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_3699),
.B(n_524),
.Y(n_3936)
);

A2O1A1Ixp33_ASAP7_75t_L g3937 ( 
.A1(n_3231),
.A2(n_525),
.B(n_556),
.C(n_555),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3594),
.A2(n_557),
.B(n_558),
.Y(n_3938)
);

OAI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3372),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_3939)
);

AND2x4_ASAP7_75t_L g3940 ( 
.A(n_3372),
.B(n_559),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3410),
.B(n_560),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3550),
.B(n_560),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3526),
.Y(n_3943)
);

OAI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_3656),
.A2(n_561),
.B(n_562),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3596),
.A2(n_561),
.B(n_563),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3681),
.A2(n_563),
.B(n_564),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3373),
.Y(n_3947)
);

OAI21x1_ASAP7_75t_L g3948 ( 
.A1(n_3447),
.A2(n_564),
.B(n_565),
.Y(n_3948)
);

AOI211x1_ASAP7_75t_L g3949 ( 
.A1(n_3225),
.A2(n_567),
.B(n_565),
.C(n_566),
.Y(n_3949)
);

AOI21x1_ASAP7_75t_L g3950 ( 
.A1(n_3335),
.A2(n_566),
.B(n_568),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_3474),
.A2(n_568),
.B(n_569),
.Y(n_3951)
);

A2O1A1Ixp33_ASAP7_75t_L g3952 ( 
.A1(n_3326),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3373),
.B(n_3450),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3251),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3499),
.B(n_570),
.Y(n_3955)
);

OAI21x1_ASAP7_75t_L g3956 ( 
.A1(n_3456),
.A2(n_3374),
.B(n_3276),
.Y(n_3956)
);

NOR2xp33_ASAP7_75t_L g3957 ( 
.A(n_3673),
.B(n_3438),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3268),
.Y(n_3958)
);

AO31x2_ASAP7_75t_L g3959 ( 
.A1(n_3312),
.A2(n_573),
.A3(n_571),
.B(n_572),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3436),
.B(n_574),
.Y(n_3960)
);

AO21x1_ASAP7_75t_L g3961 ( 
.A1(n_3678),
.A2(n_574),
.B(n_576),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3484),
.B(n_576),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3295),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3247),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3491),
.A2(n_577),
.B(n_578),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3503),
.B(n_961),
.Y(n_3966)
);

AOI22xp33_ASAP7_75t_L g3967 ( 
.A1(n_3559),
.A2(n_580),
.B1(n_577),
.B2(n_579),
.Y(n_3967)
);

BUFx2_ASAP7_75t_L g3968 ( 
.A(n_3514),
.Y(n_3968)
);

O2A1O1Ixp33_ASAP7_75t_SL g3969 ( 
.A1(n_3551),
.A2(n_582),
.B(n_580),
.C(n_581),
.Y(n_3969)
);

CKINVDCx5p33_ASAP7_75t_R g3970 ( 
.A(n_3343),
.Y(n_3970)
);

BUFx12f_ASAP7_75t_L g3971 ( 
.A(n_3434),
.Y(n_3971)
);

HB1xp67_ASAP7_75t_L g3972 ( 
.A(n_3375),
.Y(n_3972)
);

OAI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3419),
.A2(n_581),
.B(n_582),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3503),
.B(n_583),
.Y(n_3974)
);

AO31x2_ASAP7_75t_L g3975 ( 
.A1(n_3320),
.A2(n_586),
.A3(n_583),
.B(n_584),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3674),
.B(n_961),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3380),
.B(n_3414),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3510),
.A2(n_584),
.B(n_586),
.Y(n_3978)
);

AO31x2_ASAP7_75t_L g3979 ( 
.A1(n_3339),
.A2(n_3344),
.A3(n_3376),
.B(n_3574),
.Y(n_3979)
);

OAI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_3542),
.A2(n_588),
.B(n_589),
.Y(n_3980)
);

AOI21xp5_ASAP7_75t_L g3981 ( 
.A1(n_3521),
.A2(n_588),
.B(n_590),
.Y(n_3981)
);

OA21x2_ASAP7_75t_L g3982 ( 
.A1(n_3318),
.A2(n_590),
.B(n_591),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3449),
.B(n_960),
.Y(n_3983)
);

OAI22xp5_ASAP7_75t_L g3984 ( 
.A1(n_3654),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3501),
.A2(n_592),
.B(n_594),
.Y(n_3985)
);

OAI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3279),
.A2(n_597),
.B1(n_594),
.B2(n_595),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3466),
.B(n_595),
.Y(n_3987)
);

NOR2xp33_ASAP7_75t_L g3988 ( 
.A(n_3520),
.B(n_598),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3585),
.B(n_599),
.Y(n_3989)
);

OAI22x1_ASAP7_75t_L g3990 ( 
.A1(n_3404),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_3990)
);

AOI22xp33_ASAP7_75t_L g3991 ( 
.A1(n_3559),
.A2(n_604),
.B1(n_600),
.B2(n_603),
.Y(n_3991)
);

OAI21xp5_ASAP7_75t_L g3992 ( 
.A1(n_3516),
.A2(n_604),
.B(n_605),
.Y(n_3992)
);

OAI21x1_ASAP7_75t_L g3993 ( 
.A1(n_3456),
.A2(n_605),
.B(n_606),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3265),
.Y(n_3994)
);

AOI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3579),
.A2(n_607),
.B(n_608),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3659),
.B(n_960),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3298),
.Y(n_3997)
);

O2A1O1Ixp33_ASAP7_75t_SL g3998 ( 
.A1(n_3591),
.A2(n_610),
.B(n_607),
.C(n_609),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3300),
.Y(n_3999)
);

OAI22xp5_ASAP7_75t_L g4000 ( 
.A1(n_3291),
.A2(n_612),
.B1(n_610),
.B2(n_611),
.Y(n_4000)
);

A2O1A1Ixp33_ASAP7_75t_L g4001 ( 
.A1(n_3228),
.A2(n_613),
.B(n_611),
.C(n_612),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3303),
.Y(n_4002)
);

AOI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3604),
.A2(n_613),
.B(n_614),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3307),
.Y(n_4004)
);

CKINVDCx20_ASAP7_75t_R g4005 ( 
.A(n_3588),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3244),
.B(n_615),
.Y(n_4006)
);

OAI21xp33_ASAP7_75t_L g4007 ( 
.A1(n_3543),
.A2(n_615),
.B(n_616),
.Y(n_4007)
);

OAI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3354),
.A2(n_616),
.B(n_618),
.Y(n_4008)
);

OAI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3480),
.A2(n_618),
.B(n_619),
.Y(n_4009)
);

OAI21x1_ASAP7_75t_L g4010 ( 
.A1(n_3274),
.A2(n_619),
.B(n_620),
.Y(n_4010)
);

INVxp67_ASAP7_75t_SL g4011 ( 
.A(n_3739),
.Y(n_4011)
);

BUFx8_ASAP7_75t_SL g4012 ( 
.A(n_3342),
.Y(n_4012)
);

INVxp67_ASAP7_75t_L g4013 ( 
.A(n_3328),
.Y(n_4013)
);

HB1xp67_ASAP7_75t_L g4014 ( 
.A(n_3492),
.Y(n_4014)
);

OAI21x1_ASAP7_75t_L g4015 ( 
.A1(n_3274),
.A2(n_621),
.B(n_622),
.Y(n_4015)
);

AOI21x1_ASAP7_75t_L g4016 ( 
.A1(n_3335),
.A2(n_621),
.B(n_622),
.Y(n_4016)
);

INVx2_ASAP7_75t_SL g4017 ( 
.A(n_3345),
.Y(n_4017)
);

OAI21x1_ASAP7_75t_L g4018 ( 
.A1(n_3276),
.A2(n_623),
.B(n_624),
.Y(n_4018)
);

AOI221xp5_ASAP7_75t_SL g4019 ( 
.A1(n_3364),
.A2(n_626),
.B1(n_623),
.B2(n_625),
.C(n_627),
.Y(n_4019)
);

AND2x2_ASAP7_75t_SL g4020 ( 
.A(n_3739),
.B(n_625),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3665),
.A2(n_3676),
.B(n_3624),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3664),
.B(n_626),
.Y(n_4022)
);

O2A1O1Ixp33_ASAP7_75t_L g4023 ( 
.A1(n_3544),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_3608),
.A2(n_628),
.B(n_629),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3310),
.Y(n_4025)
);

O2A1O1Ixp33_ASAP7_75t_SL g4026 ( 
.A1(n_3509),
.A2(n_632),
.B(n_630),
.C(n_631),
.Y(n_4026)
);

AO31x2_ASAP7_75t_L g4027 ( 
.A1(n_3670),
.A2(n_634),
.A3(n_632),
.B(n_633),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_3631),
.A2(n_3641),
.B(n_3638),
.Y(n_4028)
);

CKINVDCx16_ASAP7_75t_R g4029 ( 
.A(n_3386),
.Y(n_4029)
);

OAI21x1_ASAP7_75t_L g4030 ( 
.A1(n_3351),
.A2(n_633),
.B(n_634),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3269),
.B(n_635),
.Y(n_4031)
);

BUFx3_ASAP7_75t_L g4032 ( 
.A(n_3470),
.Y(n_4032)
);

OAI21x1_ASAP7_75t_L g4033 ( 
.A1(n_3282),
.A2(n_635),
.B(n_636),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3420),
.B(n_959),
.Y(n_4034)
);

BUFx12f_ASAP7_75t_L g4035 ( 
.A(n_3698),
.Y(n_4035)
);

HB1xp67_ASAP7_75t_L g4036 ( 
.A(n_3614),
.Y(n_4036)
);

A2O1A1Ixp33_ASAP7_75t_L g4037 ( 
.A1(n_3518),
.A2(n_638),
.B(n_636),
.C(n_637),
.Y(n_4037)
);

O2A1O1Ixp33_ASAP7_75t_SL g4038 ( 
.A1(n_3554),
.A2(n_640),
.B(n_637),
.C(n_639),
.Y(n_4038)
);

CKINVDCx20_ASAP7_75t_R g4039 ( 
.A(n_3262),
.Y(n_4039)
);

A2O1A1Ixp33_ASAP7_75t_L g4040 ( 
.A1(n_3702),
.A2(n_644),
.B(n_642),
.C(n_643),
.Y(n_4040)
);

AO31x2_ASAP7_75t_L g4041 ( 
.A1(n_3603),
.A2(n_645),
.A3(n_642),
.B(n_644),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3475),
.B(n_959),
.Y(n_4042)
);

AOI21x1_ASAP7_75t_L g4043 ( 
.A1(n_3617),
.A2(n_645),
.B(n_646),
.Y(n_4043)
);

AOI22xp33_ASAP7_75t_L g4044 ( 
.A1(n_3556),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_4044)
);

INVx3_ASAP7_75t_SL g4045 ( 
.A(n_3609),
.Y(n_4045)
);

OAI21x1_ASAP7_75t_L g4046 ( 
.A1(n_3296),
.A2(n_648),
.B(n_649),
.Y(n_4046)
);

OAI21x1_ASAP7_75t_L g4047 ( 
.A1(n_3341),
.A2(n_650),
.B(n_651),
.Y(n_4047)
);

AO31x2_ASAP7_75t_L g4048 ( 
.A1(n_3700),
.A2(n_653),
.A3(n_651),
.B(n_652),
.Y(n_4048)
);

AND2x4_ASAP7_75t_L g4049 ( 
.A(n_3371),
.B(n_958),
.Y(n_4049)
);

OAI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_3586),
.A2(n_654),
.B(n_655),
.Y(n_4050)
);

O2A1O1Ixp33_ASAP7_75t_L g4051 ( 
.A1(n_3346),
.A2(n_658),
.B(n_654),
.C(n_657),
.Y(n_4051)
);

AOI221x1_ASAP7_75t_L g4052 ( 
.A1(n_3512),
.A2(n_660),
.B1(n_657),
.B2(n_659),
.C(n_661),
.Y(n_4052)
);

AOI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3398),
.A2(n_659),
.B(n_660),
.Y(n_4053)
);

INVx3_ASAP7_75t_L g4054 ( 
.A(n_3536),
.Y(n_4054)
);

NOR2xp33_ASAP7_75t_L g4055 ( 
.A(n_3369),
.B(n_661),
.Y(n_4055)
);

OAI21x1_ASAP7_75t_L g4056 ( 
.A1(n_3288),
.A2(n_662),
.B(n_663),
.Y(n_4056)
);

AOI21xp5_ASAP7_75t_L g4057 ( 
.A1(n_3666),
.A2(n_663),
.B(n_664),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3429),
.B(n_664),
.Y(n_4058)
);

AO31x2_ASAP7_75t_L g4059 ( 
.A1(n_3333),
.A2(n_667),
.A3(n_665),
.B(n_666),
.Y(n_4059)
);

AOI21xp5_ASAP7_75t_L g4060 ( 
.A1(n_3669),
.A2(n_665),
.B(n_668),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3500),
.B(n_957),
.Y(n_4061)
);

A2O1A1Ixp33_ASAP7_75t_L g4062 ( 
.A1(n_3385),
.A2(n_670),
.B(n_668),
.C(n_669),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3317),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3513),
.B(n_670),
.Y(n_4064)
);

CKINVDCx6p67_ASAP7_75t_R g4065 ( 
.A(n_3329),
.Y(n_4065)
);

OAI21xp5_ASAP7_75t_L g4066 ( 
.A1(n_3353),
.A2(n_671),
.B(n_672),
.Y(n_4066)
);

INVx3_ASAP7_75t_L g4067 ( 
.A(n_3635),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3272),
.Y(n_4068)
);

INVx2_ASAP7_75t_SL g4069 ( 
.A(n_3690),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3299),
.Y(n_4070)
);

INVxp67_ASAP7_75t_SL g4071 ( 
.A(n_3614),
.Y(n_4071)
);

NOR2xp33_ASAP7_75t_L g4072 ( 
.A(n_3458),
.B(n_3462),
.Y(n_4072)
);

AOI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_3707),
.A2(n_3668),
.B(n_3657),
.Y(n_4073)
);

INVx1_ASAP7_75t_SL g4074 ( 
.A(n_3682),
.Y(n_4074)
);

INVx3_ASAP7_75t_SL g4075 ( 
.A(n_3377),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3687),
.A2(n_671),
.B(n_673),
.Y(n_4076)
);

INVx1_ASAP7_75t_SL g4077 ( 
.A(n_3757),
.Y(n_4077)
);

INVx4_ASAP7_75t_L g4078 ( 
.A(n_3786),
.Y(n_4078)
);

CKINVDCx11_ASAP7_75t_R g4079 ( 
.A(n_3790),
.Y(n_4079)
);

BUFx12f_ASAP7_75t_L g4080 ( 
.A(n_3855),
.Y(n_4080)
);

BUFx2_ASAP7_75t_L g4081 ( 
.A(n_3882),
.Y(n_4081)
);

CKINVDCx11_ASAP7_75t_R g4082 ( 
.A(n_3806),
.Y(n_4082)
);

NAND2x1p5_ASAP7_75t_L g4083 ( 
.A(n_3932),
.B(n_3697),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3764),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_3817),
.A2(n_3833),
.B1(n_4020),
.B2(n_3756),
.Y(n_4085)
);

INVx3_ASAP7_75t_L g4086 ( 
.A(n_3838),
.Y(n_4086)
);

OAI21xp5_ASAP7_75t_SL g4087 ( 
.A1(n_3968),
.A2(n_3347),
.B(n_3565),
.Y(n_4087)
);

INVx3_ASAP7_75t_L g4088 ( 
.A(n_4035),
.Y(n_4088)
);

INVx3_ASAP7_75t_SL g4089 ( 
.A(n_3891),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_4039),
.A2(n_3724),
.B1(n_3667),
.B2(n_3600),
.Y(n_4090)
);

BUFx2_ASAP7_75t_SL g4091 ( 
.A(n_3800),
.Y(n_4091)
);

OAI22xp5_ASAP7_75t_L g4092 ( 
.A1(n_3932),
.A2(n_3566),
.B1(n_3497),
.B2(n_3395),
.Y(n_4092)
);

INVxp67_ASAP7_75t_SL g4093 ( 
.A(n_4011),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3906),
.B(n_3490),
.Y(n_4094)
);

INVx4_ASAP7_75t_L g4095 ( 
.A(n_3874),
.Y(n_4095)
);

CKINVDCx11_ASAP7_75t_R g4096 ( 
.A(n_3855),
.Y(n_4096)
);

AOI22xp33_ASAP7_75t_L g4097 ( 
.A1(n_3874),
.A2(n_3701),
.B1(n_3628),
.B2(n_3730),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3773),
.Y(n_4098)
);

INVx4_ASAP7_75t_L g4099 ( 
.A(n_3784),
.Y(n_4099)
);

AOI22xp33_ASAP7_75t_SL g4100 ( 
.A1(n_3932),
.A2(n_3708),
.B1(n_3297),
.B2(n_3626),
.Y(n_4100)
);

AOI22xp33_ASAP7_75t_SL g4101 ( 
.A1(n_3923),
.A2(n_3297),
.B1(n_3686),
.B2(n_3680),
.Y(n_4101)
);

INVx6_ASAP7_75t_L g4102 ( 
.A(n_3889),
.Y(n_4102)
);

AO22x1_ASAP7_75t_L g4103 ( 
.A1(n_3819),
.A2(n_3428),
.B1(n_3330),
.B2(n_3439),
.Y(n_4103)
);

OAI22xp5_ASAP7_75t_L g4104 ( 
.A1(n_4071),
.A2(n_3334),
.B1(n_3437),
.B2(n_3445),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3876),
.A2(n_3557),
.B1(n_3451),
.B2(n_3224),
.Y(n_4105)
);

AOI22xp33_ASAP7_75t_L g4106 ( 
.A1(n_3801),
.A2(n_3766),
.B1(n_3876),
.B2(n_4055),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3791),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_3836),
.A2(n_3446),
.B1(n_3752),
.B2(n_3713),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3871),
.B(n_3547),
.Y(n_4109)
);

CKINVDCx6p67_ASAP7_75t_R g4110 ( 
.A(n_4045),
.Y(n_4110)
);

AOI22xp33_ASAP7_75t_L g4111 ( 
.A1(n_3953),
.A2(n_3401),
.B1(n_3636),
.B2(n_3595),
.Y(n_4111)
);

INVx6_ASAP7_75t_L g4112 ( 
.A(n_3920),
.Y(n_4112)
);

OAI22xp33_ASAP7_75t_L g4113 ( 
.A1(n_3904),
.A2(n_3598),
.B1(n_3644),
.B2(n_3223),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3812),
.A2(n_3639),
.B1(n_3646),
.B2(n_3738),
.Y(n_4114)
);

AOI22xp33_ASAP7_75t_L g4115 ( 
.A1(n_4065),
.A2(n_3740),
.B1(n_3743),
.B2(n_3572),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3807),
.Y(n_4116)
);

INVx6_ASAP7_75t_L g4117 ( 
.A(n_3815),
.Y(n_4117)
);

BUFx8_ASAP7_75t_SL g4118 ( 
.A(n_3971),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3898),
.Y(n_4119)
);

BUFx6f_ASAP7_75t_L g4120 ( 
.A(n_3921),
.Y(n_4120)
);

CKINVDCx20_ASAP7_75t_R g4121 ( 
.A(n_4012),
.Y(n_4121)
);

OAI21xp5_ASAP7_75t_SL g4122 ( 
.A1(n_4013),
.A2(n_3616),
.B(n_3570),
.Y(n_4122)
);

CKINVDCx11_ASAP7_75t_R g4123 ( 
.A(n_4005),
.Y(n_4123)
);

INVx1_ASAP7_75t_SL g4124 ( 
.A(n_4075),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_3902),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3964),
.Y(n_4126)
);

INVx1_ASAP7_75t_SL g4127 ( 
.A(n_3903),
.Y(n_4127)
);

AOI22xp33_ASAP7_75t_SL g4128 ( 
.A1(n_3940),
.A2(n_3671),
.B1(n_3622),
.B2(n_3602),
.Y(n_4128)
);

OAI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_3862),
.A2(n_3549),
.B1(n_3629),
.B2(n_3732),
.Y(n_4129)
);

OAI22xp5_ASAP7_75t_L g4130 ( 
.A1(n_3856),
.A2(n_3741),
.B1(n_3621),
.B2(n_3473),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3808),
.Y(n_4131)
);

BUFx6f_ASAP7_75t_L g4132 ( 
.A(n_4032),
.Y(n_4132)
);

INVx1_ASAP7_75t_SL g4133 ( 
.A(n_3846),
.Y(n_4133)
);

INVx1_ASAP7_75t_SL g4134 ( 
.A(n_3809),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_3813),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3829),
.Y(n_4136)
);

BUFx3_ASAP7_75t_L g4137 ( 
.A(n_3845),
.Y(n_4137)
);

INVxp67_ASAP7_75t_SL g4138 ( 
.A(n_4036),
.Y(n_4138)
);

OR2x2_ASAP7_75t_L g4139 ( 
.A(n_3854),
.B(n_3553),
.Y(n_4139)
);

CKINVDCx5p33_ASAP7_75t_R g4140 ( 
.A(n_3970),
.Y(n_4140)
);

NAND2x1p5_ASAP7_75t_L g4141 ( 
.A(n_3789),
.B(n_3689),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_3830),
.Y(n_4142)
);

INVx4_ASAP7_75t_L g4143 ( 
.A(n_4054),
.Y(n_4143)
);

BUFx12f_ASAP7_75t_L g4144 ( 
.A(n_4017),
.Y(n_4144)
);

OAI22xp5_ASAP7_75t_L g4145 ( 
.A1(n_3925),
.A2(n_3405),
.B1(n_3393),
.B2(n_3623),
.Y(n_4145)
);

OAI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_3822),
.A2(n_3675),
.B1(n_3625),
.B2(n_3746),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_3860),
.A2(n_3799),
.B1(n_3783),
.B2(n_3831),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3865),
.Y(n_4148)
);

INVx6_ASAP7_75t_L g4149 ( 
.A(n_4029),
.Y(n_4149)
);

OAI22xp5_ASAP7_75t_L g4150 ( 
.A1(n_3770),
.A2(n_3851),
.B1(n_3911),
.B2(n_3792),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3892),
.Y(n_4151)
);

INVx1_ASAP7_75t_SL g4152 ( 
.A(n_4014),
.Y(n_4152)
);

BUFx12f_ASAP7_75t_L g4153 ( 
.A(n_4069),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3900),
.B(n_3406),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3853),
.Y(n_4155)
);

BUFx6f_ASAP7_75t_L g4156 ( 
.A(n_4067),
.Y(n_4156)
);

AOI22xp33_ASAP7_75t_L g4157 ( 
.A1(n_4007),
.A2(n_3658),
.B1(n_3264),
.B2(n_3643),
.Y(n_4157)
);

OAI22xp5_ASAP7_75t_L g4158 ( 
.A1(n_3980),
.A2(n_3748),
.B1(n_3232),
.B2(n_3246),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_3994),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_3910),
.B(n_3377),
.Y(n_4160)
);

OAI21xp5_ASAP7_75t_L g4161 ( 
.A1(n_3779),
.A2(n_3879),
.B(n_4028),
.Y(n_4161)
);

OAI22xp5_ASAP7_75t_L g4162 ( 
.A1(n_3992),
.A2(n_4009),
.B1(n_3944),
.B2(n_3991),
.Y(n_4162)
);

OAI22x1_ASAP7_75t_L g4163 ( 
.A1(n_3821),
.A2(n_3261),
.B1(n_3289),
.B2(n_3286),
.Y(n_4163)
);

BUFx12f_ASAP7_75t_L g4164 ( 
.A(n_4049),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_4068),
.Y(n_4165)
);

BUFx6f_ASAP7_75t_L g4166 ( 
.A(n_3905),
.Y(n_4166)
);

BUFx3_ASAP7_75t_L g4167 ( 
.A(n_3933),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3915),
.Y(n_4168)
);

INVxp67_ASAP7_75t_SL g4169 ( 
.A(n_3972),
.Y(n_4169)
);

OAI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_3967),
.A2(n_3487),
.B1(n_3627),
.B2(n_3517),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3935),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_4070),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3943),
.Y(n_4173)
);

CKINVDCx6p67_ASAP7_75t_R g4174 ( 
.A(n_3926),
.Y(n_4174)
);

BUFx6f_ASAP7_75t_L g4175 ( 
.A(n_3928),
.Y(n_4175)
);

INVx6_ASAP7_75t_L g4176 ( 
.A(n_3762),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_SL g4177 ( 
.A1(n_3804),
.A2(n_3709),
.B1(n_3302),
.B2(n_3319),
.Y(n_4177)
);

CKINVDCx6p67_ASAP7_75t_R g4178 ( 
.A(n_3990),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3912),
.B(n_3396),
.Y(n_4179)
);

AOI22xp33_ASAP7_75t_L g4180 ( 
.A1(n_4006),
.A2(n_3362),
.B1(n_3744),
.B2(n_3304),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3788),
.Y(n_4181)
);

AOI21xp33_ASAP7_75t_L g4182 ( 
.A1(n_3769),
.A2(n_3647),
.B(n_3416),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_L g4183 ( 
.A1(n_4072),
.A2(n_3652),
.B1(n_3599),
.B2(n_3360),
.Y(n_4183)
);

OAI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_3952),
.A2(n_3355),
.B1(n_3361),
.B2(n_3718),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_3843),
.Y(n_4185)
);

AOI22xp33_ASAP7_75t_L g4186 ( 
.A1(n_3947),
.A2(n_4058),
.B1(n_3893),
.B2(n_4000),
.Y(n_4186)
);

INVx3_ASAP7_75t_L g4187 ( 
.A(n_4074),
.Y(n_4187)
);

AOI22xp5_ASAP7_75t_L g4188 ( 
.A1(n_3936),
.A2(n_3661),
.B1(n_3528),
.B2(n_3531),
.Y(n_4188)
);

BUFx6f_ASAP7_75t_L g4189 ( 
.A(n_3868),
.Y(n_4189)
);

INVx6_ASAP7_75t_L g4190 ( 
.A(n_3960),
.Y(n_4190)
);

CKINVDCx11_ASAP7_75t_R g4191 ( 
.A(n_3873),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3930),
.Y(n_4192)
);

OAI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_4021),
.A2(n_3840),
.B(n_3937),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_3883),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3954),
.B(n_3249),
.Y(n_4195)
);

BUFx2_ASAP7_75t_L g4196 ( 
.A(n_3885),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_3977),
.B(n_3894),
.Y(n_4197)
);

BUFx8_ASAP7_75t_L g4198 ( 
.A(n_3958),
.Y(n_4198)
);

CKINVDCx6p67_ASAP7_75t_R g4199 ( 
.A(n_3827),
.Y(n_4199)
);

AOI22xp33_ASAP7_75t_SL g4200 ( 
.A1(n_3984),
.A2(n_3302),
.B1(n_3319),
.B2(n_3288),
.Y(n_4200)
);

CKINVDCx11_ASAP7_75t_R g4201 ( 
.A(n_3872),
.Y(n_4201)
);

BUFx12f_ASAP7_75t_L g4202 ( 
.A(n_3957),
.Y(n_4202)
);

BUFx10_ASAP7_75t_L g4203 ( 
.A(n_3988),
.Y(n_4203)
);

OAI22xp5_ASAP7_75t_L g4204 ( 
.A1(n_3844),
.A2(n_3435),
.B1(n_3524),
.B2(n_3534),
.Y(n_4204)
);

BUFx10_ASAP7_75t_L g4205 ( 
.A(n_3963),
.Y(n_4205)
);

NAND2x1p5_ASAP7_75t_L g4206 ( 
.A(n_3948),
.B(n_3717),
.Y(n_4206)
);

BUFx3_ASAP7_75t_L g4207 ( 
.A(n_3976),
.Y(n_4207)
);

CKINVDCx20_ASAP7_75t_R g4208 ( 
.A(n_3929),
.Y(n_4208)
);

BUFx6f_ASAP7_75t_L g4209 ( 
.A(n_3787),
.Y(n_4209)
);

AOI22xp33_ASAP7_75t_L g4210 ( 
.A1(n_3986),
.A2(n_3754),
.B1(n_3736),
.B2(n_3391),
.Y(n_4210)
);

CKINVDCx20_ASAP7_75t_R g4211 ( 
.A(n_3955),
.Y(n_4211)
);

BUFx3_ASAP7_75t_L g4212 ( 
.A(n_3993),
.Y(n_4212)
);

OAI22xp33_ASAP7_75t_L g4213 ( 
.A1(n_3939),
.A2(n_3378),
.B1(n_3383),
.B2(n_3349),
.Y(n_4213)
);

INVx3_ASAP7_75t_L g4214 ( 
.A(n_4010),
.Y(n_4214)
);

BUFx12f_ASAP7_75t_L g4215 ( 
.A(n_3949),
.Y(n_4215)
);

INVx1_ASAP7_75t_SL g4216 ( 
.A(n_3966),
.Y(n_4216)
);

CKINVDCx20_ASAP7_75t_R g4217 ( 
.A(n_3983),
.Y(n_4217)
);

INVx6_ASAP7_75t_L g4218 ( 
.A(n_3768),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3852),
.Y(n_4219)
);

OAI22xp5_ASAP7_75t_L g4220 ( 
.A1(n_3858),
.A2(n_3541),
.B1(n_3482),
.B2(n_3493),
.Y(n_4220)
);

INVx2_ASAP7_75t_SL g4221 ( 
.A(n_3974),
.Y(n_4221)
);

INVx6_ASAP7_75t_L g4222 ( 
.A(n_3922),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_3895),
.Y(n_4223)
);

BUFx3_ASAP7_75t_L g4224 ( 
.A(n_4015),
.Y(n_4224)
);

NAND2x1p5_ASAP7_75t_L g4225 ( 
.A(n_4018),
.B(n_3496),
.Y(n_4225)
);

AOI22xp33_ASAP7_75t_L g4226 ( 
.A1(n_3767),
.A2(n_3461),
.B1(n_3472),
.B2(n_3455),
.Y(n_4226)
);

CKINVDCx11_ASAP7_75t_R g4227 ( 
.A(n_3997),
.Y(n_4227)
);

BUFx2_ASAP7_75t_L g4228 ( 
.A(n_3987),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_SL g4229 ( 
.A1(n_3973),
.A2(n_3532),
.B1(n_3555),
.B2(n_3496),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4056),
.Y(n_4230)
);

INVx2_ASAP7_75t_L g4231 ( 
.A(n_3950),
.Y(n_4231)
);

BUFx6f_ASAP7_75t_L g4232 ( 
.A(n_3956),
.Y(n_4232)
);

HB1xp67_ASAP7_75t_L g4233 ( 
.A(n_3931),
.Y(n_4233)
);

OAI22xp5_ASAP7_75t_L g4234 ( 
.A1(n_3818),
.A2(n_3452),
.B1(n_3423),
.B2(n_3448),
.Y(n_4234)
);

OAI22xp33_ASAP7_75t_L g4235 ( 
.A1(n_3989),
.A2(n_3425),
.B1(n_3722),
.B2(n_3711),
.Y(n_4235)
);

INVx6_ASAP7_75t_L g4236 ( 
.A(n_3884),
.Y(n_4236)
);

HB1xp67_ASAP7_75t_L g4237 ( 
.A(n_3962),
.Y(n_4237)
);

INVx4_ASAP7_75t_L g4238 ( 
.A(n_3982),
.Y(n_4238)
);

AOI22xp33_ASAP7_75t_L g4239 ( 
.A1(n_3913),
.A2(n_3506),
.B1(n_3527),
.B2(n_3498),
.Y(n_4239)
);

AOI22xp33_ASAP7_75t_L g4240 ( 
.A1(n_3802),
.A2(n_3561),
.B1(n_3562),
.B2(n_3546),
.Y(n_4240)
);

INVx6_ASAP7_75t_L g4241 ( 
.A(n_3917),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_3941),
.B(n_3606),
.Y(n_4242)
);

OAI22xp33_ASAP7_75t_L g4243 ( 
.A1(n_4034),
.A2(n_3684),
.B1(n_3569),
.B2(n_3555),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_L g4244 ( 
.A1(n_3890),
.A2(n_3573),
.B1(n_3577),
.B2(n_3568),
.Y(n_4244)
);

INVx2_ASAP7_75t_L g4245 ( 
.A(n_4016),
.Y(n_4245)
);

AOI22xp33_ASAP7_75t_L g4246 ( 
.A1(n_3999),
.A2(n_3589),
.B1(n_3597),
.B2(n_3583),
.Y(n_4246)
);

INVx1_ASAP7_75t_SL g4247 ( 
.A(n_3863),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_3897),
.Y(n_4248)
);

INVx1_ASAP7_75t_SL g4249 ( 
.A(n_3864),
.Y(n_4249)
);

BUFx8_ASAP7_75t_L g4250 ( 
.A(n_4002),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4004),
.B(n_3306),
.Y(n_4251)
);

INVx3_ASAP7_75t_L g4252 ( 
.A(n_3881),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_3919),
.Y(n_4253)
);

OAI22xp5_ASAP7_75t_L g4254 ( 
.A1(n_4044),
.A2(n_3753),
.B1(n_3290),
.B2(n_3442),
.Y(n_4254)
);

OAI22xp5_ASAP7_75t_L g4255 ( 
.A1(n_3870),
.A2(n_3444),
.B1(n_3464),
.B2(n_3440),
.Y(n_4255)
);

INVx6_ASAP7_75t_L g4256 ( 
.A(n_3914),
.Y(n_4256)
);

CKINVDCx14_ASAP7_75t_R g4257 ( 
.A(n_4025),
.Y(n_4257)
);

AOI22xp33_ASAP7_75t_SL g4258 ( 
.A1(n_3982),
.A2(n_3532),
.B1(n_3742),
.B2(n_3731),
.Y(n_4258)
);

BUFx3_ASAP7_75t_L g4259 ( 
.A(n_3942),
.Y(n_4259)
);

AOI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_4063),
.A2(n_3637),
.B1(n_3642),
.B2(n_3618),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_3887),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3887),
.Y(n_4262)
);

AND2x4_ASAP7_75t_L g4263 ( 
.A(n_4008),
.B(n_3716),
.Y(n_4263)
);

AOI22xp33_ASAP7_75t_L g4264 ( 
.A1(n_4066),
.A2(n_3660),
.B1(n_3411),
.B2(n_3388),
.Y(n_4264)
);

OAI21xp5_ASAP7_75t_SL g4265 ( 
.A1(n_4023),
.A2(n_3630),
.B(n_3685),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4027),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4027),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_3842),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4084),
.Y(n_4269)
);

NOR2xp33_ASAP7_75t_L g4270 ( 
.A(n_4257),
.B(n_4031),
.Y(n_4270)
);

AOI21x1_ASAP7_75t_L g4271 ( 
.A1(n_4231),
.A2(n_3816),
.B(n_3805),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4098),
.Y(n_4272)
);

HB1xp67_ASAP7_75t_L g4273 ( 
.A(n_4081),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4119),
.Y(n_4274)
);

INVx8_ASAP7_75t_L g4275 ( 
.A(n_4086),
.Y(n_4275)
);

OR2x6_ASAP7_75t_L g4276 ( 
.A(n_4091),
.B(n_4095),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4107),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4109),
.B(n_4041),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4116),
.Y(n_4279)
);

INVx3_ASAP7_75t_L g4280 ( 
.A(n_4099),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_4093),
.B(n_3841),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4131),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4135),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4136),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4125),
.Y(n_4285)
);

OAI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4085),
.A2(n_4001),
.B(n_3901),
.Y(n_4286)
);

INVx3_ASAP7_75t_L g4287 ( 
.A(n_4078),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4142),
.Y(n_4288)
);

AO21x1_ASAP7_75t_SL g4289 ( 
.A1(n_4193),
.A2(n_3859),
.B(n_3850),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4148),
.Y(n_4290)
);

OAI21x1_ASAP7_75t_L g4291 ( 
.A1(n_4161),
.A2(n_3828),
.B(n_3794),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4151),
.Y(n_4292)
);

AOI21xp5_ASAP7_75t_L g4293 ( 
.A1(n_4243),
.A2(n_3760),
.B(n_3837),
.Y(n_4293)
);

AO21x2_ASAP7_75t_L g4294 ( 
.A1(n_4245),
.A2(n_3908),
.B(n_3961),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4168),
.Y(n_4295)
);

OR2x6_ASAP7_75t_L g4296 ( 
.A(n_4149),
.B(n_3951),
.Y(n_4296)
);

OR2x2_ASAP7_75t_L g4297 ( 
.A(n_4133),
.B(n_3875),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_4167),
.Y(n_4298)
);

OAI21x1_ASAP7_75t_L g4299 ( 
.A1(n_4214),
.A2(n_3759),
.B(n_3755),
.Y(n_4299)
);

INVx3_ASAP7_75t_L g4300 ( 
.A(n_4205),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4126),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_4261),
.B(n_3841),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4159),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4171),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_4174),
.Y(n_4305)
);

OAI21x1_ASAP7_75t_L g4306 ( 
.A1(n_4225),
.A2(n_3847),
.B(n_3763),
.Y(n_4306)
);

OAI21x1_ASAP7_75t_L g4307 ( 
.A1(n_4230),
.A2(n_3761),
.B(n_3774),
.Y(n_4307)
);

AOI21xp5_ASAP7_75t_L g4308 ( 
.A1(n_4162),
.A2(n_3782),
.B(n_4073),
.Y(n_4308)
);

BUFx2_ASAP7_75t_L g4309 ( 
.A(n_4143),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4173),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4181),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4185),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4165),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4169),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4155),
.Y(n_4315)
);

AND2x4_ASAP7_75t_L g4316 ( 
.A(n_4262),
.B(n_4041),
.Y(n_4316)
);

HB1xp67_ASAP7_75t_L g4317 ( 
.A(n_4189),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4147),
.B(n_4048),
.Y(n_4318)
);

AOI22xp33_ASAP7_75t_L g4319 ( 
.A1(n_4201),
.A2(n_3857),
.B1(n_3778),
.B2(n_3798),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4172),
.Y(n_4320)
);

CKINVDCx5p33_ASAP7_75t_R g4321 ( 
.A(n_4123),
.Y(n_4321)
);

OAI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_4106),
.A2(n_3880),
.B1(n_4037),
.B2(n_4040),
.Y(n_4322)
);

CKINVDCx5p33_ASAP7_75t_R g4323 ( 
.A(n_4110),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4196),
.Y(n_4324)
);

INVx2_ASAP7_75t_L g4325 ( 
.A(n_4189),
.Y(n_4325)
);

BUFx6f_ASAP7_75t_L g4326 ( 
.A(n_4156),
.Y(n_4326)
);

HB1xp67_ASAP7_75t_L g4327 ( 
.A(n_4152),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4139),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4138),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4251),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4266),
.Y(n_4331)
);

HB1xp67_ASAP7_75t_L g4332 ( 
.A(n_4187),
.Y(n_4332)
);

HB1xp67_ASAP7_75t_L g4333 ( 
.A(n_4134),
.Y(n_4333)
);

BUFx4f_ASAP7_75t_SL g4334 ( 
.A(n_4121),
.Y(n_4334)
);

HB1xp67_ASAP7_75t_L g4335 ( 
.A(n_4233),
.Y(n_4335)
);

HB1xp67_ASAP7_75t_L g4336 ( 
.A(n_4190),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_4267),
.Y(n_4337)
);

BUFx2_ASAP7_75t_L g4338 ( 
.A(n_4112),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_4219),
.B(n_4094),
.Y(n_4339)
);

CKINVDCx11_ASAP7_75t_R g4340 ( 
.A(n_4079),
.Y(n_4340)
);

BUFx12f_ASAP7_75t_L g4341 ( 
.A(n_4082),
.Y(n_4341)
);

HB1xp67_ASAP7_75t_L g4342 ( 
.A(n_4190),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4194),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4237),
.Y(n_4344)
);

INVx2_ASAP7_75t_L g4345 ( 
.A(n_4223),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4160),
.B(n_4059),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4197),
.Y(n_4347)
);

INVx3_ASAP7_75t_L g4348 ( 
.A(n_4209),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4268),
.Y(n_4349)
);

OR2x6_ASAP7_75t_L g4350 ( 
.A(n_4149),
.B(n_3965),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4242),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4195),
.Y(n_4352)
);

OAI22xp33_ASAP7_75t_L g4353 ( 
.A1(n_4178),
.A2(n_4052),
.B1(n_3777),
.B2(n_4050),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4248),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4192),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4154),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4253),
.Y(n_4357)
);

AOI22xp33_ASAP7_75t_L g4358 ( 
.A1(n_4215),
.A2(n_3765),
.B1(n_3823),
.B2(n_3938),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4247),
.Y(n_4359)
);

INVx3_ASAP7_75t_L g4360 ( 
.A(n_4209),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4249),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4198),
.Y(n_4362)
);

INVx1_ASAP7_75t_SL g4363 ( 
.A(n_4117),
.Y(n_4363)
);

OAI21x1_ASAP7_75t_L g4364 ( 
.A1(n_4252),
.A2(n_3780),
.B(n_3776),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4250),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4238),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4212),
.Y(n_4367)
);

AND2x4_ASAP7_75t_L g4368 ( 
.A(n_4263),
.B(n_4059),
.Y(n_4368)
);

CKINVDCx11_ASAP7_75t_R g4369 ( 
.A(n_4089),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4228),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_4179),
.B(n_4048),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_4224),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4236),
.Y(n_4373)
);

BUFx2_ASAP7_75t_L g4374 ( 
.A(n_4112),
.Y(n_4374)
);

OAI21x1_ASAP7_75t_L g4375 ( 
.A1(n_4206),
.A2(n_3771),
.B(n_3775),
.Y(n_4375)
);

HB1xp67_ASAP7_75t_L g4376 ( 
.A(n_4156),
.Y(n_4376)
);

BUFx2_ASAP7_75t_L g4377 ( 
.A(n_4153),
.Y(n_4377)
);

AND2x2_ASAP7_75t_L g4378 ( 
.A(n_4216),
.B(n_4221),
.Y(n_4378)
);

AOI22xp5_ASAP7_75t_L g4379 ( 
.A1(n_4208),
.A2(n_4019),
.B1(n_3758),
.B2(n_3934),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4259),
.B(n_3996),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4236),
.Y(n_4381)
);

AND2x4_ASAP7_75t_L g4382 ( 
.A(n_4137),
.B(n_3793),
.Y(n_4382)
);

AOI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4234),
.A2(n_3772),
.B(n_3869),
.Y(n_4383)
);

OAI21x1_ASAP7_75t_L g4384 ( 
.A1(n_4255),
.A2(n_3866),
.B(n_3849),
.Y(n_4384)
);

AOI21x1_ASAP7_75t_L g4385 ( 
.A1(n_4163),
.A2(n_3832),
.B(n_4043),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4141),
.Y(n_4386)
);

INVxp33_ASAP7_75t_L g4387 ( 
.A(n_4191),
.Y(n_4387)
);

BUFx10_ASAP7_75t_L g4388 ( 
.A(n_4102),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4207),
.B(n_4227),
.Y(n_4389)
);

OAI22xp5_ASAP7_75t_L g4390 ( 
.A1(n_4097),
.A2(n_4062),
.B1(n_3985),
.B2(n_3981),
.Y(n_4390)
);

AOI22xp33_ASAP7_75t_L g4391 ( 
.A1(n_4113),
.A2(n_3946),
.B1(n_3945),
.B2(n_3899),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4127),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4176),
.Y(n_4393)
);

HB1xp67_ASAP7_75t_L g4394 ( 
.A(n_4176),
.Y(n_4394)
);

NAND3xp33_ASAP7_75t_L g4395 ( 
.A(n_4100),
.B(n_3861),
.C(n_3888),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4144),
.Y(n_4396)
);

OR2x2_ASAP7_75t_L g4397 ( 
.A(n_4077),
.B(n_4124),
.Y(n_4397)
);

AND2x2_ASAP7_75t_L g4398 ( 
.A(n_4132),
.B(n_3795),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4132),
.Y(n_4399)
);

AND2x4_ASAP7_75t_L g4400 ( 
.A(n_4309),
.B(n_4298),
.Y(n_4400)
);

NOR2x1_ASAP7_75t_R g4401 ( 
.A(n_4340),
.B(n_4323),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4351),
.B(n_4199),
.Y(n_4402)
);

AND2x4_ASAP7_75t_L g4403 ( 
.A(n_4382),
.B(n_4232),
.Y(n_4403)
);

AND2x2_ASAP7_75t_L g4404 ( 
.A(n_4273),
.B(n_4120),
.Y(n_4404)
);

INVxp67_ASAP7_75t_SL g4405 ( 
.A(n_4335),
.Y(n_4405)
);

NOR2x1_ASAP7_75t_SL g4406 ( 
.A(n_4276),
.B(n_4164),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4347),
.B(n_4120),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4274),
.Y(n_4408)
);

OAI21xp5_ASAP7_75t_L g4409 ( 
.A1(n_4383),
.A2(n_4101),
.B(n_4092),
.Y(n_4409)
);

INVxp67_ASAP7_75t_L g4410 ( 
.A(n_4327),
.Y(n_4410)
);

AND2x4_ASAP7_75t_L g4411 ( 
.A(n_4276),
.B(n_4088),
.Y(n_4411)
);

AND2x4_ASAP7_75t_L g4412 ( 
.A(n_4300),
.B(n_4166),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4344),
.Y(n_4413)
);

AND2x4_ASAP7_75t_L g4414 ( 
.A(n_4300),
.B(n_4166),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4278),
.B(n_4150),
.Y(n_4415)
);

AND2x2_ASAP7_75t_L g4416 ( 
.A(n_4378),
.B(n_4128),
.Y(n_4416)
);

AOI22xp5_ASAP7_75t_L g4417 ( 
.A1(n_4319),
.A2(n_4087),
.B1(n_4105),
.B2(n_4122),
.Y(n_4417)
);

NOR2xp67_ASAP7_75t_L g4418 ( 
.A(n_4280),
.B(n_4287),
.Y(n_4418)
);

AOI21xp5_ASAP7_75t_SL g4419 ( 
.A1(n_4373),
.A2(n_4130),
.B(n_4083),
.Y(n_4419)
);

NOR2xp33_ASAP7_75t_L g4420 ( 
.A(n_4363),
.B(n_4117),
.Y(n_4420)
);

O2A1O1Ixp33_ASAP7_75t_SL g4421 ( 
.A1(n_4362),
.A2(n_4217),
.B(n_4104),
.C(n_4213),
.Y(n_4421)
);

NOR2xp33_ASAP7_75t_L g4422 ( 
.A(n_4387),
.B(n_4202),
.Y(n_4422)
);

O2A1O1Ixp33_ASAP7_75t_SL g4423 ( 
.A1(n_4365),
.A2(n_4211),
.B(n_4170),
.C(n_4096),
.Y(n_4423)
);

AND2x2_ASAP7_75t_L g4424 ( 
.A(n_4328),
.B(n_4175),
.Y(n_4424)
);

BUFx2_ASAP7_75t_L g4425 ( 
.A(n_4382),
.Y(n_4425)
);

OAI211xp5_ASAP7_75t_L g4426 ( 
.A1(n_4286),
.A2(n_4090),
.B(n_4115),
.C(n_4114),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4324),
.B(n_4175),
.Y(n_4427)
);

OAI21x1_ASAP7_75t_SL g4428 ( 
.A1(n_4293),
.A2(n_3916),
.B(n_4053),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4314),
.B(n_4332),
.Y(n_4429)
);

NOR2xp33_ASAP7_75t_L g4430 ( 
.A(n_4369),
.B(n_4376),
.Y(n_4430)
);

NAND2xp33_ASAP7_75t_L g4431 ( 
.A(n_4275),
.B(n_4140),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4346),
.B(n_4392),
.Y(n_4432)
);

AND2x2_ASAP7_75t_L g4433 ( 
.A(n_4336),
.B(n_4203),
.Y(n_4433)
);

INVx1_ASAP7_75t_SL g4434 ( 
.A(n_4377),
.Y(n_4434)
);

NAND2x1p5_ASAP7_75t_L g4435 ( 
.A(n_4305),
.B(n_4102),
.Y(n_4435)
);

AND2x4_ASAP7_75t_L g4436 ( 
.A(n_4317),
.B(n_4232),
.Y(n_4436)
);

NOR2xp33_ASAP7_75t_L g4437 ( 
.A(n_4338),
.B(n_4080),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4342),
.B(n_4218),
.Y(n_4438)
);

AND2x4_ASAP7_75t_L g4439 ( 
.A(n_4374),
.B(n_4188),
.Y(n_4439)
);

AOI21xp5_ASAP7_75t_L g4440 ( 
.A1(n_4308),
.A2(n_4229),
.B(n_4258),
.Y(n_4440)
);

AND2x4_ASAP7_75t_L g4441 ( 
.A(n_4398),
.B(n_3886),
.Y(n_4441)
);

AND2x4_ASAP7_75t_L g4442 ( 
.A(n_4333),
.B(n_4186),
.Y(n_4442)
);

O2A1O1Ixp33_ASAP7_75t_SL g4443 ( 
.A1(n_4397),
.A2(n_4146),
.B(n_4129),
.C(n_4235),
.Y(n_4443)
);

INVx1_ASAP7_75t_SL g4444 ( 
.A(n_4388),
.Y(n_4444)
);

NOR2x1_ASAP7_75t_SL g4445 ( 
.A(n_4289),
.B(n_4145),
.Y(n_4445)
);

NAND4xp25_ASAP7_75t_L g4446 ( 
.A(n_4391),
.B(n_4108),
.C(n_4183),
.D(n_4111),
.Y(n_4446)
);

NOR2x1_ASAP7_75t_SL g4447 ( 
.A(n_4296),
.B(n_4218),
.Y(n_4447)
);

NAND2x1p5_ASAP7_75t_L g4448 ( 
.A(n_4326),
.B(n_3640),
.Y(n_4448)
);

CKINVDCx5p33_ASAP7_75t_R g4449 ( 
.A(n_4341),
.Y(n_4449)
);

AOI22xp5_ASAP7_75t_L g4450 ( 
.A1(n_4379),
.A2(n_4103),
.B1(n_4180),
.B2(n_4158),
.Y(n_4450)
);

O2A1O1Ixp33_ASAP7_75t_L g4451 ( 
.A1(n_4380),
.A2(n_4220),
.B(n_4265),
.C(n_4061),
.Y(n_4451)
);

AND2x2_ASAP7_75t_L g4452 ( 
.A(n_4370),
.B(n_4200),
.Y(n_4452)
);

HB1xp67_ASAP7_75t_L g4453 ( 
.A(n_4329),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4359),
.B(n_4177),
.Y(n_4454)
);

AO21x2_ASAP7_75t_L g4455 ( 
.A1(n_4385),
.A2(n_4182),
.B(n_3867),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4269),
.Y(n_4456)
);

BUFx10_ASAP7_75t_L g4457 ( 
.A(n_4321),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4361),
.B(n_4222),
.Y(n_4458)
);

AND2x4_ASAP7_75t_L g4459 ( 
.A(n_4325),
.B(n_4389),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4272),
.Y(n_4460)
);

AO21x2_ASAP7_75t_L g4461 ( 
.A1(n_4385),
.A2(n_4022),
.B(n_3978),
.Y(n_4461)
);

AND2x2_ASAP7_75t_L g4462 ( 
.A(n_4356),
.B(n_4222),
.Y(n_4462)
);

INVx1_ASAP7_75t_SL g4463 ( 
.A(n_4388),
.Y(n_4463)
);

AOI211xp5_ASAP7_75t_L g4464 ( 
.A1(n_4322),
.A2(n_4184),
.B(n_4204),
.C(n_4254),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4352),
.B(n_4315),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4277),
.Y(n_4466)
);

AND2x2_ASAP7_75t_L g4467 ( 
.A(n_4279),
.B(n_4241),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4282),
.B(n_4241),
.Y(n_4468)
);

OAI22xp5_ASAP7_75t_L g4469 ( 
.A1(n_4296),
.A2(n_4256),
.B1(n_4157),
.B2(n_4226),
.Y(n_4469)
);

O2A1O1Ixp33_ASAP7_75t_L g4470 ( 
.A1(n_4353),
.A2(n_4042),
.B(n_4064),
.C(n_3878),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4283),
.Y(n_4471)
);

A2O1A1Ixp33_ASAP7_75t_L g4472 ( 
.A1(n_4270),
.A2(n_3848),
.B(n_3877),
.C(n_4051),
.Y(n_4472)
);

OA21x2_ASAP7_75t_L g4473 ( 
.A1(n_4291),
.A2(n_3814),
.B(n_3781),
.Y(n_4473)
);

NOR2xp33_ASAP7_75t_L g4474 ( 
.A(n_4399),
.B(n_4118),
.Y(n_4474)
);

AND2x4_ASAP7_75t_L g4475 ( 
.A(n_4326),
.B(n_3825),
.Y(n_4475)
);

AO32x2_ASAP7_75t_L g4476 ( 
.A1(n_4390),
.A2(n_4256),
.A3(n_3795),
.B1(n_3975),
.B2(n_3959),
.Y(n_4476)
);

OAI21x1_ASAP7_75t_SL g4477 ( 
.A1(n_4371),
.A2(n_3909),
.B(n_3907),
.Y(n_4477)
);

AND2x4_ASAP7_75t_L g4478 ( 
.A(n_4326),
.B(n_3826),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_4405),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4408),
.Y(n_4480)
);

AOI22xp33_ASAP7_75t_L g4481 ( 
.A1(n_4446),
.A2(n_4395),
.B1(n_4350),
.B2(n_4368),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4465),
.B(n_4330),
.Y(n_4482)
);

AOI22xp33_ASAP7_75t_SL g4483 ( 
.A1(n_4445),
.A2(n_4381),
.B1(n_4394),
.B2(n_4368),
.Y(n_4483)
);

OR2x2_ASAP7_75t_L g4484 ( 
.A(n_4432),
.B(n_4339),
.Y(n_4484)
);

INVx3_ASAP7_75t_L g4485 ( 
.A(n_4400),
.Y(n_4485)
);

AND2x2_ASAP7_75t_L g4486 ( 
.A(n_4404),
.B(n_4284),
.Y(n_4486)
);

AND2x4_ASAP7_75t_SL g4487 ( 
.A(n_4411),
.B(n_4386),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_4453),
.B(n_4318),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4429),
.B(n_4288),
.Y(n_4489)
);

INVx1_ASAP7_75t_SL g4490 ( 
.A(n_4434),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4456),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4415),
.B(n_4290),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4413),
.B(n_4292),
.Y(n_4493)
);

OR2x2_ASAP7_75t_L g4494 ( 
.A(n_4410),
.B(n_4295),
.Y(n_4494)
);

OAI21xp33_ASAP7_75t_L g4495 ( 
.A1(n_4417),
.A2(n_4358),
.B(n_4297),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4460),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4466),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4471),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4441),
.B(n_4304),
.Y(n_4499)
);

INVx2_ASAP7_75t_SL g4500 ( 
.A(n_4444),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4467),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_4458),
.B(n_4310),
.Y(n_4502)
);

OR2x2_ASAP7_75t_L g4503 ( 
.A(n_4441),
.B(n_4285),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_4442),
.B(n_4452),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4425),
.Y(n_4505)
);

INVx2_ASAP7_75t_L g4506 ( 
.A(n_4425),
.Y(n_4506)
);

NOR2x1_ASAP7_75t_L g4507 ( 
.A(n_4419),
.B(n_4348),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4468),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4459),
.B(n_4393),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4416),
.B(n_4367),
.Y(n_4510)
);

INVx2_ASAP7_75t_SL g4511 ( 
.A(n_4463),
.Y(n_4511)
);

AND2x2_ASAP7_75t_L g4512 ( 
.A(n_4427),
.B(n_4372),
.Y(n_4512)
);

AOI22xp33_ASAP7_75t_L g4513 ( 
.A1(n_4409),
.A2(n_4350),
.B1(n_4316),
.B2(n_4244),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4462),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4439),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4407),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4454),
.B(n_4311),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4424),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4438),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4464),
.B(n_4312),
.Y(n_4520)
);

INVx1_ASAP7_75t_SL g4521 ( 
.A(n_4402),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4440),
.B(n_4320),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4418),
.Y(n_4523)
);

INVx2_ASAP7_75t_SL g4524 ( 
.A(n_4435),
.Y(n_4524)
);

BUFx2_ASAP7_75t_L g4525 ( 
.A(n_4412),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4433),
.B(n_4436),
.Y(n_4526)
);

AND2x4_ASAP7_75t_SL g4527 ( 
.A(n_4437),
.B(n_4396),
.Y(n_4527)
);

BUFx2_ASAP7_75t_L g4528 ( 
.A(n_4414),
.Y(n_4528)
);

AND2x2_ASAP7_75t_L g4529 ( 
.A(n_4420),
.B(n_4366),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4476),
.Y(n_4530)
);

OAI22xp5_ASAP7_75t_L g4531 ( 
.A1(n_4450),
.A2(n_4281),
.B1(n_4303),
.B2(n_4301),
.Y(n_4531)
);

NOR2x1_ASAP7_75t_L g4532 ( 
.A(n_4431),
.B(n_4469),
.Y(n_4532)
);

INVxp67_ASAP7_75t_SL g4533 ( 
.A(n_4447),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4476),
.Y(n_4534)
);

INVx2_ASAP7_75t_SL g4535 ( 
.A(n_4457),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4451),
.Y(n_4536)
);

BUFx2_ASAP7_75t_L g4537 ( 
.A(n_4403),
.Y(n_4537)
);

AND2x2_ASAP7_75t_L g4538 ( 
.A(n_4403),
.B(n_4316),
.Y(n_4538)
);

OR2x2_ASAP7_75t_L g4539 ( 
.A(n_4475),
.B(n_4313),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4455),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4426),
.B(n_4348),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4478),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4430),
.B(n_4360),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4474),
.B(n_4360),
.Y(n_4544)
);

OAI221xp5_ASAP7_75t_SL g4545 ( 
.A1(n_4472),
.A2(n_4240),
.B1(n_4239),
.B2(n_4260),
.C(n_4246),
.Y(n_4545)
);

OAI21xp5_ASAP7_75t_L g4546 ( 
.A1(n_4532),
.A2(n_4443),
.B(n_4421),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4499),
.Y(n_4547)
);

OAI22xp33_ASAP7_75t_SL g4548 ( 
.A1(n_4532),
.A2(n_4449),
.B1(n_4422),
.B2(n_4423),
.Y(n_4548)
);

INVx2_ASAP7_75t_SL g4549 ( 
.A(n_4487),
.Y(n_4549)
);

INVx2_ASAP7_75t_SL g4550 ( 
.A(n_4527),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4522),
.B(n_4281),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4485),
.B(n_4302),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4499),
.Y(n_4553)
);

INVx3_ASAP7_75t_SL g4554 ( 
.A(n_4490),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4485),
.B(n_4302),
.Y(n_4555)
);

AOI21xp5_ASAP7_75t_SL g4556 ( 
.A1(n_4533),
.A2(n_4406),
.B(n_4531),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4496),
.Y(n_4557)
);

INVx1_ASAP7_75t_SL g4558 ( 
.A(n_4490),
.Y(n_4558)
);

NAND2x1_ASAP7_75t_L g4559 ( 
.A(n_4507),
.B(n_4473),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4498),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4491),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4538),
.B(n_4473),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4497),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4522),
.B(n_4331),
.Y(n_4564)
);

OAI22xp33_ASAP7_75t_L g4565 ( 
.A1(n_4521),
.A2(n_4275),
.B1(n_4334),
.B2(n_4448),
.Y(n_4565)
);

INVx3_ASAP7_75t_L g4566 ( 
.A(n_4524),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4493),
.Y(n_4567)
);

OR2x2_ASAP7_75t_L g4568 ( 
.A(n_4484),
.B(n_4488),
.Y(n_4568)
);

AND2x4_ASAP7_75t_L g4569 ( 
.A(n_4523),
.B(n_4299),
.Y(n_4569)
);

CKINVDCx20_ASAP7_75t_R g4570 ( 
.A(n_4535),
.Y(n_4570)
);

OAI33xp33_ASAP7_75t_L g4571 ( 
.A1(n_4536),
.A2(n_4470),
.A3(n_3834),
.B1(n_3835),
.B2(n_3820),
.B3(n_4401),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4479),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4494),
.Y(n_4573)
);

BUFx3_ASAP7_75t_L g4574 ( 
.A(n_4500),
.Y(n_4574)
);

AND2x4_ASAP7_75t_L g4575 ( 
.A(n_4507),
.B(n_4271),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4526),
.B(n_4337),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4482),
.Y(n_4577)
);

BUFx4f_ASAP7_75t_L g4578 ( 
.A(n_4511),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_4503),
.Y(n_4579)
);

OR2x2_ASAP7_75t_L g4580 ( 
.A(n_4492),
.B(n_4355),
.Y(n_4580)
);

INVx4_ASAP7_75t_L g4581 ( 
.A(n_4525),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4489),
.Y(n_4582)
);

NOR2xp67_ASAP7_75t_L g4583 ( 
.A(n_4530),
.B(n_673),
.Y(n_4583)
);

HB1xp67_ASAP7_75t_L g4584 ( 
.A(n_4521),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4520),
.B(n_4461),
.Y(n_4585)
);

AOI221xp5_ASAP7_75t_L g4586 ( 
.A1(n_4495),
.A2(n_4428),
.B1(n_4477),
.B2(n_3924),
.C(n_4038),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4515),
.B(n_4357),
.Y(n_4587)
);

AOI221xp5_ASAP7_75t_L g4588 ( 
.A1(n_4495),
.A2(n_4428),
.B1(n_4477),
.B2(n_4060),
.C(n_4057),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4480),
.Y(n_4589)
);

AOI322xp5_ASAP7_75t_L g4590 ( 
.A1(n_4534),
.A2(n_4481),
.A3(n_4513),
.B1(n_4541),
.B2(n_4504),
.C1(n_4517),
.C2(n_4510),
.Y(n_4590)
);

AOI22xp33_ASAP7_75t_L g4591 ( 
.A1(n_4501),
.A2(n_4294),
.B1(n_4384),
.B2(n_4210),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4519),
.B(n_4364),
.Y(n_4592)
);

OAI33xp33_ASAP7_75t_L g4593 ( 
.A1(n_4531),
.A2(n_3459),
.A3(n_3505),
.B1(n_3465),
.B2(n_4354),
.B3(n_4345),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4502),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4486),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4537),
.B(n_4343),
.Y(n_4596)
);

OR2x2_ASAP7_75t_L g4597 ( 
.A(n_4505),
.B(n_4349),
.Y(n_4597)
);

BUFx6f_ASAP7_75t_L g4598 ( 
.A(n_4528),
.Y(n_4598)
);

AND2x2_ASAP7_75t_L g4599 ( 
.A(n_4512),
.B(n_4306),
.Y(n_4599)
);

BUFx3_ASAP7_75t_L g4600 ( 
.A(n_4543),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4539),
.Y(n_4601)
);

OR2x2_ASAP7_75t_L g4602 ( 
.A(n_4506),
.B(n_4307),
.Y(n_4602)
);

HB1xp67_ASAP7_75t_L g4603 ( 
.A(n_4516),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4581),
.B(n_4518),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4562),
.B(n_4529),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_L g4606 ( 
.A(n_4590),
.B(n_4540),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4581),
.B(n_4509),
.Y(n_4607)
);

AND3x2_ASAP7_75t_L g4608 ( 
.A(n_4556),
.B(n_4544),
.C(n_4483),
.Y(n_4608)
);

AND2x4_ASAP7_75t_SL g4609 ( 
.A(n_4570),
.B(n_4514),
.Y(n_4609)
);

AND2x2_ASAP7_75t_L g4610 ( 
.A(n_4598),
.B(n_4508),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4598),
.B(n_4542),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4598),
.B(n_4271),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4584),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4547),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4553),
.Y(n_4615)
);

NAND2xp5_ASAP7_75t_L g4616 ( 
.A(n_4567),
.B(n_4561),
.Y(n_4616)
);

OAI22xp5_ASAP7_75t_L g4617 ( 
.A1(n_4554),
.A2(n_4545),
.B1(n_4264),
.B2(n_3927),
.Y(n_4617)
);

INVx3_ASAP7_75t_L g4618 ( 
.A(n_4575),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4563),
.B(n_3886),
.Y(n_4619)
);

NAND2x1p5_ASAP7_75t_L g4620 ( 
.A(n_4578),
.B(n_3226),
.Y(n_4620)
);

NOR2x1_ASAP7_75t_L g4621 ( 
.A(n_4546),
.B(n_3995),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4552),
.B(n_4375),
.Y(n_4622)
);

INVxp67_ASAP7_75t_SL g4623 ( 
.A(n_4583),
.Y(n_4623)
);

AOI22xp33_ASAP7_75t_L g4624 ( 
.A1(n_4571),
.A2(n_4024),
.B1(n_3797),
.B2(n_4076),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4580),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4555),
.B(n_3795),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4603),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4599),
.B(n_4558),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4557),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4566),
.B(n_3959),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4560),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4564),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4585),
.B(n_3975),
.Y(n_4633)
);

NAND2xp5_ASAP7_75t_L g4634 ( 
.A(n_4577),
.B(n_4573),
.Y(n_4634)
);

OR2x2_ASAP7_75t_L g4635 ( 
.A(n_4568),
.B(n_3918),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4572),
.Y(n_4636)
);

INVxp67_ASAP7_75t_L g4637 ( 
.A(n_4623),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4604),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4616),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4616),
.Y(n_4640)
);

OR2x2_ASAP7_75t_L g4641 ( 
.A(n_4635),
.B(n_4551),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4606),
.B(n_4591),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4606),
.B(n_4582),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4634),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4634),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4625),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4632),
.Y(n_4647)
);

AND2x2_ASAP7_75t_L g4648 ( 
.A(n_4628),
.B(n_4549),
.Y(n_4648)
);

INVxp67_ASAP7_75t_SL g4649 ( 
.A(n_4621),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4629),
.Y(n_4650)
);

INVxp33_ASAP7_75t_L g4651 ( 
.A(n_4620),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_SL g4652 ( 
.A(n_4618),
.B(n_4548),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4605),
.B(n_4569),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4631),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4613),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4627),
.B(n_4588),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4614),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_4615),
.B(n_4619),
.Y(n_4658)
);

NOR2xp33_ASAP7_75t_L g4659 ( 
.A(n_4609),
.B(n_4550),
.Y(n_4659)
);

INVx2_ASAP7_75t_L g4660 ( 
.A(n_4607),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4636),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4630),
.B(n_4595),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4610),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4619),
.Y(n_4664)
);

AND2x2_ASAP7_75t_L g4665 ( 
.A(n_4611),
.B(n_4569),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4633),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4626),
.B(n_4594),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4618),
.Y(n_4668)
);

INVx1_ASAP7_75t_SL g4669 ( 
.A(n_4612),
.Y(n_4669)
);

OR2x2_ASAP7_75t_L g4670 ( 
.A(n_4622),
.B(n_4579),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4608),
.B(n_4574),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4617),
.B(n_4600),
.Y(n_4672)
);

INVx3_ASAP7_75t_L g4673 ( 
.A(n_4617),
.Y(n_4673)
);

OR2x2_ASAP7_75t_L g4674 ( 
.A(n_4624),
.B(n_4601),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4616),
.Y(n_4675)
);

AND2x4_ASAP7_75t_SL g4676 ( 
.A(n_4607),
.B(n_4576),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4616),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4614),
.B(n_4589),
.Y(n_4678)
);

OR2x2_ASAP7_75t_L g4679 ( 
.A(n_4635),
.B(n_4597),
.Y(n_4679)
);

OAI22xp33_ASAP7_75t_L g4680 ( 
.A1(n_4642),
.A2(n_4559),
.B1(n_4565),
.B2(n_4575),
.Y(n_4680)
);

AOI21xp33_ASAP7_75t_L g4681 ( 
.A1(n_4637),
.A2(n_4559),
.B(n_4602),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4678),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4639),
.B(n_4592),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4671),
.B(n_4672),
.Y(n_4684)
);

AND2x2_ASAP7_75t_L g4685 ( 
.A(n_4648),
.B(n_4665),
.Y(n_4685)
);

NOR2x1_ASAP7_75t_L g4686 ( 
.A(n_4652),
.B(n_3896),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4653),
.B(n_4596),
.Y(n_4687)
);

NAND4xp25_ASAP7_75t_SL g4688 ( 
.A(n_4643),
.B(n_4586),
.C(n_4587),
.D(n_4593),
.Y(n_4688)
);

AND2x2_ASAP7_75t_L g4689 ( 
.A(n_4660),
.B(n_3918),
.Y(n_4689)
);

AND2x2_ASAP7_75t_L g4690 ( 
.A(n_4659),
.B(n_3803),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4673),
.B(n_3824),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4673),
.B(n_3824),
.Y(n_4692)
);

NAND2xp33_ASAP7_75t_SL g4693 ( 
.A(n_4651),
.B(n_3226),
.Y(n_4693)
);

AOI21xp33_ASAP7_75t_L g4694 ( 
.A1(n_4649),
.A2(n_675),
.B(n_676),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4644),
.B(n_3979),
.Y(n_4695)
);

INVx2_ASAP7_75t_L g4696 ( 
.A(n_4638),
.Y(n_4696)
);

OR2x2_ASAP7_75t_L g4697 ( 
.A(n_4674),
.B(n_3979),
.Y(n_4697)
);

AND2x2_ASAP7_75t_L g4698 ( 
.A(n_4663),
.B(n_3803),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4678),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4645),
.B(n_4003),
.Y(n_4700)
);

INVx2_ASAP7_75t_L g4701 ( 
.A(n_4676),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4669),
.B(n_3803),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4640),
.B(n_3810),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4675),
.B(n_3785),
.Y(n_4704)
);

BUFx3_ASAP7_75t_L g4705 ( 
.A(n_4668),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4677),
.B(n_3969),
.Y(n_4706)
);

AOI21xp5_ASAP7_75t_L g4707 ( 
.A1(n_4656),
.A2(n_4026),
.B(n_3998),
.Y(n_4707)
);

NOR2xp67_ASAP7_75t_L g4708 ( 
.A(n_4664),
.B(n_676),
.Y(n_4708)
);

OR2x2_ASAP7_75t_L g4709 ( 
.A(n_4666),
.B(n_3796),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4647),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4646),
.B(n_4030),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4657),
.B(n_4033),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4650),
.B(n_4046),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4655),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4654),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4661),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4658),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4669),
.B(n_3796),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4641),
.B(n_3811),
.Y(n_4719)
);

OR2x2_ASAP7_75t_L g4720 ( 
.A(n_4667),
.B(n_677),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4696),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4706),
.Y(n_4722)
);

O2A1O1Ixp5_ASAP7_75t_L g4723 ( 
.A1(n_4680),
.A2(n_4684),
.B(n_4681),
.C(n_4701),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4682),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4699),
.Y(n_4725)
);

AOI322xp5_ASAP7_75t_L g4726 ( 
.A1(n_4686),
.A2(n_4658),
.A3(n_4662),
.B1(n_4679),
.B2(n_4670),
.C1(n_3366),
.C2(n_3365),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4690),
.B(n_677),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4705),
.Y(n_4728)
);

O2A1O1Ixp5_ASAP7_75t_L g4729 ( 
.A1(n_4681),
.A2(n_3402),
.B(n_3392),
.C(n_3337),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4700),
.Y(n_4730)
);

OAI21xp33_ASAP7_75t_L g4731 ( 
.A1(n_4688),
.A2(n_4047),
.B(n_3357),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4710),
.Y(n_4732)
);

INVx1_ASAP7_75t_SL g4733 ( 
.A(n_4720),
.Y(n_4733)
);

AOI32xp33_ASAP7_75t_L g4734 ( 
.A1(n_4693),
.A2(n_3432),
.A3(n_3476),
.B1(n_3415),
.B2(n_3322),
.Y(n_4734)
);

HB1xp67_ASAP7_75t_L g4735 ( 
.A(n_4714),
.Y(n_4735)
);

NOR2xp33_ASAP7_75t_L g4736 ( 
.A(n_4685),
.B(n_678),
.Y(n_4736)
);

INVx1_ASAP7_75t_SL g4737 ( 
.A(n_4704),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4716),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_SL g4739 ( 
.A(n_4708),
.B(n_3226),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4715),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4717),
.B(n_678),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4711),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4687),
.B(n_679),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4712),
.Y(n_4744)
);

OAI22xp5_ASAP7_75t_L g4745 ( 
.A1(n_4697),
.A2(n_3728),
.B1(n_3266),
.B2(n_3325),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4713),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4708),
.B(n_679),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4703),
.B(n_680),
.Y(n_4748)
);

NOR2xp33_ASAP7_75t_L g4749 ( 
.A(n_4683),
.B(n_681),
.Y(n_4749)
);

OR2x2_ASAP7_75t_L g4750 ( 
.A(n_4691),
.B(n_4692),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4707),
.B(n_681),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4689),
.Y(n_4752)
);

OAI221xp5_ASAP7_75t_L g4753 ( 
.A1(n_4694),
.A2(n_3839),
.B1(n_3728),
.B2(n_3515),
.C(n_3523),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4683),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4728),
.B(n_4698),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4737),
.B(n_4719),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4733),
.B(n_4722),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4754),
.B(n_4695),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4721),
.Y(n_4759)
);

INVxp67_ASAP7_75t_L g4760 ( 
.A(n_4749),
.Y(n_4760)
);

NAND3xp33_ASAP7_75t_SL g4761 ( 
.A(n_4723),
.B(n_4702),
.C(n_4718),
.Y(n_4761)
);

INVx2_ASAP7_75t_L g4762 ( 
.A(n_4735),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4730),
.B(n_4751),
.Y(n_4763)
);

AO21x1_ASAP7_75t_L g4764 ( 
.A1(n_4732),
.A2(n_4694),
.B(n_4709),
.Y(n_4764)
);

BUFx2_ASAP7_75t_L g4765 ( 
.A(n_4724),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4743),
.Y(n_4766)
);

OAI22xp33_ASAP7_75t_L g4767 ( 
.A1(n_4727),
.A2(n_3266),
.B1(n_3325),
.B2(n_3260),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4747),
.Y(n_4768)
);

OAI211xp5_ASAP7_75t_SL g4769 ( 
.A1(n_4731),
.A2(n_684),
.B(n_682),
.C(n_683),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4725),
.B(n_683),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4752),
.B(n_684),
.Y(n_4771)
);

NOR2xp33_ASAP7_75t_SL g4772 ( 
.A(n_4736),
.B(n_3260),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4738),
.Y(n_4773)
);

OAI22xp33_ASAP7_75t_SL g4774 ( 
.A1(n_4740),
.A2(n_3504),
.B1(n_3530),
.B2(n_3481),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4748),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4741),
.Y(n_4776)
);

OAI22xp5_ASAP7_75t_L g4777 ( 
.A1(n_4750),
.A2(n_3540),
.B1(n_3266),
.B2(n_3325),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4742),
.B(n_685),
.Y(n_4778)
);

INVxp67_ASAP7_75t_L g4779 ( 
.A(n_4739),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_L g4780 ( 
.A(n_4744),
.B(n_685),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4746),
.Y(n_4781)
);

AOI22xp5_ASAP7_75t_L g4782 ( 
.A1(n_4753),
.A2(n_3381),
.B1(n_3426),
.B2(n_3260),
.Y(n_4782)
);

OAI221xp5_ASAP7_75t_L g4783 ( 
.A1(n_4729),
.A2(n_688),
.B1(n_686),
.B2(n_687),
.C(n_689),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4745),
.Y(n_4784)
);

CKINVDCx14_ASAP7_75t_R g4785 ( 
.A(n_4757),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4762),
.B(n_4726),
.Y(n_4786)
);

O2A1O1Ixp33_ASAP7_75t_L g4787 ( 
.A1(n_4761),
.A2(n_4726),
.B(n_4734),
.C(n_690),
.Y(n_4787)
);

OAI22xp5_ASAP7_75t_L g4788 ( 
.A1(n_4760),
.A2(n_3426),
.B1(n_3463),
.B2(n_3381),
.Y(n_4788)
);

INVxp67_ASAP7_75t_L g4789 ( 
.A(n_4765),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4755),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4759),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4766),
.B(n_688),
.Y(n_4792)
);

AOI221xp5_ASAP7_75t_L g4793 ( 
.A1(n_4781),
.A2(n_691),
.B1(n_689),
.B2(n_690),
.C(n_692),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_SL g4794 ( 
.A(n_4764),
.B(n_3381),
.Y(n_4794)
);

NOR2xp33_ASAP7_75t_L g4795 ( 
.A(n_4784),
.B(n_693),
.Y(n_4795)
);

OAI221xp5_ASAP7_75t_SL g4796 ( 
.A1(n_4779),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.C(n_696),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4771),
.Y(n_4797)
);

INVxp33_ASAP7_75t_SL g4798 ( 
.A(n_4770),
.Y(n_4798)
);

AND2x2_ASAP7_75t_L g4799 ( 
.A(n_4756),
.B(n_694),
.Y(n_4799)
);

INVx8_ASAP7_75t_L g4800 ( 
.A(n_4778),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4780),
.Y(n_4801)
);

XNOR2x1_ASAP7_75t_L g4802 ( 
.A(n_4768),
.B(n_4775),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4776),
.B(n_695),
.Y(n_4803)
);

INVx1_ASAP7_75t_SL g4804 ( 
.A(n_4763),
.Y(n_4804)
);

INVxp67_ASAP7_75t_SL g4805 ( 
.A(n_4773),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4774),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4774),
.Y(n_4807)
);

AOI22xp5_ASAP7_75t_L g4808 ( 
.A1(n_4772),
.A2(n_3463),
.B1(n_3538),
.B2(n_3426),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4758),
.Y(n_4809)
);

INVx1_ASAP7_75t_SL g4810 ( 
.A(n_4777),
.Y(n_4810)
);

NOR2xp33_ASAP7_75t_L g4811 ( 
.A(n_4783),
.B(n_696),
.Y(n_4811)
);

NOR2xp33_ASAP7_75t_L g4812 ( 
.A(n_4769),
.B(n_697),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_4767),
.B(n_697),
.Y(n_4813)
);

AOI21xp5_ASAP7_75t_L g4814 ( 
.A1(n_4782),
.A2(n_699),
.B(n_700),
.Y(n_4814)
);

OAI21xp33_ASAP7_75t_SL g4815 ( 
.A1(n_4782),
.A2(n_701),
.B(n_702),
.Y(n_4815)
);

OA22x2_ASAP7_75t_L g4816 ( 
.A1(n_4762),
.A2(n_705),
.B1(n_703),
.B2(n_704),
.Y(n_4816)
);

XNOR2xp5_ASAP7_75t_L g4817 ( 
.A(n_4771),
.B(n_703),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4755),
.B(n_704),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4816),
.Y(n_4819)
);

NAND3xp33_ASAP7_75t_L g4820 ( 
.A(n_4785),
.B(n_3538),
.C(n_3463),
.Y(n_4820)
);

INVx1_ASAP7_75t_L g4821 ( 
.A(n_4790),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4818),
.B(n_706),
.Y(n_4822)
);

NAND3xp33_ASAP7_75t_L g4823 ( 
.A(n_4795),
.B(n_3578),
.C(n_3538),
.Y(n_4823)
);

AOI21xp33_ASAP7_75t_L g4824 ( 
.A1(n_4789),
.A2(n_706),
.B(n_707),
.Y(n_4824)
);

NOR2x1_ASAP7_75t_L g4825 ( 
.A(n_4803),
.B(n_707),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4799),
.B(n_708),
.Y(n_4826)
);

AOI221xp5_ASAP7_75t_L g4827 ( 
.A1(n_4787),
.A2(n_711),
.B1(n_709),
.B2(n_710),
.C(n_712),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4812),
.B(n_4817),
.Y(n_4828)
);

OAI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4815),
.A2(n_711),
.B(n_712),
.Y(n_4829)
);

AOI21xp5_ASAP7_75t_L g4830 ( 
.A1(n_4794),
.A2(n_713),
.B(n_714),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4805),
.Y(n_4831)
);

INVx1_ASAP7_75t_SL g4832 ( 
.A(n_4810),
.Y(n_4832)
);

NOR3x1_ASAP7_75t_L g4833 ( 
.A(n_4786),
.B(n_713),
.C(n_714),
.Y(n_4833)
);

AOI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4792),
.A2(n_715),
.B(n_716),
.Y(n_4834)
);

NOR3xp33_ASAP7_75t_L g4835 ( 
.A(n_4796),
.B(n_4813),
.C(n_4793),
.Y(n_4835)
);

HB1xp67_ASAP7_75t_L g4836 ( 
.A(n_4791),
.Y(n_4836)
);

O2A1O1Ixp5_ASAP7_75t_L g4837 ( 
.A1(n_4809),
.A2(n_717),
.B(n_715),
.C(n_716),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_L g4838 ( 
.A(n_4811),
.B(n_717),
.Y(n_4838)
);

NOR2xp33_ASAP7_75t_L g4839 ( 
.A(n_4798),
.B(n_718),
.Y(n_4839)
);

OR2x2_ASAP7_75t_L g4840 ( 
.A(n_4804),
.B(n_718),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4797),
.Y(n_4841)
);

INVx2_ASAP7_75t_L g4842 ( 
.A(n_4800),
.Y(n_4842)
);

O2A1O1Ixp33_ASAP7_75t_SL g4843 ( 
.A1(n_4806),
.A2(n_722),
.B(n_719),
.C(n_720),
.Y(n_4843)
);

NAND3xp33_ASAP7_75t_L g4844 ( 
.A(n_4814),
.B(n_3581),
.C(n_3578),
.Y(n_4844)
);

NOR2x1_ASAP7_75t_SL g4845 ( 
.A(n_4801),
.B(n_3578),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4807),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4802),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4800),
.Y(n_4848)
);

NAND3xp33_ASAP7_75t_L g4849 ( 
.A(n_4788),
.B(n_3584),
.C(n_3581),
.Y(n_4849)
);

OAI21xp5_ASAP7_75t_L g4850 ( 
.A1(n_4830),
.A2(n_4808),
.B(n_719),
.Y(n_4850)
);

AOI221xp5_ASAP7_75t_L g4851 ( 
.A1(n_4843),
.A2(n_724),
.B1(n_722),
.B2(n_723),
.C(n_725),
.Y(n_4851)
);

AOI21xp33_ASAP7_75t_L g4852 ( 
.A1(n_4832),
.A2(n_724),
.B(n_725),
.Y(n_4852)
);

AOI22xp5_ASAP7_75t_L g4853 ( 
.A1(n_4827),
.A2(n_4819),
.B1(n_4835),
.B2(n_4839),
.Y(n_4853)
);

AOI221xp5_ASAP7_75t_L g4854 ( 
.A1(n_4831),
.A2(n_4848),
.B1(n_4846),
.B2(n_4836),
.C(n_4847),
.Y(n_4854)
);

OAI221xp5_ASAP7_75t_L g4855 ( 
.A1(n_4829),
.A2(n_729),
.B1(n_727),
.B2(n_728),
.C(n_730),
.Y(n_4855)
);

INVx2_ASAP7_75t_SL g4856 ( 
.A(n_4842),
.Y(n_4856)
);

A2O1A1Ixp33_ASAP7_75t_L g4857 ( 
.A1(n_4837),
.A2(n_730),
.B(n_727),
.C(n_729),
.Y(n_4857)
);

AOI221xp5_ASAP7_75t_L g4858 ( 
.A1(n_4821),
.A2(n_734),
.B1(n_731),
.B2(n_733),
.C(n_735),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4840),
.Y(n_4859)
);

AOI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_4838),
.A2(n_3584),
.B1(n_3587),
.B2(n_3581),
.Y(n_4860)
);

AOI322xp5_ASAP7_75t_L g4861 ( 
.A1(n_4841),
.A2(n_733),
.A3(n_735),
.B1(n_736),
.B2(n_737),
.C1(n_738),
.C2(n_739),
.Y(n_4861)
);

OR2x2_ASAP7_75t_L g4862 ( 
.A(n_4826),
.B(n_736),
.Y(n_4862)
);

OAI211xp5_ASAP7_75t_SL g4863 ( 
.A1(n_4828),
.A2(n_740),
.B(n_737),
.C(n_739),
.Y(n_4863)
);

OAI21x1_ASAP7_75t_SL g4864 ( 
.A1(n_4845),
.A2(n_4834),
.B(n_4825),
.Y(n_4864)
);

OAI22xp33_ASAP7_75t_L g4865 ( 
.A1(n_4820),
.A2(n_3587),
.B1(n_3640),
.B2(n_3584),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4833),
.B(n_742),
.Y(n_4866)
);

AOI211x1_ASAP7_75t_SL g4867 ( 
.A1(n_4824),
.A2(n_745),
.B(n_743),
.C(n_744),
.Y(n_4867)
);

NAND4xp25_ASAP7_75t_L g4868 ( 
.A(n_4822),
.B(n_747),
.C(n_744),
.D(n_746),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4844),
.B(n_748),
.Y(n_4869)
);

NAND4xp75_ASAP7_75t_L g4870 ( 
.A(n_4823),
.B(n_753),
.C(n_751),
.D(n_752),
.Y(n_4870)
);

AOI211xp5_ASAP7_75t_L g4871 ( 
.A1(n_4849),
.A2(n_755),
.B(n_752),
.C(n_754),
.Y(n_4871)
);

AOI321xp33_ASAP7_75t_L g4872 ( 
.A1(n_4831),
.A2(n_756),
.A3(n_758),
.B1(n_754),
.B2(n_755),
.C(n_757),
.Y(n_4872)
);

OAI211xp5_ASAP7_75t_L g4873 ( 
.A1(n_4854),
.A2(n_758),
.B(n_756),
.C(n_757),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4856),
.Y(n_4874)
);

HB1xp67_ASAP7_75t_L g4875 ( 
.A(n_4869),
.Y(n_4875)
);

AOI211xp5_ASAP7_75t_L g4876 ( 
.A1(n_4852),
.A2(n_761),
.B(n_759),
.C(n_760),
.Y(n_4876)
);

AOI221xp5_ASAP7_75t_L g4877 ( 
.A1(n_4855),
.A2(n_3662),
.B1(n_3663),
.B2(n_3640),
.C(n_3587),
.Y(n_4877)
);

OAI21xp33_ASAP7_75t_L g4878 ( 
.A1(n_4853),
.A2(n_4859),
.B(n_4850),
.Y(n_4878)
);

NAND3xp33_ASAP7_75t_L g4879 ( 
.A(n_4858),
.B(n_759),
.C(n_760),
.Y(n_4879)
);

OR2x2_ASAP7_75t_L g4880 ( 
.A(n_4866),
.B(n_762),
.Y(n_4880)
);

O2A1O1Ixp33_ASAP7_75t_L g4881 ( 
.A1(n_4857),
.A2(n_764),
.B(n_762),
.C(n_763),
.Y(n_4881)
);

BUFx6f_ASAP7_75t_L g4882 ( 
.A(n_4862),
.Y(n_4882)
);

NAND4xp25_ASAP7_75t_SL g4883 ( 
.A(n_4851),
.B(n_766),
.C(n_764),
.D(n_765),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4870),
.Y(n_4884)
);

NAND4xp75_ASAP7_75t_L g4885 ( 
.A(n_4867),
.B(n_768),
.C(n_765),
.D(n_766),
.Y(n_4885)
);

NOR3xp33_ASAP7_75t_L g4886 ( 
.A(n_4863),
.B(n_769),
.C(n_770),
.Y(n_4886)
);

AOI211x1_ASAP7_75t_L g4887 ( 
.A1(n_4868),
.A2(n_772),
.B(n_769),
.C(n_771),
.Y(n_4887)
);

AOI21xp5_ASAP7_75t_L g4888 ( 
.A1(n_4864),
.A2(n_772),
.B(n_773),
.Y(n_4888)
);

AOI221xp5_ASAP7_75t_L g4889 ( 
.A1(n_4871),
.A2(n_3679),
.B1(n_3696),
.B2(n_3663),
.C(n_3662),
.Y(n_4889)
);

AOI22xp33_ASAP7_75t_L g4890 ( 
.A1(n_4865),
.A2(n_3663),
.B1(n_3679),
.B2(n_3662),
.Y(n_4890)
);

AOI221x1_ASAP7_75t_L g4891 ( 
.A1(n_4861),
.A2(n_775),
.B1(n_773),
.B2(n_774),
.C(n_776),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4860),
.B(n_774),
.Y(n_4892)
);

NOR2x1_ASAP7_75t_L g4893 ( 
.A(n_4872),
.B(n_776),
.Y(n_4893)
);

OAI21xp33_ASAP7_75t_L g4894 ( 
.A1(n_4856),
.A2(n_777),
.B(n_778),
.Y(n_4894)
);

NAND2x1p5_ASAP7_75t_L g4895 ( 
.A(n_4874),
.B(n_3679),
.Y(n_4895)
);

NOR2x1_ASAP7_75t_L g4896 ( 
.A(n_4873),
.B(n_4888),
.Y(n_4896)
);

OAI21xp5_ASAP7_75t_L g4897 ( 
.A1(n_4893),
.A2(n_777),
.B(n_779),
.Y(n_4897)
);

HB1xp67_ASAP7_75t_L g4898 ( 
.A(n_4884),
.Y(n_4898)
);

XNOR2xp5_ASAP7_75t_L g4899 ( 
.A(n_4887),
.B(n_780),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4894),
.Y(n_4900)
);

AND2x2_ASAP7_75t_L g4901 ( 
.A(n_4882),
.B(n_781),
.Y(n_4901)
);

INVx2_ASAP7_75t_L g4902 ( 
.A(n_4882),
.Y(n_4902)
);

OR2x2_ASAP7_75t_L g4903 ( 
.A(n_4880),
.B(n_781),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4882),
.B(n_782),
.Y(n_4904)
);

NOR2x1_ASAP7_75t_L g4905 ( 
.A(n_4879),
.B(n_782),
.Y(n_4905)
);

OR2x2_ASAP7_75t_L g4906 ( 
.A(n_4892),
.B(n_783),
.Y(n_4906)
);

NAND4xp75_ASAP7_75t_L g4907 ( 
.A(n_4891),
.B(n_786),
.C(n_783),
.D(n_784),
.Y(n_4907)
);

NOR2x1p5_ASAP7_75t_L g4908 ( 
.A(n_4885),
.B(n_4883),
.Y(n_4908)
);

NOR2x1_ASAP7_75t_L g4909 ( 
.A(n_4878),
.B(n_786),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4881),
.Y(n_4910)
);

NOR3xp33_ASAP7_75t_L g4911 ( 
.A(n_4902),
.B(n_4876),
.C(n_4886),
.Y(n_4911)
);

NOR3x1_ASAP7_75t_L g4912 ( 
.A(n_4907),
.B(n_4875),
.C(n_4877),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4901),
.B(n_4890),
.Y(n_4913)
);

NAND4xp75_ASAP7_75t_L g4914 ( 
.A(n_4909),
.B(n_4889),
.C(n_789),
.D(n_787),
.Y(n_4914)
);

AOI322xp5_ASAP7_75t_L g4915 ( 
.A1(n_4898),
.A2(n_3737),
.A3(n_3735),
.B1(n_3696),
.B2(n_790),
.C1(n_791),
.C2(n_792),
.Y(n_4915)
);

OAI211xp5_ASAP7_75t_SL g4916 ( 
.A1(n_4896),
.A2(n_789),
.B(n_787),
.C(n_788),
.Y(n_4916)
);

AND2x4_ASAP7_75t_L g4917 ( 
.A(n_4904),
.B(n_788),
.Y(n_4917)
);

NOR2xp67_ASAP7_75t_L g4918 ( 
.A(n_4900),
.B(n_790),
.Y(n_4918)
);

NOR3xp33_ASAP7_75t_L g4919 ( 
.A(n_4897),
.B(n_791),
.C(n_793),
.Y(n_4919)
);

OAI211xp5_ASAP7_75t_SL g4920 ( 
.A1(n_4910),
.A2(n_795),
.B(n_793),
.C(n_794),
.Y(n_4920)
);

OAI21xp5_ASAP7_75t_L g4921 ( 
.A1(n_4899),
.A2(n_795),
.B(n_796),
.Y(n_4921)
);

XOR2xp5_ASAP7_75t_L g4922 ( 
.A(n_4914),
.B(n_4903),
.Y(n_4922)
);

AOI211xp5_ASAP7_75t_L g4923 ( 
.A1(n_4920),
.A2(n_4906),
.B(n_4908),
.C(n_4905),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_4917),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4918),
.B(n_4895),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4917),
.B(n_4915),
.Y(n_4926)
);

OAI22xp5_ASAP7_75t_L g4927 ( 
.A1(n_4921),
.A2(n_3735),
.B1(n_3737),
.B2(n_3696),
.Y(n_4927)
);

AO22x2_ASAP7_75t_L g4928 ( 
.A1(n_4922),
.A2(n_4911),
.B1(n_4913),
.B2(n_4919),
.Y(n_4928)
);

AOI22x1_ASAP7_75t_SL g4929 ( 
.A1(n_4924),
.A2(n_4912),
.B1(n_4916),
.B2(n_799),
.Y(n_4929)
);

OAI22xp5_ASAP7_75t_SL g4930 ( 
.A1(n_4926),
.A2(n_799),
.B1(n_796),
.B2(n_797),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4925),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4931),
.Y(n_4932)
);

NOR2xp33_ASAP7_75t_L g4933 ( 
.A(n_4930),
.B(n_4927),
.Y(n_4933)
);

OR2x6_ASAP7_75t_L g4934 ( 
.A(n_4928),
.B(n_4923),
.Y(n_4934)
);

AO22x2_ASAP7_75t_L g4935 ( 
.A1(n_4932),
.A2(n_4929),
.B1(n_4934),
.B2(n_4933),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4932),
.Y(n_4936)
);

OAI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4936),
.A2(n_3737),
.B1(n_3735),
.B2(n_801),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4935),
.A2(n_797),
.B(n_800),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_SL g4939 ( 
.A(n_4936),
.B(n_802),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4939),
.Y(n_4940)
);

OAI21xp5_ASAP7_75t_L g4941 ( 
.A1(n_4938),
.A2(n_802),
.B(n_803),
.Y(n_4941)
);

AOI21xp33_ASAP7_75t_SL g4942 ( 
.A1(n_4937),
.A2(n_803),
.B(n_804),
.Y(n_4942)
);

OAI21x1_ASAP7_75t_SL g4943 ( 
.A1(n_4940),
.A2(n_806),
.B(n_807),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4941),
.B(n_807),
.Y(n_4944)
);

AOI22xp33_ASAP7_75t_L g4945 ( 
.A1(n_4942),
.A2(n_810),
.B1(n_808),
.B2(n_809),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_L g4946 ( 
.A(n_4945),
.B(n_808),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4943),
.Y(n_4947)
);

AOI221xp5_ASAP7_75t_L g4948 ( 
.A1(n_4947),
.A2(n_4944),
.B1(n_812),
.B2(n_809),
.C(n_811),
.Y(n_4948)
);

AOI211xp5_ASAP7_75t_L g4949 ( 
.A1(n_4948),
.A2(n_4946),
.B(n_814),
.C(n_812),
.Y(n_4949)
);


endmodule