module real_jpeg_32511_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_244;
wire n_202;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_0),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_0),
.Y(n_154)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_0),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_0),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_34),
.B1(n_39),
.B2(n_44),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_1),
.A2(n_44),
.B1(n_167),
.B2(n_171),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_2),
.A2(n_102),
.B1(n_107),
.B2(n_108),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_2),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_107),
.B1(n_133),
.B2(n_137),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_107),
.B1(n_187),
.B2(n_191),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_69),
.B1(n_74),
.B2(n_77),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_3),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_3),
.A2(n_176),
.B(n_177),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_5),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_6),
.A2(n_157),
.B1(n_161),
.B2(n_163),
.Y(n_156)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_8),
.A2(n_58),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_196),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_194),
.Y(n_12)
);

INVxp33_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_164),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_15),
.B(n_164),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_113),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_67),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_32),
.B1(n_45),
.B2(n_56),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_20),
.Y(n_184)
);

OAI22x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_22),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_23),
.Y(n_145)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_28),
.Y(n_175)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_29),
.Y(n_136)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_29),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_29),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_31),
.Y(n_225)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_45),
.B(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_46),
.A2(n_57),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

BUFx4f_ASAP7_75t_SL g214 ( 
.A(n_48),
.Y(n_214)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_50),
.Y(n_190)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_55),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_66),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_78),
.B(n_99),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_116),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_126),
.C(n_128),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_R g180 ( 
.A(n_77),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_77),
.B(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_77),
.A2(n_226),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_77),
.B(n_183),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_77),
.B(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

AOI22x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_86),
.B2(n_89),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_130),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_119),
.B(n_125),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_128),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_148),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_131),
.A2(n_245),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_143),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_142),
.Y(n_249)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_143),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_180),
.C(n_182),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_176),
.B(n_177),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_233),
.B(n_273),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_201),
.B(n_206),
.Y(n_274)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_228),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_207),
.A2(n_228),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

AO221x1_ASAP7_75t_L g272 ( 
.A1(n_207),
.A2(n_228),
.B1(n_238),
.B2(n_252),
.C(n_253),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_220),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_224),
.B(n_226),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_254),
.B(n_272),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_251),
.Y(n_237)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_262),
.B(n_271),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_257),
.B(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);


endmodule