module fake_jpeg_18578_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_33),
.B1(n_32),
.B2(n_18),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_23),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_32),
.Y(n_76)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_62),
.B(n_78),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_60),
.B1(n_55),
.B2(n_24),
.Y(n_103)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_92),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_33),
.B1(n_43),
.B2(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_86),
.B1(n_91),
.B2(n_65),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_81),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_35),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_94),
.B1(n_30),
.B2(n_29),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_33),
.B1(n_16),
.B2(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_21),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_44),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_46),
.C(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_21),
.B1(n_27),
.B2(n_18),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_93),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_96),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_46),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_116),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_44),
.B1(n_40),
.B2(n_39),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_102),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_118),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_55),
.B1(n_24),
.B2(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_28),
.B1(n_44),
.B2(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_39),
.B1(n_40),
.B2(n_58),
.Y(n_118)
);

OAI22x1_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_29),
.B1(n_30),
.B2(n_20),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_92),
.B1(n_83),
.B2(n_90),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_38),
.B1(n_41),
.B2(n_46),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_128),
.A2(n_46),
.B(n_85),
.Y(n_133)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_134),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_30),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_133),
.A2(n_139),
.B(n_146),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_67),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_38),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_154),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_30),
.B(n_29),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_72),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_142),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_70),
.B1(n_93),
.B2(n_69),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_15),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_63),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_38),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_70),
.B1(n_69),
.B2(n_63),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

AND2x4_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_101),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_153),
.B(n_133),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_63),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_22),
.Y(n_152)
);

OR2x2_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_22),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_22),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_38),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_165),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_108),
.B1(n_119),
.B2(n_97),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_162),
.A2(n_166),
.B1(n_167),
.B2(n_181),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_155),
.A2(n_119),
.B1(n_112),
.B2(n_117),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_185),
.B1(n_129),
.B2(n_151),
.Y(n_189)
);

AO21x2_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_100),
.B(n_73),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_146),
.B1(n_149),
.B2(n_131),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_149),
.B1(n_131),
.B2(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_121),
.C(n_107),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_170),
.B(n_179),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_121),
.C(n_107),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_134),
.B(n_20),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_184),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_142),
.B1(n_130),
.B2(n_140),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_126),
.B(n_121),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_188),
.B(n_143),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_117),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_126),
.B1(n_71),
.B2(n_41),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_38),
.C(n_100),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_20),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_189),
.A2(n_164),
.B1(n_159),
.B2(n_187),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_191),
.A2(n_197),
.B(n_220),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_195),
.Y(n_230)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_204),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_207),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_10),
.B(n_1),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_10),
.B(n_1),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_34),
.Y(n_201)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_34),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_206),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_34),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_31),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_214),
.Y(n_244)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_31),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_216),
.Y(n_225)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_184),
.C(n_167),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_245),
.C(n_199),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_235),
.B1(n_241),
.B2(n_232),
.Y(n_257)
);

AO22x1_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_165),
.B1(n_175),
.B2(n_161),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_183),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_243),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_200),
.A2(n_175),
.B1(n_165),
.B2(n_31),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_11),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_207),
.A2(n_165),
.B(n_0),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_193),
.B(n_195),
.C(n_215),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_31),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_189),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_209),
.B1(n_211),
.B2(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_203),
.B(n_9),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_26),
.C(n_3),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_220),
.B1(n_197),
.B2(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_252),
.A2(n_254),
.B1(n_257),
.B2(n_234),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_212),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_262),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_202),
.C(n_196),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_258),
.C(n_260),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_196),
.C(n_191),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_203),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_204),
.C(n_198),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_261),
.B(n_237),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_194),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_8),
.B1(n_3),
.B2(n_5),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_266),
.Y(n_273)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_248),
.B(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_221),
.B1(n_235),
.B2(n_242),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_270),
.B1(n_267),
.B2(n_280),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_221),
.B1(n_252),
.B2(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_283),
.Y(n_290)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_282),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_253),
.C(n_258),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_292),
.C(n_298),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_228),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_246),
.C(n_231),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_274),
.B(n_279),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_278),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_232),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_0),
.B(n_5),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_239),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_231),
.C(n_236),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_304),
.Y(n_313)
);

XOR2x2_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_283),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_296),
.B(n_288),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_289),
.A2(n_270),
.B1(n_281),
.B2(n_239),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_272),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_26),
.C(n_7),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_290),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_299),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_285),
.C(n_290),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_317),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_314),
.B(n_310),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_315),
.A2(n_301),
.B(n_300),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_26),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_319),
.B(n_6),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_6),
.Y(n_319)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_322),
.B(n_323),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_301),
.C(n_11),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_6),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_314),
.B(n_14),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_324),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

AOI21xp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_330),
.B(n_326),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_12),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_12),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_335)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_14),
.B(n_15),
.Y(n_336)
);


endmodule