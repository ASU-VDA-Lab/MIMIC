module fake_ibex_856_n_921 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_921);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_921;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_849;
wire n_857;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_696;
wire n_837;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_564;
wire n_562;
wire n_506;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_894;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_50),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_20),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_70),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_46),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_12),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_124),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_45),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_44),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_81),
.B(n_140),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_59),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_85),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_136),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_47),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_7),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_64),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_67),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_5),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_60),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_128),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_103),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_52),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_100),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_145),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_123),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_141),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_94),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_65),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_109),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_17),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_88),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_119),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_132),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_24),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_54),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_126),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_155),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_112),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_99),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_86),
.B(n_19),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_16),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_39),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_40),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_17),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_18),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_101),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_18),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_78),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_16),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_69),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_12),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_142),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_36),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_61),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_171),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_51),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_133),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_0),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_104),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_27),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_7),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_71),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_80),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_8),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_56),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_37),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_113),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_167),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_161),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_117),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_110),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_43),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_116),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_160),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_74),
.B(n_91),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_107),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_134),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_146),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_102),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_55),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_89),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_127),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_42),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_53),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_62),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_66),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_192),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx6p67_ASAP7_75t_R g299 ( 
.A(n_238),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_0),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_293),
.B1(n_181),
.B2(n_201),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_181),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_235),
.Y(n_305)
);

AOI22x1_ASAP7_75t_SL g306 ( 
.A1(n_250),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_306)
);

BUFx8_ASAP7_75t_SL g307 ( 
.A(n_250),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_216),
.B(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_200),
.B(n_6),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_241),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_183),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_210),
.B(n_6),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_235),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_267),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_179),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_193),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_317)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_235),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_235),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_202),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_205),
.B(n_11),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_184),
.A2(n_84),
.B(n_174),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_235),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_13),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_222),
.B(n_13),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_197),
.B(n_14),
.Y(n_330)
);

BUFx8_ASAP7_75t_SL g331 ( 
.A(n_190),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_184),
.A2(n_90),
.B(n_172),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_235),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_194),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_177),
.Y(n_336)
);

AOI22x1_ASAP7_75t_SL g337 ( 
.A1(n_190),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_201),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_219),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_182),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_279),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_15),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_271),
.B(n_21),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_219),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_271),
.B(n_21),
.Y(n_346)
);

OAI22x1_ASAP7_75t_SL g347 ( 
.A1(n_220),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_347)
);

OAI22x1_ASAP7_75t_L g348 ( 
.A1(n_282),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_186),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_191),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_296),
.B(n_25),
.Y(n_351)
);

OA22x2_ASAP7_75t_SL g352 ( 
.A1(n_220),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_196),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_279),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_279),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_206),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_279),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_203),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_229),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_203),
.A2(n_98),
.B(n_169),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_233),
.B(n_29),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_226),
.B(n_30),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g364 ( 
.A1(n_226),
.A2(n_270),
.B(n_263),
.Y(n_364)
);

BUFx12f_ASAP7_75t_L g365 ( 
.A(n_178),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_204),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_180),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_263),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_215),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_232),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_243),
.A2(n_268),
.B1(n_265),
.B2(n_249),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_329),
.Y(n_372)
);

BUFx6f_ASAP7_75t_SL g373 ( 
.A(n_308),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_299),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_364),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

AND2x2_ASAP7_75t_SL g377 ( 
.A(n_302),
.B(n_240),
.Y(n_377)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_209),
.Y(n_379)
);

BUFx16f_ASAP7_75t_R g380 ( 
.A(n_307),
.Y(n_380)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_342),
.B(n_232),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_306),
.A2(n_244),
.B1(n_248),
.B2(n_274),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_312),
.B(n_270),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_328),
.B(n_256),
.C(n_252),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_299),
.A2(n_234),
.B1(n_258),
.B2(n_276),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_312),
.B(n_291),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_257),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_363),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_315),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_302),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g395 ( 
.A1(n_303),
.A2(n_234),
.B1(n_258),
.B2(n_276),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

AND3x2_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_255),
.C(n_289),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_321),
.B(n_259),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_302),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_300),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_301),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_298),
.Y(n_405)
);

INVx11_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_324),
.B(n_272),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_298),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_L g415 ( 
.A(n_328),
.B(n_322),
.C(n_309),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_353),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_353),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

XNOR2x2_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_189),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_326),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_311),
.B(n_280),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_305),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_344),
.B(n_291),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_297),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_297),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_351),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_329),
.B(n_185),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_313),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_L g432 ( 
.A(n_336),
.B(n_195),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_318),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_313),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_301),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_351),
.B(n_207),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_329),
.B(n_188),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_316),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_316),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_336),
.B(n_214),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_319),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_362),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_319),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_330),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g445 ( 
.A(n_342),
.B(n_187),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_300),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

CKINVDCx6p67_ASAP7_75t_R g448 ( 
.A(n_335),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_340),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_340),
.B(n_221),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_331),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_320),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_349),
.B(n_228),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_325),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_338),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_325),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_367),
.B(n_198),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_367),
.B(n_199),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_350),
.B(n_354),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_333),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_333),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_310),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_308),
.A2(n_247),
.B1(n_273),
.B2(n_231),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_341),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_343),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_343),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_366),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_300),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_334),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_366),
.B(n_355),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_357),
.B(n_369),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_355),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_365),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_365),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_356),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_371),
.B(n_247),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_304),
.A2(n_260),
.B1(n_237),
.B2(n_242),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_327),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_358),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_300),
.B(n_295),
.Y(n_482)
);

AND3x2_ASAP7_75t_L g483 ( 
.A(n_352),
.B(n_290),
.C(n_245),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_327),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_439),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_413),
.B(n_208),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_377),
.A2(n_370),
.B1(n_314),
.B2(n_317),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_398),
.B(n_393),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_444),
.B(n_212),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_420),
.B(n_213),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_L g493 ( 
.A(n_422),
.B(n_217),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_464),
.B(n_218),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_408),
.B(n_223),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_404),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_390),
.B(n_246),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_464),
.B(n_224),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_449),
.A2(n_323),
.B(n_288),
.C(n_283),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_225),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_391),
.A2(n_348),
.B1(n_360),
.B2(n_361),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_415),
.B(n_275),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_377),
.B(n_227),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_429),
.B(n_230),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_372),
.B(n_430),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_406),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_435),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_429),
.B(n_236),
.Y(n_510)
);

OAI22x1_ASAP7_75t_L g511 ( 
.A1(n_480),
.A2(n_337),
.B1(n_306),
.B2(n_347),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_432),
.A2(n_337),
.B1(n_281),
.B2(n_287),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_410),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_471),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_437),
.B(n_211),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_454),
.B(n_239),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_389),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_461),
.B(n_251),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_323),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_392),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_469),
.B(n_253),
.Y(n_523)
);

NOR3xp33_ASAP7_75t_L g524 ( 
.A(n_381),
.B(n_266),
.C(n_261),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_438),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_379),
.B(n_262),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_457),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_442),
.B(n_269),
.Y(n_529)
);

NOR3xp33_ASAP7_75t_L g530 ( 
.A(n_381),
.B(n_285),
.C(n_277),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_448),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_373),
.A2(n_479),
.B1(n_399),
.B2(n_426),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_292),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_459),
.B(n_294),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_401),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_384),
.B(n_332),
.Y(n_537)
);

OAI21xp33_ASAP7_75t_L g538 ( 
.A1(n_465),
.A2(n_460),
.B(n_436),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_401),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_374),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_433),
.B(n_284),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_402),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_436),
.B(n_332),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_373),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_402),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

O2A1O1Ixp33_ASAP7_75t_L g548 ( 
.A1(n_478),
.A2(n_361),
.B(n_32),
.C(n_33),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_425),
.B(n_31),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_386),
.B(n_475),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_375),
.B(n_376),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_383),
.B(n_339),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_375),
.B(n_339),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_472),
.Y(n_554)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_421),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_468),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_387),
.B(n_345),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_387),
.B(n_345),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_376),
.B(n_345),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_424),
.B(n_345),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_378),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_472),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_475),
.B(n_34),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_419),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_440),
.B(n_48),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_378),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_423),
.B(n_431),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_450),
.B(n_38),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_476),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_453),
.B(n_115),
.Y(n_570)
);

AOI21xp33_ASAP7_75t_L g571 ( 
.A1(n_514),
.A2(n_456),
.B(n_427),
.Y(n_571)
);

AOI21xp33_ASAP7_75t_L g572 ( 
.A1(n_519),
.A2(n_456),
.B(n_395),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_507),
.B(n_397),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_507),
.B(n_483),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_488),
.B(n_445),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_519),
.B(n_474),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_530),
.A2(n_524),
.B1(n_490),
.B2(n_502),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_L g578 ( 
.A1(n_490),
.A2(n_463),
.B(n_441),
.C(n_481),
.Y(n_578)
);

AO32x1_ASAP7_75t_L g579 ( 
.A1(n_569),
.A2(n_414),
.A3(n_418),
.B1(n_417),
.B2(n_416),
.Y(n_579)
);

OAI21xp33_ASAP7_75t_L g580 ( 
.A1(n_555),
.A2(n_434),
.B(n_431),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_544),
.A2(n_441),
.B(n_447),
.Y(n_581)
);

NOR2x1_ASAP7_75t_L g582 ( 
.A(n_540),
.B(n_406),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_504),
.B(n_527),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_553),
.A2(n_443),
.B(n_434),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_561),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_559),
.A2(n_452),
.B(n_455),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_537),
.A2(n_452),
.B(n_455),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_545),
.B(n_447),
.Y(n_590)
);

O2A1O1Ixp5_ASAP7_75t_L g591 ( 
.A1(n_537),
.A2(n_482),
.B(n_477),
.C(n_462),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_532),
.A2(n_382),
.B1(n_484),
.B2(n_477),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_499),
.A2(n_462),
.B(n_466),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

AO21x1_ASAP7_75t_L g595 ( 
.A1(n_548),
.A2(n_396),
.B(n_412),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_535),
.B(n_382),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_515),
.B(n_382),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_567),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_L g599 ( 
.A(n_505),
.B(n_451),
.C(n_380),
.Y(n_599)
);

AOI21x1_ASAP7_75t_L g600 ( 
.A1(n_521),
.A2(n_407),
.B(n_385),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_530),
.B(n_524),
.C(n_487),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_561),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_497),
.B(n_378),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_L g604 ( 
.A(n_512),
.B(n_451),
.C(n_419),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_495),
.B(n_501),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_545),
.B(n_57),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_536),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_550),
.B(n_388),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_489),
.A2(n_543),
.B(n_542),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_518),
.B(n_522),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_538),
.A2(n_409),
.B(n_396),
.C(n_403),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_550),
.B(n_412),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_546),
.Y(n_613)
);

BUFx8_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

OAI321xp33_ASAP7_75t_L g615 ( 
.A1(n_564),
.A2(n_411),
.A3(n_388),
.B1(n_470),
.B2(n_446),
.C(n_400),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_567),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_531),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_563),
.B(n_63),
.C(n_68),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_550),
.B(n_72),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_561),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_485),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_529),
.B(n_73),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_503),
.B(n_76),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_513),
.B(n_79),
.Y(n_624)
);

AOI21x1_ASAP7_75t_L g625 ( 
.A1(n_560),
.A2(n_446),
.B(n_400),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_549),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_567),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_554),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_566),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_562),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_565),
.A2(n_105),
.B(n_106),
.C(n_111),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_516),
.B(n_520),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_523),
.B(n_175),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_486),
.A2(n_118),
.B(n_120),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_492),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_494),
.B(n_121),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_491),
.B(n_166),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_493),
.A2(n_533),
.B(n_534),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_511),
.B(n_165),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_506),
.A2(n_125),
.B(n_129),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_526),
.B(n_159),
.Y(n_641)
);

AND2x2_ASAP7_75t_SL g642 ( 
.A(n_564),
.B(n_130),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_510),
.B(n_131),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_498),
.B(n_568),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_570),
.A2(n_552),
.B(n_558),
.Y(n_645)
);

A2O1A1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_638),
.A2(n_558),
.B(n_557),
.C(n_570),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_605),
.A2(n_632),
.B(n_609),
.C(n_583),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_601),
.B(n_496),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_577),
.A2(n_509),
.B1(n_525),
.B2(n_517),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_575),
.B(n_500),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_628),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_610),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_572),
.A2(n_528),
.B1(n_556),
.B2(n_547),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_597),
.B(n_541),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_586),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_614),
.Y(n_656)
);

A2O1A1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_578),
.A2(n_148),
.B(n_150),
.C(n_151),
.Y(n_657)
);

AO31x2_ASAP7_75t_L g658 ( 
.A1(n_595),
.A2(n_152),
.A3(n_157),
.B(n_158),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_581),
.A2(n_588),
.B(n_584),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_626),
.B(n_571),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_573),
.B(n_596),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_606),
.B(n_627),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_574),
.B(n_592),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_606),
.B(n_582),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_593),
.A2(n_645),
.B(n_587),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_576),
.B(n_580),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_617),
.B(n_614),
.Y(n_667)
);

AO32x2_ASAP7_75t_L g668 ( 
.A1(n_579),
.A2(n_616),
.A3(n_585),
.B1(n_615),
.B2(n_642),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_613),
.B(n_644),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_619),
.B(n_604),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_611),
.A2(n_623),
.B(n_624),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_608),
.A2(n_612),
.B1(n_639),
.B2(n_622),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_620),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_633),
.A2(n_603),
.B(n_590),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_629),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_621),
.A2(n_635),
.B(n_641),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_594),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_636),
.A2(n_640),
.B(n_634),
.C(n_618),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_643),
.A2(n_637),
.B(n_631),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_599),
.B(n_629),
.Y(n_680)
);

AO31x2_ASAP7_75t_L g681 ( 
.A1(n_579),
.A2(n_630),
.A3(n_598),
.B(n_602),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_579),
.A2(n_589),
.B(n_602),
.Y(n_682)
);

CKINVDCx11_ASAP7_75t_R g683 ( 
.A(n_629),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_602),
.A2(n_377),
.B1(n_577),
.B2(n_610),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_601),
.B(n_488),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_601),
.B(n_488),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_601),
.B(n_488),
.Y(n_687)
);

AOI211x1_ASAP7_75t_L g688 ( 
.A1(n_595),
.A2(n_583),
.B(n_597),
.C(n_596),
.Y(n_688)
);

OAI21xp33_ASAP7_75t_L g689 ( 
.A1(n_605),
.A2(n_473),
.B(n_456),
.Y(n_689)
);

BUFx4f_ASAP7_75t_L g690 ( 
.A(n_642),
.Y(n_690)
);

AOI21x1_ASAP7_75t_L g691 ( 
.A1(n_625),
.A2(n_600),
.B(n_595),
.Y(n_691)
);

AO31x2_ASAP7_75t_L g692 ( 
.A1(n_595),
.A2(n_499),
.A3(n_537),
.B(n_544),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_586),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_601),
.B(n_488),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_604),
.B(n_456),
.C(n_577),
.Y(n_695)
);

OAI21xp33_ASAP7_75t_L g696 ( 
.A1(n_605),
.A2(n_473),
.B(n_456),
.Y(n_696)
);

AOI21x1_ASAP7_75t_L g697 ( 
.A1(n_625),
.A2(n_600),
.B(n_595),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_601),
.B(n_488),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_601),
.B(n_488),
.Y(n_699)
);

AO31x2_ASAP7_75t_L g700 ( 
.A1(n_595),
.A2(n_499),
.A3(n_537),
.B(n_544),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_601),
.B(n_488),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_591),
.A2(n_537),
.B(n_544),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_628),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_601),
.B(n_488),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_572),
.B(n_555),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_638),
.A2(n_605),
.B(n_632),
.C(n_507),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_575),
.B(n_480),
.Y(n_707)
);

AOI21x1_ASAP7_75t_L g708 ( 
.A1(n_625),
.A2(n_600),
.B(n_595),
.Y(n_708)
);

AO22x2_ASAP7_75t_L g709 ( 
.A1(n_592),
.A2(n_386),
.B1(n_337),
.B2(n_601),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_614),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_601),
.A2(n_642),
.B1(n_487),
.B2(n_592),
.Y(n_711)
);

CKINVDCx11_ASAP7_75t_R g712 ( 
.A(n_617),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_601),
.B(n_488),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_601),
.B(n_488),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_585),
.B(n_616),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_628),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_614),
.Y(n_717)
);

NAND2x1p5_ASAP7_75t_L g718 ( 
.A(n_617),
.B(n_540),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_586),
.Y(n_719)
);

AO31x2_ASAP7_75t_L g720 ( 
.A1(n_595),
.A2(n_499),
.A3(n_537),
.B(n_544),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_607),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_638),
.A2(n_605),
.B(n_632),
.C(n_507),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_601),
.B(n_488),
.Y(n_723)
);

AO31x2_ASAP7_75t_L g724 ( 
.A1(n_595),
.A2(n_499),
.A3(n_537),
.B(n_544),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_628),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_601),
.B(n_488),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_651),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_706),
.A2(n_722),
.B(n_647),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_682),
.A2(n_691),
.B(n_697),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_685),
.B(n_686),
.Y(n_731)
);

NOR2x1_ASAP7_75t_R g732 ( 
.A(n_712),
.B(n_717),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_673),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_690),
.A2(n_709),
.B1(n_711),
.B2(n_705),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_656),
.Y(n_735)
);

AOI21xp5_ASAP7_75t_L g736 ( 
.A1(n_678),
.A2(n_671),
.B(n_679),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_SL g737 ( 
.A1(n_687),
.A2(n_698),
.B1(n_701),
.B2(n_726),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_694),
.B(n_699),
.Y(n_738)
);

AO21x2_ASAP7_75t_L g739 ( 
.A1(n_708),
.A2(n_665),
.B(n_702),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_704),
.B(n_713),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_718),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_684),
.A2(n_714),
.B1(n_723),
.B2(n_672),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_689),
.A2(n_696),
.B1(n_695),
.B2(n_670),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_710),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_664),
.B(n_721),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_703),
.Y(n_746)
);

CKINVDCx8_ASAP7_75t_R g747 ( 
.A(n_667),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_664),
.B(n_715),
.Y(n_748)
);

AOI32xp33_ASAP7_75t_L g749 ( 
.A1(n_660),
.A2(n_648),
.A3(n_663),
.B1(n_654),
.B2(n_707),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_683),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_669),
.B(n_725),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_661),
.B(n_716),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_672),
.A2(n_662),
.B1(n_688),
.B2(n_653),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_666),
.A2(n_650),
.B1(n_676),
.B2(n_680),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_675),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_655),
.B(n_719),
.Y(n_756)
);

AO31x2_ASAP7_75t_L g757 ( 
.A1(n_646),
.A2(n_657),
.A3(n_674),
.B(n_649),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_677),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_693),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_693),
.B(n_719),
.Y(n_760)
);

AOI222xp33_ASAP7_75t_L g761 ( 
.A1(n_668),
.A2(n_692),
.B1(n_700),
.B2(n_720),
.C1(n_724),
.C2(n_658),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_724),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_681),
.B(n_652),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_678),
.A2(n_551),
.B(n_671),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_652),
.B(n_664),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_683),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_652),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_693),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_656),
.Y(n_769)
);

BUFx8_ASAP7_75t_L g770 ( 
.A(n_717),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_656),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_683),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_683),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_690),
.A2(n_711),
.B1(n_652),
.B2(n_642),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_651),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_690),
.A2(n_711),
.B1(n_652),
.B2(n_642),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_652),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_693),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_718),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_685),
.B(n_480),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_682),
.A2(n_659),
.A3(n_595),
.B(n_499),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_685),
.B(n_480),
.Y(n_782)
);

AO21x1_ASAP7_75t_L g783 ( 
.A1(n_684),
.A2(n_711),
.B(n_670),
.Y(n_783)
);

OR2x6_ASAP7_75t_L g784 ( 
.A(n_717),
.B(n_386),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_652),
.B(n_490),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_767),
.Y(n_786)
);

AO21x2_ASAP7_75t_L g787 ( 
.A1(n_729),
.A2(n_736),
.B(n_764),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_760),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_740),
.B(n_742),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_739),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_731),
.B(n_738),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_763),
.B(n_748),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_730),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_727),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_746),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_740),
.B(n_752),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_785),
.B(n_749),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_775),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_733),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_751),
.Y(n_801)
);

INVx6_ASAP7_75t_L g802 ( 
.A(n_759),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_728),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_777),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_781),
.Y(n_805)
);

HB1xp67_ASAP7_75t_SL g806 ( 
.A(n_770),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_784),
.B(n_737),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_781),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_750),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_781),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_758),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_762),
.Y(n_813)
);

INVxp33_ASAP7_75t_L g814 ( 
.A(n_732),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_743),
.A2(n_780),
.B(n_782),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_770),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_774),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_741),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_742),
.B(n_734),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_754),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_779),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_807),
.A2(n_737),
.B1(n_774),
.B2(n_776),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_808),
.B(n_761),
.Y(n_823)
);

AND2x4_ASAP7_75t_SL g824 ( 
.A(n_788),
.B(n_778),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_795),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_808),
.B(n_761),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_789),
.B(n_801),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_789),
.B(n_776),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_805),
.B(n_783),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_786),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_811),
.B(n_753),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_817),
.B(n_743),
.Y(n_832)
);

OR2x2_ASAP7_75t_L g833 ( 
.A(n_798),
.B(n_792),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_813),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_787),
.B(n_757),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_825),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_830),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_833),
.B(n_816),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_823),
.B(n_793),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_830),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_823),
.B(n_826),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_833),
.B(n_814),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_826),
.B(n_790),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_827),
.B(n_820),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_834),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_835),
.B(n_787),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_834),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_835),
.B(n_787),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_836),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_845),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_846),
.B(n_831),
.Y(n_851)
);

AND2x4_ASAP7_75t_SL g852 ( 
.A(n_837),
.B(n_788),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_841),
.B(n_819),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_840),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_841),
.B(n_819),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_848),
.B(n_829),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_838),
.B(n_732),
.Y(n_857)
);

NAND2x1p5_ASAP7_75t_L g858 ( 
.A(n_847),
.B(n_788),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_840),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_841),
.B(n_832),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_860),
.B(n_839),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_854),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_856),
.B(n_848),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_856),
.B(n_848),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_849),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_852),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_860),
.B(n_851),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_850),
.B(n_843),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_857),
.A2(n_822),
.B1(n_842),
.B2(n_815),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_863),
.B(n_864),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_863),
.B(n_843),
.Y(n_871)
);

OAI21xp33_ASAP7_75t_L g872 ( 
.A1(n_868),
.A2(n_855),
.B(n_853),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_865),
.Y(n_873)
);

AOI32xp33_ASAP7_75t_L g874 ( 
.A1(n_866),
.A2(n_852),
.A3(n_847),
.B1(n_850),
.B2(n_800),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_865),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_862),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_864),
.B(n_859),
.Y(n_877)
);

O2A1O1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_867),
.A2(n_784),
.B(n_791),
.C(n_810),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_861),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_868),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_876),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_875),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_879),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_877),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_884),
.B(n_872),
.Y(n_885)
);

AOI211xp5_ASAP7_75t_SL g886 ( 
.A1(n_883),
.A2(n_869),
.B(n_806),
.C(n_828),
.Y(n_886)
);

AOI211x1_ASAP7_75t_SL g887 ( 
.A1(n_882),
.A2(n_878),
.B(n_874),
.C(n_844),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_SL g888 ( 
.A(n_887),
.B(n_772),
.C(n_809),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_L g889 ( 
.A(n_886),
.B(n_772),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_889),
.B(n_885),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_L g891 ( 
.A(n_888),
.B(n_881),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_890),
.B(n_880),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_891),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_892),
.Y(n_894)
);

NOR2x1_ASAP7_75t_SL g895 ( 
.A(n_893),
.B(n_766),
.Y(n_895)
);

AOI22x1_ASAP7_75t_L g896 ( 
.A1(n_894),
.A2(n_735),
.B1(n_771),
.B2(n_769),
.Y(n_896)
);

XNOR2xp5_ASAP7_75t_L g897 ( 
.A(n_895),
.B(n_773),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_894),
.B(n_882),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_896),
.B(n_898),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_897),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_897),
.B(n_802),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_897),
.Y(n_902)
);

XNOR2x1_ASAP7_75t_L g903 ( 
.A(n_897),
.B(n_784),
.Y(n_903)
);

XOR2xp5_ASAP7_75t_L g904 ( 
.A(n_903),
.B(n_747),
.Y(n_904)
);

OAI21xp33_ASAP7_75t_L g905 ( 
.A1(n_901),
.A2(n_870),
.B(n_818),
.Y(n_905)
);

OAI22x1_ASAP7_75t_L g906 ( 
.A1(n_902),
.A2(n_802),
.B1(n_821),
.B2(n_870),
.Y(n_906)
);

NOR4xp25_ASAP7_75t_L g907 ( 
.A(n_900),
.B(n_899),
.C(n_802),
.D(n_794),
.Y(n_907)
);

AOI222xp33_ASAP7_75t_L g908 ( 
.A1(n_900),
.A2(n_802),
.B1(n_873),
.B2(n_794),
.C1(n_799),
.C2(n_796),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_901),
.A2(n_875),
.B1(n_858),
.B2(n_788),
.Y(n_909)
);

OAI22x1_ASAP7_75t_L g910 ( 
.A1(n_902),
.A2(n_765),
.B1(n_745),
.B2(n_858),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_907),
.A2(n_904),
.B(n_908),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_906),
.A2(n_871),
.B1(n_745),
.B2(n_755),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_905),
.A2(n_871),
.B1(n_797),
.B2(n_824),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_910),
.B(n_768),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_911),
.A2(n_909),
.B(n_756),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_914),
.A2(n_803),
.B(n_804),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_912),
.A2(n_796),
.B(n_799),
.Y(n_917)
);

OAI21xp33_ASAP7_75t_L g918 ( 
.A1(n_915),
.A2(n_916),
.B(n_913),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_917),
.B(n_812),
.Y(n_919)
);

OR2x6_ASAP7_75t_L g920 ( 
.A(n_918),
.B(n_919),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_920),
.A2(n_812),
.B(n_768),
.Y(n_921)
);


endmodule