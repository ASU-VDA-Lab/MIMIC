module fake_jpeg_31808_n_400 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_400);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_400;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_12),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_49),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_11),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_67),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_62),
.B(n_78),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_25),
.A2(n_33),
.B(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_0),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_74),
.B(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_39),
.B(n_0),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_86),
.C(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_79),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_81),
.Y(n_122)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_83),
.Y(n_124)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_87),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_1),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_89),
.Y(n_147)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_32),
.A2(n_1),
.B(n_2),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_28),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_37),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_19),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_32),
.B(n_21),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_107),
.B(n_64),
.C(n_68),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_29),
.B1(n_35),
.B2(n_37),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_126),
.B1(n_146),
.B2(n_74),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_116),
.Y(n_158)
);

INVx2_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_110),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_29),
.B(n_5),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_21),
.B(n_6),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_65),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_52),
.A2(n_38),
.B1(n_22),
.B2(n_15),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_84),
.A2(n_42),
.B1(n_22),
.B2(n_17),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_127),
.A2(n_141),
.B1(n_144),
.B2(n_131),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_42),
.B(n_17),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_68),
.B(n_8),
.C(n_9),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_79),
.A2(n_16),
.B1(n_36),
.B2(n_19),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_83),
.A2(n_42),
.B1(n_16),
.B2(n_18),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_72),
.A2(n_36),
.B1(n_18),
.B2(n_21),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_150),
.B1(n_77),
.B2(n_85),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_49),
.A2(n_21),
.B1(n_6),
.B2(n_7),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_51),
.A2(n_21),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_59),
.B1(n_53),
.B2(n_57),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_167),
.B1(n_169),
.B2(n_179),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_156),
.A2(n_174),
.B1(n_186),
.B2(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_69),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_157),
.B(n_163),
.Y(n_206)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_65),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_164),
.Y(n_207)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_140),
.B1(n_150),
.B2(n_143),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_177),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_110),
.B(n_4),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_190),
.C(n_138),
.Y(n_208)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_98),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_8),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_8),
.B1(n_9),
.B2(n_141),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_137),
.A2(n_8),
.B1(n_125),
.B2(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_188),
.B1(n_132),
.B2(n_102),
.Y(n_204)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_111),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_184),
.B(n_100),
.Y(n_219)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_185),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_106),
.A2(n_125),
.B1(n_124),
.B2(n_142),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_121),
.A2(n_118),
.B1(n_129),
.B2(n_136),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_191),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_113),
.B(n_145),
.C(n_130),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_98),
.A2(n_136),
.B1(n_130),
.B2(n_105),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_102),
.C(n_138),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_202),
.C(n_153),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_132),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_203),
.B(n_220),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_208),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_128),
.B1(n_144),
.B2(n_100),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

INVx11_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_128),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_128),
.B1(n_114),
.B2(n_100),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_215),
.A2(n_159),
.B1(n_164),
.B2(n_204),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_165),
.B(n_114),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_114),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_177),
.B(n_149),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_160),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_149),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_190),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_196),
.A2(n_156),
.B1(n_154),
.B2(n_186),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_253),
.B1(n_210),
.B2(n_199),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_246),
.C(n_249),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_225),
.B(n_194),
.C(n_154),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_237),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_179),
.B(n_174),
.C(n_170),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_152),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_242),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_167),
.B1(n_188),
.B2(n_172),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_196),
.B1(n_217),
.B2(n_210),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_171),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_182),
.B(n_189),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_184),
.B(n_185),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_178),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_191),
.C(n_181),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_168),
.B(n_160),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_200),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_259),
.B1(n_268),
.B2(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_257),
.A2(n_235),
.B1(n_251),
.B2(n_227),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_210),
.B1(n_195),
.B2(n_164),
.Y(n_259)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_265),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_210),
.B1(n_201),
.B2(n_207),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_233),
.A2(n_207),
.B1(n_201),
.B2(n_222),
.Y(n_270)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_220),
.B1(n_207),
.B2(n_205),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_235),
.B1(n_253),
.B2(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_278),
.Y(n_288)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_226),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_228),
.C(n_230),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_246),
.C(n_249),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_228),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_295),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_287),
.A2(n_298),
.B1(n_264),
.B2(n_257),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_254),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_294),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_234),
.C(n_245),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_252),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_272),
.B1(n_262),
.B2(n_264),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_261),
.A2(n_232),
.B(n_247),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_249),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_261),
.A2(n_232),
.B(n_247),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

AO21x2_ASAP7_75t_L g298 ( 
.A1(n_255),
.A2(n_248),
.B(n_233),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_255),
.A2(n_235),
.B(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_263),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_314),
.C(n_318),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_280),
.A2(n_259),
.B1(n_256),
.B2(n_268),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_303),
.A2(n_305),
.B1(n_298),
.B2(n_297),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_288),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_319),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_308),
.B(n_320),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_270),
.B1(n_298),
.B2(n_287),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_274),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_310),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_311),
.A2(n_298),
.B(n_294),
.Y(n_335)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_262),
.C(n_276),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_231),
.B1(n_241),
.B2(n_227),
.Y(n_315)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_281),
.A2(n_275),
.B1(n_263),
.B2(n_250),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_321),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_295),
.C(n_276),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_335),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_307),
.Y(n_323)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_323),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_311),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_338),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_300),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_316),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_301),
.B(n_318),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_332),
.B(n_334),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_309),
.A2(n_298),
.B(n_290),
.C(n_279),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_336),
.A2(n_279),
.B(n_284),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_289),
.Y(n_337)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_R g338 ( 
.A(n_313),
.B(n_265),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_340),
.B(n_325),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_302),
.C(n_305),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_347),
.C(n_330),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_313),
.B(n_303),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_345),
.A2(n_336),
.B(n_334),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_310),
.C(n_236),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_333),
.Y(n_348)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_310),
.Y(n_350)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_325),
.Y(n_353)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_353),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_344),
.B(n_324),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_358),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_342),
.C(n_340),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_341),
.B(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_363),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_361),
.A2(n_364),
.B(n_351),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_347),
.B(n_306),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_345),
.A2(n_322),
.B(n_336),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_350),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_365),
.Y(n_368)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_366),
.A2(n_373),
.B(n_364),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_356),
.A2(n_346),
.B(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_367),
.Y(n_377)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_375),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_374),
.C(n_355),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_361),
.A2(n_348),
.B(n_343),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_343),
.C(n_349),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_362),
.B(n_283),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_380),
.C(n_382),
.Y(n_388)
);

AOI31xp33_ASAP7_75t_L g385 ( 
.A1(n_379),
.A2(n_271),
.A3(n_277),
.B(n_265),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_355),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_365),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_372),
.B(n_336),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_339),
.C(n_289),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_368),
.A2(n_312),
.B1(n_236),
.B2(n_269),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_376),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_386),
.Y(n_391)
);

AO21x1_ASAP7_75t_L g392 ( 
.A1(n_385),
.A2(n_389),
.B(n_277),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_377),
.A2(n_273),
.B(n_267),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_387),
.A2(n_376),
.B(n_260),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_381),
.A2(n_260),
.B(n_271),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_390),
.A2(n_393),
.B(n_222),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_392),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_226),
.C(n_221),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_218),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_213),
.B(n_221),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_395),
.B(n_200),
.Y(n_397)
);

OAI321xp33_ASAP7_75t_L g399 ( 
.A1(n_397),
.A2(n_398),
.A3(n_396),
.B1(n_216),
.B2(n_193),
.C(n_218),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_399),
.B(n_193),
.C(n_216),
.Y(n_400)
);


endmodule