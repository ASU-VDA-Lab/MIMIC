module fake_jpeg_20289_n_308 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_20),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_29),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_49),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_32),
.B1(n_25),
.B2(n_28),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_19),
.B1(n_34),
.B2(n_32),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_60),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_23),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_40),
.CI(n_39),
.CON(n_83),
.SN(n_83)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_24),
.B1(n_29),
.B2(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_65),
.B1(n_42),
.B2(n_43),
.Y(n_81)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_24),
.B1(n_21),
.B2(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_39),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_69),
.C(n_87),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_39),
.C(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_24),
.B1(n_21),
.B2(n_20),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_70),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_91),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_79),
.B1(n_19),
.B2(n_34),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_28),
.B1(n_25),
.B2(n_32),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_90),
.B(n_52),
.C(n_35),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_57),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_89),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_39),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_95),
.Y(n_144)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_114),
.B1(n_86),
.B2(n_68),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_109),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_106),
.A2(n_86),
.B1(n_76),
.B2(n_35),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_116),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_43),
.C(n_46),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_72),
.C(n_94),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_38),
.B1(n_35),
.B2(n_19),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_75),
.C(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_22),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_80),
.B(n_38),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_22),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_22),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_23),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_23),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_83),
.B(n_77),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_140),
.B(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_66),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_135),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_88),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_72),
.C(n_76),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_97),
.B(n_33),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_141),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_86),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_95),
.B1(n_102),
.B2(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_107),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_26),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_30),
.B1(n_26),
.B2(n_23),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_33),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_106),
.B1(n_112),
.B2(n_68),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_26),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_151),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_121),
.B(n_95),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_153),
.A2(n_163),
.B(n_165),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_172),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_99),
.B(n_116),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_99),
.B(n_106),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_106),
.B(n_108),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_170),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_106),
.B1(n_100),
.B2(n_112),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_122),
.A2(n_96),
.B1(n_38),
.B2(n_62),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_172),
.A2(n_139),
.B1(n_147),
.B2(n_128),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_26),
.B(n_30),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_181),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_177),
.B(n_31),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_30),
.B(n_26),
.C(n_23),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_126),
.A2(n_30),
.B(n_26),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_31),
.B(n_23),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_126),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_142),
.C(n_137),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_192),
.C(n_154),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_140),
.B1(n_143),
.B2(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_175),
.B1(n_159),
.B2(n_181),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_170),
.B1(n_155),
.B2(n_169),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_179),
.B(n_159),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_141),
.C(n_123),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_131),
.Y(n_193)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_123),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_201),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_151),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_125),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_33),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_18),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_18),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_208),
.B(n_210),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_23),
.Y(n_209)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_216),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_204),
.A2(n_165),
.B1(n_182),
.B2(n_152),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_196),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_215),
.C(n_223),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_162),
.C(n_164),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_162),
.C(n_155),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_229),
.B(n_195),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_159),
.C(n_160),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_215),
.C(n_213),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_160),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_233),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_31),
.B(n_2),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_201),
.B(n_5),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_206),
.B(n_5),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_205),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_212),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_186),
.Y(n_244)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_198),
.C(n_204),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_247),
.C(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_251),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_196),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_191),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_227),
.B1(n_195),
.B2(n_221),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_189),
.B1(n_202),
.B2(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_266),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_259),
.B1(n_262),
.B2(n_261),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_211),
.B(n_189),
.C(n_244),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_225),
.B1(n_232),
.B2(n_207),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_253),
.A2(n_229),
.B1(n_203),
.B2(n_9),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_7),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_203),
.B1(n_8),
.B2(n_9),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_237),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_237),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_268),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_242),
.B(n_245),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_275),
.B(n_10),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_242),
.B(n_247),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_281),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_7),
.B(n_8),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_254),
.C(n_257),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_286),
.C(n_12),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_261),
.C(n_267),
.Y(n_286)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_11),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_278),
.B(n_270),
.Y(n_293)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_296),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_11),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_283),
.A3(n_291),
.B1(n_287),
.B2(n_286),
.C1(n_284),
.C2(n_13),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_295),
.A3(n_299),
.B1(n_303),
.B2(n_300),
.C1(n_298),
.C2(n_16),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_12),
.B(n_13),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_14),
.B(n_15),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_304),
.A2(n_305),
.B(n_301),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_14),
.B(n_15),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_15),
.Y(n_308)
);


endmodule