module fake_jpeg_30798_n_534 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_63),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_0),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_76),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_20),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_96),
.Y(n_105)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_83),
.B(n_21),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_32),
.B(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_100),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_30),
.B1(n_43),
.B2(n_42),
.Y(n_160)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_2),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_28),
.B(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_35),
.Y(n_138)
);

NOR2x1_ASAP7_75t_R g112 ( 
.A(n_93),
.B(n_47),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_138),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_47),
.B1(n_38),
.B2(n_44),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_122),
.B1(n_88),
.B2(n_43),
.Y(n_169)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_50),
.A2(n_47),
.B1(n_38),
.B2(n_44),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_60),
.A2(n_45),
.B1(n_28),
.B2(n_35),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_123),
.A2(n_41),
.B1(n_26),
.B2(n_25),
.Y(n_221)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_132),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_54),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_142),
.B(n_148),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_55),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_66),
.A2(n_3),
.B(n_4),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_45),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_98),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_160),
.A2(n_41),
.B1(n_26),
.B2(n_25),
.Y(n_218)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_75),
.A2(n_30),
.B1(n_29),
.B2(n_43),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_61),
.B1(n_53),
.B2(n_95),
.Y(n_187)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_165),
.Y(n_245)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_105),
.B(n_30),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_189),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_177),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_192),
.Y(n_243)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_79),
.B1(n_86),
.B2(n_84),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_182),
.A2(n_218),
.B1(n_225),
.B2(n_141),
.Y(n_240)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_185),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_130),
.A2(n_80),
.B1(n_70),
.B2(n_69),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g248 ( 
.A1(n_186),
.A2(n_163),
.B1(n_161),
.B2(n_139),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_164),
.B(n_113),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_29),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_125),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_102),
.B(n_58),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_191),
.B(n_194),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_108),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_102),
.B(n_61),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_116),
.A2(n_38),
.B1(n_24),
.B2(n_44),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_200),
.B(n_49),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_133),
.B(n_53),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_214),
.Y(n_254)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_114),
.B(n_42),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_114),
.B(n_42),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_124),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_133),
.B(n_29),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_219),
.Y(n_269)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_216),
.Y(n_261)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_222),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_154),
.B(n_41),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_154),
.B(n_49),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_21),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_108),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_224),
.Y(n_267)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_121),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_143),
.A2(n_51),
.B1(n_26),
.B2(n_25),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_233),
.A2(n_250),
.B(n_215),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_141),
.B1(n_130),
.B2(n_163),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_248),
.B1(n_173),
.B2(n_179),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_122),
.B(n_21),
.C(n_49),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_237),
.B(n_268),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_240),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_241),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_183),
.A2(n_146),
.B1(n_129),
.B2(n_126),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_244),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_174),
.A2(n_103),
.B1(n_49),
.B2(n_158),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_174),
.B(n_103),
.C(n_158),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_252),
.B(n_260),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_185),
.A2(n_151),
.B1(n_161),
.B2(n_147),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_255),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_200),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_182),
.A2(n_147),
.B1(n_81),
.B2(n_5),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_272),
.B1(n_186),
.B2(n_187),
.Y(n_276)
);

AO22x1_ASAP7_75t_L g271 ( 
.A1(n_221),
.A2(n_49),
.B1(n_4),
.B2(n_5),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_212),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_225),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_209),
.B(n_6),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_243),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_233),
.B1(n_232),
.B2(n_250),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_221),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_277),
.B(n_278),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_177),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_170),
.B1(n_171),
.B2(n_195),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_279),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_288),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_261),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_234),
.B(n_167),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_284),
.B(n_285),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_234),
.B(n_208),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_227),
.B(n_241),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_286),
.B(n_289),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_287),
.A2(n_302),
.B(n_253),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_198),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_267),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_297),
.Y(n_322)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_260),
.B(n_175),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_293),
.B(n_294),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_184),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_228),
.B(n_211),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_295),
.B(n_299),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_197),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_228),
.B(n_188),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_226),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_271),
.A2(n_190),
.B(n_223),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_268),
.A2(n_181),
.B1(n_176),
.B2(n_199),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_303),
.A2(n_313),
.B1(n_266),
.B2(n_251),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_214),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_306),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_252),
.B(n_224),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_228),
.B(n_203),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_314),
.Y(n_321)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_312),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_248),
.A2(n_165),
.B1(n_178),
.B2(n_166),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_239),
.B1(n_247),
.B2(n_226),
.Y(n_350)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_240),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_9),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_237),
.B(n_9),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_318),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_232),
.B(n_273),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_245),
.B(n_9),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_230),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_323),
.A2(n_324),
.B1(n_333),
.B2(n_337),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_296),
.A2(n_232),
.B1(n_265),
.B2(n_259),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_259),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_315),
.C(n_283),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_295),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_330),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_275),
.A2(n_263),
.B(n_242),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_329),
.A2(n_336),
.B(n_340),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_299),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_276),
.A2(n_263),
.B1(n_256),
.B2(n_242),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_287),
.A2(n_253),
.B(n_245),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_334),
.A2(n_347),
.B(n_312),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_318),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_338),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_282),
.A2(n_256),
.B1(n_231),
.B2(n_249),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_310),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_247),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_339),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_275),
.A2(n_231),
.B(n_249),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_291),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_346),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_302),
.A2(n_239),
.B(n_258),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_307),
.B1(n_311),
.B2(n_303),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_351),
.A2(n_288),
.B1(n_311),
.B2(n_300),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_317),
.A2(n_230),
.B(n_258),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_353),
.A2(n_306),
.B(n_294),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_356),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

A2O1A1O1Ixp25_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_286),
.B(n_278),
.C(n_289),
.D(n_293),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_383),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_SL g362 ( 
.A1(n_334),
.A2(n_314),
.B(n_316),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_362),
.A2(n_368),
.B1(n_385),
.B2(n_348),
.Y(n_399)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_364),
.A2(n_333),
.B1(n_337),
.B2(n_351),
.Y(n_397)
);

OAI21xp33_ASAP7_75t_SL g368 ( 
.A1(n_336),
.A2(n_342),
.B(n_353),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_358),
.Y(n_369)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_371),
.A2(n_329),
.B(n_353),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_373),
.C(n_377),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_281),
.C(n_284),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_320),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_375),
.Y(n_400)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_322),
.B(n_285),
.C(n_290),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_339),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_390),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_309),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_301),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_382),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_379),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_321),
.B(n_343),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_386),
.C(n_377),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_320),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_381),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_321),
.B(n_298),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_307),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_332),
.C(n_331),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_305),
.Y(n_387)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_388),
.A2(n_391),
.B(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_389),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_328),
.B(n_292),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_348),
.A2(n_266),
.B1(n_251),
.B2(n_229),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_328),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_370),
.A2(n_323),
.B1(n_351),
.B2(n_339),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_397),
.B1(n_367),
.B2(n_354),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_399),
.A2(n_403),
.B(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_384),
.A2(n_348),
.B1(n_332),
.B2(n_326),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_404),
.A2(n_410),
.B1(n_414),
.B2(n_419),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_388),
.A2(n_348),
.B(n_340),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_390),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_341),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_330),
.Y(n_409)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

OAI22x1_ASAP7_75t_L g410 ( 
.A1(n_391),
.A2(n_376),
.B1(n_367),
.B2(n_392),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_338),
.B1(n_350),
.B2(n_344),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_322),
.Y(n_415)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_415),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_343),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_421),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_392),
.A2(n_335),
.B1(n_352),
.B2(n_327),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_329),
.C(n_327),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_423),
.C(n_421),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_345),
.C(n_352),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_365),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_369),
.C(n_363),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_398),
.B(n_386),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_426),
.B(n_417),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_437),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_450),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_382),
.C(n_378),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_435),
.C(n_422),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_404),
.A2(n_413),
.B1(n_399),
.B2(n_410),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_434),
.A2(n_438),
.B1(n_420),
.B2(n_414),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_371),
.C(n_365),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_400),
.B(n_345),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_413),
.A2(n_364),
.B1(n_379),
.B2(n_324),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_395),
.A2(n_383),
.B1(n_389),
.B2(n_393),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_444),
.Y(n_455)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_440),
.Y(n_454)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_405),
.Y(n_444)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_360),
.B1(n_341),
.B2(n_355),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_446),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_407),
.B(n_355),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_447),
.Y(n_465)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

BUFx12_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_449),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_409),
.B(n_346),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_451),
.B(n_467),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_443),
.C(n_432),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_423),
.C(n_394),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_458),
.C(n_459),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_394),
.C(n_416),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_406),
.C(n_398),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_428),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_419),
.C(n_401),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_434),
.C(n_443),
.Y(n_483)
);

FAx1_ASAP7_75t_SL g463 ( 
.A(n_441),
.B(n_415),
.CI(n_420),
.CON(n_463),
.SN(n_463)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_446),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_412),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_408),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_469),
.B(n_470),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_439),
.B(n_418),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_464),
.A2(n_427),
.B1(n_425),
.B2(n_432),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_476),
.Y(n_491)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_475),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_441),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_477),
.B(n_483),
.Y(n_498)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_480),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_465),
.B(n_436),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_486),
.Y(n_499)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_454),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_484),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g485 ( 
.A1(n_455),
.A2(n_444),
.B(n_430),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_487),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_438),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_457),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_450),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_478),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_463),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_10),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_467),
.C(n_459),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_492),
.B(n_12),
.C(n_14),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_17),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_486),
.B(n_470),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_501),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_481),
.A2(n_462),
.B1(n_468),
.B2(n_460),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_497),
.A2(n_472),
.B1(n_449),
.B2(n_11),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_469),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_485),
.A2(n_456),
.B(n_445),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_502),
.B(n_9),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_490),
.A2(n_463),
.B1(n_473),
.B2(n_349),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_508),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_498),
.A2(n_473),
.B(n_471),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_509),
.C(n_510),
.Y(n_514)
);

OAI321xp33_ASAP7_75t_L g506 ( 
.A1(n_493),
.A2(n_449),
.A3(n_472),
.B1(n_451),
.B2(n_349),
.C(n_229),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_506),
.A2(n_507),
.B1(n_494),
.B2(n_16),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_10),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_499),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_512),
.C(n_513),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_509),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_515),
.B(n_520),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_497),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_500),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_518),
.B(n_505),
.Y(n_524)
);

BUFx4f_ASAP7_75t_SL g520 ( 
.A(n_512),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_519),
.A2(n_491),
.B(n_495),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_523),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_524),
.B(n_514),
.C(n_492),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_521),
.B(n_501),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_528),
.B(n_519),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_525),
.Y(n_528)
);

NAND4xp25_ASAP7_75t_SL g530 ( 
.A(n_529),
.B(n_520),
.C(n_516),
.D(n_499),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_530),
.A2(n_510),
.B(n_16),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_531),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_15),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_17),
.B(n_400),
.Y(n_534)
);


endmodule