module fake_jpeg_26921_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_24),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_60),
.Y(n_67)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_22),
.B1(n_29),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_22),
.B1(n_29),
.B2(n_28),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_23),
.B1(n_39),
.B2(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_61),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_55),
.Y(n_81)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_23),
.B1(n_20),
.B2(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_77),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_23),
.B1(n_40),
.B2(n_18),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_81),
.B1(n_52),
.B2(n_62),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_16),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_78),
.Y(n_106)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_90),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_25),
.B1(n_19),
.B2(n_16),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_32),
.B1(n_30),
.B2(n_40),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_40),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_56),
.B(n_54),
.Y(n_96)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_19),
.B1(n_40),
.B2(n_32),
.Y(n_87)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_88),
.A2(n_61),
.B1(n_30),
.B2(n_32),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_52),
.B1(n_62),
.B2(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_97),
.B1(n_105),
.B2(n_66),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_65),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_96),
.B(n_41),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_69),
.B(n_14),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_100),
.B(n_104),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_64),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_50),
.C(n_37),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_69),
.B(n_13),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_50),
.B1(n_62),
.B2(n_52),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_81),
.B1(n_77),
.B2(n_84),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_115),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_42),
.B1(n_37),
.B2(n_41),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_42),
.B1(n_41),
.B2(n_34),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_41),
.A3(n_34),
.B1(n_31),
.B2(n_17),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_78),
.B(n_41),
.C(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_92),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_41),
.B1(n_34),
.B2(n_33),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_128),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_34),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_130),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_107),
.B(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_138),
.B(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_134),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_136),
.B1(n_139),
.B2(n_74),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_79),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_96),
.A2(n_90),
.B1(n_70),
.B2(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_90),
.B1(n_70),
.B2(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_113),
.C(n_95),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_137),
.C(n_127),
.Y(n_173)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_150),
.B1(n_155),
.B2(n_161),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_95),
.B1(n_92),
.B2(n_114),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_110),
.B(n_106),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_106),
.B(n_107),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_116),
.B1(n_75),
.B2(n_31),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_33),
.A3(n_27),
.B1(n_34),
.B2(n_17),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_17),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_165),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_70),
.B1(n_66),
.B2(n_89),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_116),
.B1(n_89),
.B2(n_33),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_164),
.B(n_74),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_31),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_74),
.B1(n_27),
.B2(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_33),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_120),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_172),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_124),
.C(n_119),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_188),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_124),
.C(n_120),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_129),
.B(n_117),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_182),
.B(n_154),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_129),
.B(n_136),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

AO22x2_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_122),
.B1(n_132),
.B2(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_157),
.B1(n_146),
.B2(n_148),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_135),
.CI(n_143),
.CON(n_188),
.SN(n_188)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_166),
.B1(n_150),
.B2(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_74),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_167),
.B1(n_170),
.B2(n_166),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_27),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_148),
.B(n_8),
.Y(n_198)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

AO21x1_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_192),
.B(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_191),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_207),
.B1(n_210),
.B2(n_213),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_219),
.B1(n_221),
.B2(n_185),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_149),
.B1(n_160),
.B2(n_156),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_160),
.B1(n_171),
.B2(n_165),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_8),
.B(n_15),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_220),
.B(n_10),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_74),
.B1(n_27),
.B2(n_2),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_15),
.C(n_14),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_177),
.C(n_184),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_15),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_189),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_174),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_0),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_179),
.B(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_174),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_223),
.B1(n_232),
.B2(n_239),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_216),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_210),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_176),
.C(n_184),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_236),
.C(n_238),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_182),
.C(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_190),
.C(n_188),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_183),
.B1(n_190),
.B2(n_181),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_183),
.B1(n_188),
.B2(n_6),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_220),
.B1(n_221),
.B2(n_219),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_250),
.C(n_252),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_249),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_213),
.B1(n_207),
.B2(n_247),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_211),
.Y(n_250)
);

FAx1_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_227),
.CI(n_238),
.CON(n_255),
.SN(n_255)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_260),
.B(n_263),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_237),
.B(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_236),
.B(n_233),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_264),
.B(n_243),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_228),
.B(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_229),
.C(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_262),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_205),
.B(n_212),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_226),
.C(n_229),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_214),
.C(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_259),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_248),
.B1(n_245),
.B2(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_276),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_8),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_9),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_9),
.B(n_11),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_10),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_264),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_4),
.B(n_6),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_11),
.B1(n_12),
.B2(n_6),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_271),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_267),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_287),
.B(n_288),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_271),
.C(n_12),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_286),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_4),
.B(n_7),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_280),
.B(n_281),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_289),
.C(n_291),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_4),
.B(n_7),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_7),
.Y(n_296)
);


endmodule