module real_jpeg_29261_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_0),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_107),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_0),
.A2(n_53),
.B1(n_54),
.B2(n_107),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_0),
.A2(n_58),
.B1(n_60),
.B2(n_107),
.Y(n_241)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_1),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_1),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_27),
.B1(n_31),
.B2(n_37),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_37),
.B1(n_58),
.B2(n_60),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_3),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_25),
.B1(n_58),
.B2(n_60),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_5),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_48),
.B1(n_58),
.B2(n_60),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_48),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_7),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_7),
.A2(n_27),
.B1(n_31),
.B2(n_168),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_7),
.A2(n_53),
.B1(n_54),
.B2(n_168),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_7),
.A2(n_58),
.B1(n_60),
.B2(n_168),
.Y(n_254)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_9),
.B(n_26),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_9),
.B(n_31),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_9),
.A2(n_31),
.B(n_206),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_166),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_55),
.B(n_58),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_75),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_9),
.A2(n_92),
.B1(n_111),
.B2(n_254),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_10),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_27),
.B1(n_31),
.B2(n_46),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_10),
.A2(n_46),
.B1(n_58),
.B2(n_60),
.Y(n_181)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_12),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_12),
.A2(n_27),
.B1(n_31),
.B2(n_133),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_133),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_12),
.A2(n_58),
.B1(n_60),
.B2(n_133),
.Y(n_246)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_14),
.A2(n_27),
.B1(n_31),
.B2(n_66),
.Y(n_71)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_14),
.Y(n_205)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_15),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_340),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_80),
.B(n_338),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_20),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_21),
.A2(n_44),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_22),
.A2(n_33),
.B(n_79),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_29),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_29),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g165 ( 
.A(n_23),
.B(n_166),
.CON(n_165),
.SN(n_165)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_26),
.A2(n_33),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_27),
.A2(n_34),
.B1(n_165),
.B2(n_179),
.Y(n_178)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_27),
.A2(n_53),
.A3(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_29),
.B(n_31),
.Y(n_179)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_32),
.A2(n_45),
.B(n_49),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_33),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_39),
.B(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_72),
.C(n_77),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_40),
.A2(n_41),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.C(n_63),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_42),
.A2(n_43),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_44),
.A2(n_49),
.B1(n_106),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_44),
.A2(n_49),
.B1(n_132),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_50),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_50),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_50),
.A2(n_63),
.B1(n_306),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_61),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_57),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_99),
.B(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_51),
.A2(n_61),
.B(n_115),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_51),
.A2(n_57),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_51),
.A2(n_139),
.B(n_214),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_51),
.A2(n_57),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_51),
.A2(n_57),
.B1(n_213),
.B2(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_54),
.B(n_204),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_54),
.A2(n_56),
.B(n_166),
.C(n_233),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_98),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_57),
.B(n_166),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_60),
.B(n_259),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_62),
.B(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_63),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_64),
.A2(n_74),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_69),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_65),
.A2(n_70),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_65),
.A2(n_70),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_65),
.A2(n_70),
.B1(n_162),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_65),
.A2(n_70),
.B1(n_190),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_75),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_74),
.A2(n_76),
.B(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_74),
.A2(n_129),
.B(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_77),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_331),
.B(n_337),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_301),
.A3(n_323),
.B1(n_329),
.B2(n_330),
.C(n_342),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_151),
.B(n_300),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_134),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_84),
.B(n_134),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_108),
.C(n_119),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_85),
.A2(n_86),
.B1(n_108),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_100),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_102),
.C(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_97),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_88),
.B(n_97),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_89),
.A2(n_112),
.B(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_90),
.A2(n_96),
.B(n_124),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_90),
.A2(n_91),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_96),
.Y(n_95)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_91),
.Y(n_255)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_92),
.A2(n_111),
.B1(n_122),
.B2(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_112),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_95),
.A2(n_111),
.B(n_241),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_108),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_118),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_110),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_114),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_110),
.A2(n_145),
.B(n_148),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B(n_113),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_111),
.A2(n_246),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_119),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_128),
.C(n_130),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_120),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_125),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_128),
.A2(n_130),
.B1(n_131),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_128),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_149),
.B2(n_150),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_137),
.B(n_144),
.C(n_150),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_140),
.B(n_143),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_142),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_143),
.B(n_303),
.C(n_313),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_143),
.A2(n_303),
.B1(n_304),
.B2(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_143),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_294),
.B(n_299),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_194),
.B(n_280),
.C(n_293),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_182),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_154),
.B(n_182),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_169),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_156),
.B(n_157),
.C(n_169),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_164),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_166),
.B(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_171),
.B(n_175),
.C(n_177),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_183),
.A2(n_184),
.B1(n_275),
.B2(n_277),
.Y(n_274)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_188),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_193),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_193),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_279),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_272),
.B(n_278),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_224),
.B(n_271),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_215),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_198),
.B(n_215),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_208),
.C(n_211),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_199),
.A2(n_200),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_222),
.C(n_223),
.Y(n_273)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_265),
.B(n_270),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_242),
.B(n_264),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_227),
.B(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_232),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_241),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_250),
.B(n_263),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_248),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_256),
.B(n_262),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_273),
.B(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_282),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_291),
.B2(n_292),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_288),
.C(n_292),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_315),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_310),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_312),
.B1(n_317),
.B2(n_321),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_321),
.C(n_322),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_314),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_322),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_334),
.Y(n_336)
);


endmodule