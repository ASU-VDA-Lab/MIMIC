module real_jpeg_32769_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_57;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_50;
wire n_33;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_58;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_59;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_SL g59 ( 
.A(n_0),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_2),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx2_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

NAND2x1p5_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_10),
.Y(n_9)
);

AND2x4_ASAP7_75t_SL g21 ( 
.A(n_4),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_4),
.B(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_6),
.A2(n_7),
.B1(n_12),
.B2(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_18),
.Y(n_49)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_19),
.B1(n_32),
.B2(n_34),
.C(n_41),
.Y(n_8)
);

AO21x1_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_13),
.B(n_17),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_45),
.Y(n_44)
);

OA21x2_ASAP7_75t_L g48 ( 
.A1(n_12),
.A2(n_49),
.B(n_50),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_45),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_28),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_35),
.B(n_38),
.Y(n_34)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_31),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

AOI211xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_46),
.C(n_55),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_45),
.B(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_48),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);


endmodule