module fake_netlist_1_9987_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g12 ( .A(n_10), .B(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_3), .B(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_11), .A2(n_7), .B1(n_1), .B2(n_2), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_14), .B(n_0), .Y(n_18) );
OAI22xp5_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_19) );
BUFx4f_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
OAI22xp33_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_17), .B1(n_16), .B2(n_13), .Y(n_22) );
OAI21x1_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_12), .B(n_14), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_20), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_22), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_17), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AOI21xp33_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_18), .B(n_4), .Y(n_31) );
OAI21xp5_ASAP7_75t_L g32 ( .A1(n_28), .A2(n_24), .B(n_20), .Y(n_32) );
AND2x4_ASAP7_75t_L g33 ( .A(n_30), .B(n_24), .Y(n_33) );
A2O1A1Ixp33_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_15), .B(n_24), .C(n_12), .Y(n_34) );
OAI311xp33_ASAP7_75t_L g35 ( .A1(n_30), .A2(n_15), .A3(n_24), .B1(n_4), .C1(n_6), .Y(n_35) );
AOI22xp33_ASAP7_75t_SL g36 ( .A1(n_33), .A2(n_32), .B1(n_6), .B2(n_8), .Y(n_36) );
BUFx2_ASAP7_75t_L g37 ( .A(n_33), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
AOI22xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_36), .B1(n_35), .B2(n_34), .Y(n_39) );
endmodule