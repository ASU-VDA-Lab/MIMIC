module fake_jpeg_1163_n_452 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_452);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_47),
.Y(n_129)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_50),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_52),
.Y(n_113)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_53),
.Y(n_150)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_65),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_88),
.Y(n_97)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_21),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_15),
.B(n_9),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_83),
.Y(n_109)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_15),
.B(n_9),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_90),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_9),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_95),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_94),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_102),
.A2(n_103),
.B1(n_124),
.B2(n_133),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_42),
.B1(n_21),
.B2(n_43),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_32),
.B1(n_25),
.B2(n_27),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_134),
.B1(n_141),
.B2(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_39),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_112),
.B(n_119),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_39),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_52),
.A2(n_42),
.B1(n_43),
.B2(n_41),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_41),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_136),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_34),
.B1(n_38),
.B2(n_29),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_71),
.A2(n_34),
.B1(n_38),
.B2(n_29),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_30),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_27),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_42),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_72),
.A2(n_76),
.B1(n_49),
.B2(n_45),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_46),
.A2(n_25),
.B1(n_19),
.B2(n_42),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_167),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_115),
.B1(n_110),
.B2(n_125),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_154),
.A2(n_145),
.B(n_99),
.C(n_104),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_157),
.Y(n_196)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_160),
.Y(n_207)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_114),
.Y(n_161)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_120),
.A2(n_42),
.B1(n_70),
.B2(n_67),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_168),
.B1(n_180),
.B2(n_183),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_97),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_163),
.B(n_177),
.Y(n_202)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_57),
.B1(n_50),
.B2(n_19),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_113),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_174),
.Y(n_205)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_176),
.Y(n_209)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_108),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_179),
.Y(n_211)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_53),
.B1(n_93),
.B2(n_24),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_182),
.Y(n_217)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_109),
.B(n_0),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_189),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_116),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_194),
.B1(n_145),
.B2(n_123),
.Y(n_213)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_137),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_103),
.B(n_24),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_142),
.C(n_133),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_123),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_193),
.B(n_132),
.CI(n_124),
.CON(n_195),
.SN(n_195)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_195),
.B(n_99),
.Y(n_250)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_98),
.B1(n_150),
.B2(n_131),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_215),
.B1(n_219),
.B2(n_220),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_206),
.B(n_157),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_152),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_153),
.A2(n_150),
.B1(n_98),
.B2(n_131),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_153),
.A2(n_137),
.B1(n_130),
.B2(n_147),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_130),
.B1(n_151),
.B2(n_128),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_106),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_165),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_180),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_154),
.A2(n_122),
.B1(n_151),
.B2(n_128),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_177),
.B1(n_183),
.B2(n_166),
.Y(n_243)
);

NAND2x1_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_171),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_236),
.B(n_247),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_167),
.C(n_177),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_235),
.C(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_251),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_206),
.C(n_201),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_237),
.A2(n_226),
.B1(n_196),
.B2(n_217),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_161),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_241),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_218),
.B1(n_217),
.B2(n_205),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_176),
.C(n_178),
.Y(n_244)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_250),
.C(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_164),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_195),
.B(n_158),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_159),
.C(n_170),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_227),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_196),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_251),
.A2(n_204),
.B1(n_215),
.B2(n_219),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_256),
.A2(n_260),
.B1(n_266),
.B2(n_272),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_223),
.B(n_198),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_258),
.A2(n_271),
.B(n_278),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_198),
.B1(n_202),
.B2(n_220),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_234),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_264),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_244),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_228),
.A2(n_213),
.B(n_224),
.Y(n_271)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_218),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_268),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_247),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_235),
.C(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_290),
.C(n_275),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_232),
.B(n_228),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_285),
.A2(n_259),
.B1(n_277),
.B2(n_271),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_292),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_287),
.B(n_265),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_231),
.C(n_242),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_269),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_301),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_297),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_233),
.B(n_237),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_302),
.A2(n_243),
.B(n_255),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_252),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_278),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_310),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_315),
.C(n_320),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_265),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_311),
.B(n_312),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_262),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_260),
.C(n_258),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_324),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_266),
.C(n_269),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_256),
.B1(n_229),
.B2(n_272),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_291),
.B1(n_280),
.B2(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_323),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_286),
.B(n_207),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_288),
.B(n_207),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_325),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_237),
.C(n_255),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_294),
.C(n_283),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_296),
.B(n_292),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_200),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_253),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_314),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_333),
.B(n_345),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_337),
.B(n_347),
.Y(n_357)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_316),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_354),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_296),
.B(n_302),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_338),
.A2(n_346),
.B1(n_348),
.B2(n_349),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_321),
.A2(n_280),
.B1(n_282),
.B2(n_295),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_341),
.A2(n_351),
.B1(n_274),
.B2(n_225),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_353),
.Y(n_358)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_299),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_305),
.A2(n_281),
.B1(n_297),
.B2(n_293),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_267),
.B(n_230),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_293),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_350),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_319),
.A2(n_229),
.B1(n_293),
.B2(n_267),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_226),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_312),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_371),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_326),
.C(n_311),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_364),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_334),
.A2(n_323),
.B1(n_307),
.B2(n_320),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_361),
.A2(n_344),
.B1(n_345),
.B2(n_349),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_343),
.A2(n_329),
.B1(n_315),
.B2(n_330),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_363),
.A2(n_367),
.B1(n_351),
.B2(n_354),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_340),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_310),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_370),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_333),
.A2(n_317),
.B1(n_322),
.B2(n_328),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_339),
.A2(n_317),
.B(n_208),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_373),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_203),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_203),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_372),
.A2(n_334),
.B1(n_350),
.B2(n_347),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_210),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_212),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_210),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_212),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_348),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_378),
.A2(n_394),
.B1(n_372),
.B2(n_361),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_367),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_379),
.B(n_383),
.Y(n_411)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_381),
.A2(n_388),
.B1(n_395),
.B2(n_357),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_358),
.C(n_370),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_368),
.Y(n_384)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_384),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_353),
.C(n_335),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_386),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_337),
.C(n_341),
.Y(n_386)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_216),
.C(n_224),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_371),
.C(n_356),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_393),
.B(n_363),
.Y(n_399)
);

INVx11_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_208),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_357),
.C(n_366),
.Y(n_407)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_387),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_397),
.B(n_402),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_399),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_404),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_365),
.Y(n_402)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_378),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_406),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_392),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_216),
.C(n_224),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_408),
.B(n_412),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_389),
.A2(n_200),
.B(n_169),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_409),
.A2(n_391),
.B(n_214),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_214),
.C(n_104),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_385),
.C(n_390),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_416),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_403),
.C(n_401),
.Y(n_416)
);

XOR2x2_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_386),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_417),
.A2(n_424),
.B(n_10),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_392),
.C(n_381),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_412),
.C(n_214),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_422),
.A2(n_10),
.B(n_3),
.Y(n_435)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_398),
.A2(n_394),
.B(n_396),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_393),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_425),
.B(n_11),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_428),
.B(n_429),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_122),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_430),
.B(n_431),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_155),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_435),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_421),
.A2(n_155),
.B1(n_3),
.B2(n_4),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_433),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_415),
.B(n_420),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_426),
.A2(n_413),
.B(n_418),
.Y(n_437)
);

AO21x1_ASAP7_75t_L g444 ( 
.A1(n_437),
.A2(n_433),
.B(n_428),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_414),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_442),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_417),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_444),
.C(n_446),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_11),
.Y(n_446)
);

AOI321xp33_ASAP7_75t_L g447 ( 
.A1(n_445),
.A2(n_441),
.A3(n_436),
.B1(n_6),
.B2(n_10),
.C(n_11),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_447),
.A2(n_4),
.B1(n_12),
.B2(n_13),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_SL g450 ( 
.A(n_449),
.B(n_448),
.C(n_4),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_14),
.B(n_0),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_14),
.C(n_0),
.Y(n_452)
);


endmodule