module fake_jpeg_15743_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_52),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_1),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_85),
.Y(n_107)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_64),
.B(n_46),
.C(n_53),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_92),
.B(n_59),
.C(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_59),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_97),
.Y(n_119)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_63),
.B1(n_56),
.B2(n_51),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_63),
.B1(n_56),
.B2(n_61),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_108),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_54),
.B1(n_55),
.B2(n_43),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_105),
.B1(n_110),
.B2(n_112),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_60),
.B1(n_45),
.B2(n_43),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_45),
.B1(n_62),
.B2(n_22),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_107),
.C(n_110),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_113),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_117),
.B1(n_5),
.B2(n_6),
.Y(n_129)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_105),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_93),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_137),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_102),
.B1(n_94),
.B2(n_104),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_124),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_140),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_132),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_134),
.B(n_126),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_144),
.B(n_146),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_134),
.B(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_127),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_138),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_7),
.B(n_8),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_145),
.A2(n_127),
.B1(n_121),
.B2(n_123),
.Y(n_151)
);

AOI22x1_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_122),
.B1(n_131),
.B2(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_154),
.Y(n_156)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_155),
.B1(n_115),
.B2(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_151),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_148),
.B(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_118),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_7),
.B(n_8),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_10),
.B(n_11),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_29),
.B1(n_40),
.B2(n_39),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_42),
.B(n_25),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_19),
.C(n_37),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_38),
.B1(n_18),
.B2(n_27),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_17),
.B(n_36),
.Y(n_169)
);


endmodule