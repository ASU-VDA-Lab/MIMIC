module fake_ariane_1080_n_1035 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_1035);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1035;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_752;
wire n_1029;
wire n_341;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_586;
wire n_443;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_597;
wire n_269;
wire n_816;
wire n_1018;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_553;
wire n_446;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_485;
wire n_401;
wire n_495;
wire n_267;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_529;
wire n_502;
wire n_561;
wire n_253;
wire n_770;
wire n_839;
wire n_821;
wire n_928;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_612;
wire n_449;
wire n_333;
wire n_388;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_543;
wire n_260;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_262;
wire n_490;
wire n_743;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_527;
wire n_741;
wire n_290;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_673;
wire n_452;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_534;
wire n_249;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_1027;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_580;
wire n_358;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_718;
wire n_329;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_650;
wire n_258;
wire n_364;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_233),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_26),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_87),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_106),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_55),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_96),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_31),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_21),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_76),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_81),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_157),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_166),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_71),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_0),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_3),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_191),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_130),
.Y(n_259)
);

CKINVDCx12_ASAP7_75t_R g260 ( 
.A(n_51),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_117),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_156),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_172),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_73),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_95),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_4),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_153),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_97),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_192),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_80),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_85),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_2),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_147),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_19),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_18),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_24),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_52),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_127),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_18),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_25),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_145),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_88),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_58),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_209),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_115),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_121),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_102),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_222),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_61),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_232),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_177),
.Y(n_296)
);

BUFx2_ASAP7_75t_SL g297 ( 
.A(n_198),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_194),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_202),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_105),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_77),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_215),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_10),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_1),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_112),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_190),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_143),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_37),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_69),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_75),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_3),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_184),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_201),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_56),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_23),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_163),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_142),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_220),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_134),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_53),
.Y(n_322)
);

BUFx8_ASAP7_75t_SL g323 ( 
.A(n_152),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_64),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_182),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_148),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_47),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_99),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_181),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_70),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_216),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_160),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_155),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_193),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_37),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_33),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_224),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_5),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_27),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_54),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_150),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_90),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_33),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_227),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_137),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_189),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_125),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_98),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_42),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_151),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_113),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_44),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_200),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_180),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_135),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_93),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_161),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_84),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_1),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_9),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_40),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_83),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_176),
.B(n_230),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_183),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_178),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_168),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_179),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_57),
.Y(n_369)
);

HB1xp67_ASAP7_75t_SL g370 ( 
.A(n_221),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_27),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_207),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_154),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_146),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_111),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_32),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_5),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_10),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_219),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_79),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_103),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_185),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_228),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_11),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_229),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_167),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_223),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_158),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_173),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_144),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_86),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_138),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_15),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_199),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_128),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_238),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_323),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_247),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_245),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_243),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_238),
.B(n_2),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_284),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_348),
.B(n_4),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_243),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_236),
.A2(n_246),
.B(n_242),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_298),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_292),
.B(n_45),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_251),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_263),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_248),
.A2(n_6),
.B(n_7),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_310),
.B(n_8),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_310),
.B(n_9),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_11),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_247),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_255),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_244),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_263),
.Y(n_421)
);

BUFx12f_ASAP7_75t_L g422 ( 
.A(n_294),
.Y(n_422)
);

OAI22x1_ASAP7_75t_SL g423 ( 
.A1(n_235),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_247),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_276),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_256),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_285),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_330),
.B(n_46),
.Y(n_428)
);

AOI22x1_ASAP7_75t_SL g429 ( 
.A1(n_268),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_313),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_317),
.B(n_16),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_294),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_340),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_361),
.B(n_16),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_20),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_307),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_283),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_20),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_266),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_307),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_247),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_254),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_250),
.B(n_21),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_258),
.B(n_22),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_254),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_254),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_317),
.B(n_22),
.Y(n_448)
);

CKINVDCx11_ASAP7_75t_R g449 ( 
.A(n_274),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_254),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_262),
.B(n_23),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_261),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_261),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_261),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_384),
.B(n_24),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_308),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_261),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_288),
.B(n_25),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_332),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_264),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_289),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_270),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_374),
.B(n_26),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_324),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_289),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_386),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_272),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_289),
.B(n_48),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_289),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_271),
.B(n_28),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_299),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_279),
.B(n_28),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_277),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_299),
.Y(n_475)
);

NOR2x1_ASAP7_75t_L g476 ( 
.A(n_280),
.B(n_50),
.Y(n_476)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_366),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_299),
.Y(n_478)
);

BUFx8_ASAP7_75t_SL g479 ( 
.A(n_304),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_299),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_328),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_345),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_319),
.Y(n_483)
);

BUFx12f_ASAP7_75t_L g484 ( 
.A(n_366),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_278),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_319),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_281),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_293),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_282),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_295),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_302),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_303),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_306),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_305),
.Y(n_494)
);

BUFx8_ASAP7_75t_SL g495 ( 
.A(n_339),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_316),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_321),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_309),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_393),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_331),
.A2(n_60),
.B(n_59),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g501 ( 
.A1(n_327),
.A2(n_35),
.B(n_36),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_252),
.B(n_62),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_370),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_344),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_346),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g506 ( 
.A(n_311),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_347),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_354),
.B(n_38),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_355),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_356),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_357),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_335),
.B(n_39),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_275),
.B(n_41),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_336),
.Y(n_514)
);

BUFx12f_ASAP7_75t_L g515 ( 
.A(n_343),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_318),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_320),
.A2(n_42),
.B1(n_43),
.B2(n_63),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_234),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_359),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_362),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_363),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_365),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_371),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_367),
.A2(n_43),
.B(n_65),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_376),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_368),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_379),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_397),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_405),
.B(n_395),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_430),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_518),
.B(n_381),
.Y(n_533)
);

AND3x2_ASAP7_75t_L g534 ( 
.A(n_409),
.B(n_372),
.C(n_337),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_492),
.B(n_394),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_438),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_481),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_420),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_479),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_495),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_434),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_449),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_520),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_425),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_485),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_401),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_408),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_506),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_398),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_398),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_418),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_515),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_422),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_426),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_484),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_518),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_424),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_428),
.A2(n_404),
.B1(n_402),
.B2(n_396),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_478),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_421),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_433),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_411),
.B(n_389),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_437),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_459),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_519),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_519),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_411),
.B(n_390),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_478),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_411),
.B(n_382),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_R g572 ( 
.A(n_487),
.B(n_489),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_456),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_410),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_419),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_477),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_494),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_477),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_498),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_507),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_511),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_514),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_523),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_482),
.B(n_237),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_504),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_505),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_441),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_516),
.B(n_391),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_516),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_396),
.B(n_267),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_464),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_400),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_465),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_404),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_407),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_467),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_424),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_511),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_509),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_442),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_510),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_431),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_448),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_407),
.B(n_312),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_592),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_598),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_545),
.Y(n_608)
);

NOR3xp33_ASAP7_75t_L g609 ( 
.A(n_595),
.B(n_463),
.C(n_451),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_586),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_545),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_535),
.B(n_471),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_531),
.Y(n_613)
);

NOR2xp67_ASAP7_75t_L g614 ( 
.A(n_528),
.B(n_427),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_561),
.B(n_471),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_561),
.B(n_513),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_587),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_537),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_570),
.B(n_513),
.Y(n_619)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_591),
.B(n_414),
.C(n_412),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_570),
.B(n_557),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_605),
.B(n_415),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_567),
.B(n_412),
.Y(n_623)
);

BUFx5_ASAP7_75t_L g624 ( 
.A(n_532),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_577),
.B(n_445),
.C(n_444),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_533),
.B(n_415),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_534),
.B(n_416),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_562),
.B(n_458),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_560),
.B(n_493),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_548),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_550),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_588),
.B(n_414),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_544),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_529),
.B(n_403),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_563),
.B(n_565),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_603),
.A2(n_512),
.B1(n_517),
.B2(n_503),
.Y(n_636)
);

AOI221xp5_ASAP7_75t_L g637 ( 
.A1(n_596),
.A2(n_435),
.B1(n_417),
.B2(n_439),
.C(n_436),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_530),
.A2(n_508),
.B(n_473),
.C(n_439),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_555),
.B(n_522),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_550),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_547),
.B(n_496),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_582),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_529),
.B(n_497),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_566),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_550),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_568),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_550),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_539),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_594),
.B(n_597),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_589),
.B(n_460),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_572),
.B(n_462),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_546),
.B(n_502),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_552),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_571),
.B(n_462),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_604),
.A2(n_455),
.B1(n_436),
.B2(n_417),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_581),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_600),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_602),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_580),
.Y(n_660)
);

BUFx5_ASAP7_75t_L g661 ( 
.A(n_552),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_542),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_551),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_573),
.B(n_468),
.Y(n_664)
);

OR2x6_ASAP7_75t_L g665 ( 
.A(n_555),
.B(n_435),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_558),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_559),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_601),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_576),
.B(n_579),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_599),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_552),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_552),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_564),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_569),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_575),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_662),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_632),
.B(n_583),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_622),
.A2(n_584),
.B1(n_575),
.B2(n_499),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_610),
.B(n_574),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_613),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_670),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_660),
.B(n_549),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_626),
.B(n_488),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_607),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_649),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_SL g686 ( 
.A(n_637),
.B(n_543),
.C(n_593),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_617),
.B(n_553),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_618),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_638),
.A2(n_525),
.B1(n_490),
.B2(n_491),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_630),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_642),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_607),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_645),
.B(n_536),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_644),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_651),
.B(n_488),
.Y(n_695)
);

CKINVDCx8_ASAP7_75t_R g696 ( 
.A(n_634),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_623),
.Y(n_697)
);

NOR2x1p5_ASAP7_75t_L g698 ( 
.A(n_633),
.B(n_540),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_652),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_656),
.A2(n_585),
.B1(n_406),
.B2(n_526),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_631),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_625),
.A2(n_578),
.B1(n_297),
.B2(n_476),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_608),
.B(n_590),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_631),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_657),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_614),
.B(n_554),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_612),
.B(n_538),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_640),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_636),
.A2(n_240),
.B1(n_241),
.B2(n_239),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_658),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_659),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_650),
.B(n_556),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_611),
.B(n_521),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_615),
.A2(n_500),
.B(n_524),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_640),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_634),
.B(n_521),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_606),
.B(n_526),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_621),
.B(n_527),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_616),
.B(n_619),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_R g720 ( 
.A(n_647),
.B(n_541),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_629),
.B(n_527),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_R g722 ( 
.A(n_669),
.B(n_260),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_635),
.B(n_413),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_639),
.B(n_364),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_624),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_666),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_665),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_675),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_655),
.B(n_624),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_624),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_624),
.B(n_249),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_628),
.B(n_423),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_640),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_620),
.A2(n_501),
.B1(n_429),
.B2(n_524),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_667),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_663),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_668),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_609),
.B(n_469),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_627),
.B(n_253),
.Y(n_739)
);

BUFx12f_ASAP7_75t_L g740 ( 
.A(n_646),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_643),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_671),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_664),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_672),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_641),
.A2(n_259),
.B1(n_265),
.B2(n_257),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_646),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_646),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_653),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_SL g749 ( 
.A1(n_689),
.A2(n_674),
.B(n_673),
.C(n_661),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_680),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_677),
.B(n_648),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_729),
.A2(n_273),
.B(n_269),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_719),
.B(n_661),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_743),
.B(n_748),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_676),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_700),
.A2(n_734),
.B1(n_724),
.B2(n_741),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_709),
.A2(n_287),
.B(n_290),
.C(n_286),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_731),
.A2(n_296),
.B(n_291),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_740),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_SL g760 ( 
.A(n_681),
.B(n_648),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_693),
.B(n_648),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_683),
.B(n_654),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_695),
.B(n_654),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_688),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_725),
.A2(n_730),
.B(n_718),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_682),
.B(n_654),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_714),
.A2(n_469),
.B(n_300),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_733),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_715),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_SL g770 ( 
.A(n_726),
.B(n_301),
.Y(n_770)
);

CKINVDCx14_ASAP7_75t_R g771 ( 
.A(n_720),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_716),
.B(n_443),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_716),
.B(n_443),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_728),
.B(n_446),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_696),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_699),
.B(n_721),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_710),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_690),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_712),
.A2(n_360),
.B(n_314),
.C(n_315),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_727),
.B(n_322),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_702),
.A2(n_678),
.B(n_738),
.C(n_705),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_707),
.Y(n_782)
);

BUFx6f_ASAP7_75t_SL g783 ( 
.A(n_697),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_738),
.A2(n_369),
.B(n_326),
.C(n_329),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_703),
.B(n_325),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_747),
.B(n_333),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_711),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_R g788 ( 
.A(n_686),
.B(n_334),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

AOI21x1_ASAP7_75t_L g790 ( 
.A1(n_742),
.A2(n_486),
.B(n_447),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_733),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_685),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_745),
.A2(n_388),
.B1(n_341),
.B2(n_342),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_691),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_713),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_698),
.B(n_446),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_717),
.Y(n_797)
);

AOI221xp5_ASAP7_75t_L g798 ( 
.A1(n_732),
.A2(n_350),
.B1(n_351),
.B2(n_353),
.C(n_358),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_684),
.Y(n_799)
);

AOI21x1_ASAP7_75t_L g800 ( 
.A1(n_744),
.A2(n_486),
.B(n_450),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_SL g801 ( 
.A(n_722),
.B(n_375),
.C(n_373),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_739),
.A2(n_385),
.B(n_380),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_724),
.B(n_392),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_701),
.B(n_447),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_694),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_797),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_754),
.B(n_679),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_768),
.Y(n_808)
);

AO21x2_ASAP7_75t_L g809 ( 
.A1(n_767),
.A2(n_735),
.B(n_736),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_749),
.A2(n_723),
.B(n_737),
.Y(n_810)
);

OAI21x1_ASAP7_75t_L g811 ( 
.A1(n_765),
.A2(n_692),
.B(n_706),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_768),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_759),
.B(n_687),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_768),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_750),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_791),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_790),
.A2(n_708),
.B(n_704),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_778),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_777),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_763),
.A2(n_708),
.B(n_704),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_791),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_800),
.A2(n_708),
.B(n_704),
.Y(n_822)
);

AO21x2_ASAP7_75t_L g823 ( 
.A1(n_753),
.A2(n_746),
.B(n_452),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_791),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_762),
.A2(n_72),
.B(n_74),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_787),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_775),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_792),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_782),
.B(n_450),
.Y(n_829)
);

AO21x2_ASAP7_75t_L g830 ( 
.A1(n_781),
.A2(n_483),
.B(n_480),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_769),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_789),
.Y(n_832)
);

AO21x2_ASAP7_75t_L g833 ( 
.A1(n_752),
.A2(n_480),
.B(n_475),
.Y(n_833)
);

BUFx4f_ASAP7_75t_L g834 ( 
.A(n_766),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_799),
.Y(n_835)
);

INVx3_ASAP7_75t_SL g836 ( 
.A(n_796),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_764),
.Y(n_837)
);

AO21x2_ASAP7_75t_L g838 ( 
.A1(n_795),
.A2(n_475),
.B(n_472),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_774),
.B(n_772),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_776),
.B(n_453),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_789),
.A2(n_78),
.B(n_82),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_773),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_758),
.A2(n_89),
.B(n_91),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_755),
.Y(n_844)
);

AO21x2_ASAP7_75t_L g845 ( 
.A1(n_784),
.A2(n_472),
.B(n_470),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_794),
.Y(n_846)
);

AOI22x1_ASAP7_75t_L g847 ( 
.A1(n_802),
.A2(n_470),
.B1(n_466),
.B2(n_461),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_805),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_796),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_804),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_756),
.A2(n_92),
.B(n_94),
.Y(n_851)
);

AO21x2_ASAP7_75t_L g852 ( 
.A1(n_785),
.A2(n_466),
.B(n_461),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_761),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_760),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_803),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_751),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_815),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_810),
.A2(n_757),
.B(n_779),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_828),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_856),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_818),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_844),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_834),
.B(n_770),
.Y(n_863)
);

INVx6_ASAP7_75t_L g864 ( 
.A(n_835),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_807),
.B(n_771),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_819),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_848),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_855),
.A2(n_788),
.B1(n_798),
.B2(n_801),
.Y(n_868)
);

BUFx2_ASAP7_75t_R g869 ( 
.A(n_836),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_826),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_827),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_855),
.A2(n_786),
.B1(n_780),
.B2(n_793),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_839),
.A2(n_783),
.B1(n_457),
.B2(n_454),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_834),
.B(n_783),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_837),
.B(n_832),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_853),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_806),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_854),
.A2(n_457),
.B1(n_454),
.B2(n_101),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_846),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_812),
.Y(n_880)
);

AO21x1_ASAP7_75t_L g881 ( 
.A1(n_851),
.A2(n_100),
.B(n_104),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_850),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_842),
.B(n_226),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_811),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_838),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_829),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_SL g887 ( 
.A1(n_851),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_887)
);

OAI22xp33_ASAP7_75t_L g888 ( 
.A1(n_849),
.A2(n_110),
.B1(n_114),
.B2(n_116),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_838),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_825),
.A2(n_118),
.B(n_119),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_813),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_832),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_840),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_813),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_832),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_862),
.B(n_840),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_874),
.B(n_891),
.Y(n_897)
);

OR2x6_ASAP7_75t_L g898 ( 
.A(n_874),
.B(n_808),
.Y(n_898)
);

NOR2x1_ASAP7_75t_SL g899 ( 
.A(n_877),
.B(n_830),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_894),
.B(n_814),
.Y(n_900)
);

NAND2xp33_ASAP7_75t_R g901 ( 
.A(n_865),
.B(n_816),
.Y(n_901)
);

BUFx8_ASAP7_75t_L g902 ( 
.A(n_871),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_857),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_859),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_860),
.B(n_821),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_861),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_868),
.B(n_847),
.C(n_824),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_R g908 ( 
.A(n_864),
.B(n_821),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_867),
.B(n_812),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_880),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_L g911 ( 
.A(n_863),
.B(n_831),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_R g912 ( 
.A(n_883),
.B(n_841),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_869),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_886),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_880),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_876),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_875),
.B(n_809),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_875),
.B(n_830),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_866),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_870),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_873),
.B(n_872),
.Y(n_921)
);

AOI21xp33_ASAP7_75t_L g922 ( 
.A1(n_858),
.A2(n_845),
.B(n_852),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_882),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_872),
.B(n_820),
.Y(n_924)
);

AO31x2_ASAP7_75t_L g925 ( 
.A1(n_885),
.A2(n_823),
.A3(n_833),
.B(n_843),
.Y(n_925)
);

NAND2x1_ASAP7_75t_L g926 ( 
.A(n_892),
.B(n_895),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_916),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_924),
.B(n_879),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_917),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_903),
.Y(n_930)
);

AND2x2_ASAP7_75t_SL g931 ( 
.A(n_921),
.B(n_893),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_918),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_923),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_906),
.B(n_884),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_905),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_926),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_904),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_920),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_914),
.A2(n_893),
.B1(n_888),
.B2(n_887),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_915),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_919),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_909),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_896),
.B(n_889),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_925),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_910),
.B(n_887),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_899),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_900),
.B(n_878),
.Y(n_947)
);

AO21x2_ASAP7_75t_L g948 ( 
.A1(n_922),
.A2(n_881),
.B(n_890),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_900),
.B(n_817),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_897),
.B(n_817),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_911),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_913),
.B(n_822),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_898),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_902),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_897),
.B(n_822),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_898),
.Y(n_956)
);

OA211x2_ASAP7_75t_L g957 ( 
.A1(n_947),
.A2(n_907),
.B(n_912),
.C(n_901),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_928),
.B(n_908),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_933),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_942),
.B(n_935),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_933),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_937),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_927),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_941),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_930),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_934),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_932),
.B(n_929),
.Y(n_967)
);

OAI21xp33_ASAP7_75t_L g968 ( 
.A1(n_939),
.A2(n_129),
.B(n_131),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_929),
.B(n_132),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_952),
.B(n_133),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_SL g971 ( 
.A(n_931),
.B(n_136),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_SL g972 ( 
.A(n_945),
.B(n_139),
.C(n_140),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_943),
.B(n_141),
.Y(n_973)
);

NAND2x1_ASAP7_75t_L g974 ( 
.A(n_936),
.B(n_946),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_953),
.B(n_149),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_938),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_974),
.Y(n_977)
);

AND3x2_ASAP7_75t_L g978 ( 
.A(n_971),
.B(n_950),
.C(n_951),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_960),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_959),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_966),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_963),
.Y(n_982)
);

NOR2xp67_ASAP7_75t_L g983 ( 
.A(n_967),
.B(n_954),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_965),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_958),
.B(n_940),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_958),
.B(n_940),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_976),
.B(n_936),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_961),
.B(n_949),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_971),
.B(n_969),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_989),
.A2(n_968),
.B1(n_972),
.B2(n_957),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_983),
.B(n_970),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_981),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_980),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_977),
.B(n_975),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_979),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_982),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_984),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_997),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_990),
.A2(n_987),
.B(n_977),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_995),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_997),
.Y(n_1001)
);

OAI31xp33_ASAP7_75t_SL g1002 ( 
.A1(n_991),
.A2(n_978),
.A3(n_986),
.B(n_985),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_993),
.Y(n_1003)
);

OAI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_994),
.A2(n_955),
.B1(n_988),
.B2(n_973),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_998),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_999),
.Y(n_1006)
);

OAI211xp5_ASAP7_75t_SL g1007 ( 
.A1(n_1000),
.A2(n_992),
.B(n_996),
.C(n_956),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_1001),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1003),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_SL g1010 ( 
.A1(n_1002),
.A2(n_1004),
.B(n_950),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_998),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_1005),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_1010),
.B(n_948),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1008),
.Y(n_1014)
);

AOI221xp5_ASAP7_75t_L g1015 ( 
.A1(n_1006),
.A2(n_948),
.B1(n_944),
.B2(n_964),
.C(n_962),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1009),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1012),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_1014),
.B(n_1011),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1016),
.Y(n_1019)
);

O2A1O1Ixp5_ASAP7_75t_L g1020 ( 
.A1(n_1017),
.A2(n_1013),
.B(n_1015),
.C(n_1007),
.Y(n_1020)
);

AOI221xp5_ASAP7_75t_L g1021 ( 
.A1(n_1019),
.A2(n_159),
.B1(n_165),
.B2(n_169),
.C(n_170),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_SL g1022 ( 
.A1(n_1018),
.A2(n_171),
.B(n_174),
.C(n_175),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1020),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_1022),
.B(n_187),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_SL g1025 ( 
.A(n_1023),
.B(n_1021),
.C(n_188),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1025),
.B(n_1024),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1026),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_1027),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_1028),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1029),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_1030),
.Y(n_1031)
);

AOI222xp33_ASAP7_75t_L g1032 ( 
.A1(n_1031),
.A2(n_195),
.B1(n_197),
.B2(n_203),
.C1(n_204),
.C2(n_205),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1031),
.A2(n_206),
.B1(n_208),
.B2(n_210),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1034),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_1035)
);


endmodule