module real_jpeg_21151_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_40),
.B1(n_55),
.B2(n_76),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_1),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_55),
.Y(n_136)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_26),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_107),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_7),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_91)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_10),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_70),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_80),
.Y(n_123)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_14),
.A2(n_62),
.B(n_84),
.C(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_14),
.B(n_62),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_14),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_14),
.A2(n_15),
.B(n_27),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_15),
.B(n_37),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_15),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_15),
.A2(n_29),
.B1(n_33),
.B2(n_136),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_15),
.B(n_67),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_15),
.A2(n_37),
.B(n_104),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_112),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_20),
.B(n_94),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_71),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_24)
);

OAI21x1_ASAP7_75t_SL g45 ( 
.A1(n_25),
.A2(n_33),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_26),
.B(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_29),
.A2(n_111),
.B1(n_120),
.B2(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_29),
.A2(n_123),
.B(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_30),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_30),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_40),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_36),
.A2(n_40),
.B(n_42),
.C(n_51),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_58),
.Y(n_60)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_38),
.A2(n_62),
.A3(n_66),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_51),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_41),
.CON(n_39),
.SN(n_39)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_41),
.A2(n_63),
.B(n_86),
.C(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_41),
.B(n_85),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_41),
.B(n_111),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.C(n_52),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_52),
.B(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B1(n_67),
.B2(n_68),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_54),
.A2(n_57),
.B1(n_61),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_61),
.B1(n_69),
.B2(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_61)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_58),
.B(n_63),
.Y(n_105)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_93),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_87),
.B(n_90),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_83),
.A2(n_85),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_83),
.A2(n_85),
.B1(n_131),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_83),
.A2(n_85),
.B1(n_100),
.B2(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_102),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_95),
.A2(n_96),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2x2_ASAP7_75t_SL g172 ( 
.A(n_99),
.B(n_102),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_106),
.Y(n_158)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_168),
.B(n_173),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_155),
.B(n_167),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_143),
.B(n_154),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_132),
.B(n_142),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_124),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_128),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_137),
.B(n_141),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_135),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_145),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_157),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_166),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_164),
.C(n_165),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);


endmodule