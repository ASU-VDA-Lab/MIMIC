module fake_ariane_2112_n_2005 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_17, n_225, n_235, n_464, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_384, n_468, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_460, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2005);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2005;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_495;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_489;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1674;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_1913;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_1726;
wire n_1945;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_1003;
wire n_701;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_1063;
wire n_537;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1252;
wire n_1129;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_849;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_174),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_42),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_119),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_263),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_153),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_452),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_223),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_19),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_154),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_136),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_192),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_243),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_367),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_470),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_253),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_378),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_53),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_152),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_271),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_149),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_440),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_376),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_324),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_39),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_319),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_447),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_290),
.Y(n_505)
);

CKINVDCx12_ASAP7_75t_R g506 ( 
.A(n_471),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_39),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_163),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_73),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_353),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_459),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_177),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_312),
.Y(n_513)
);

BUFx5_ASAP7_75t_L g514 ( 
.A(n_59),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_46),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_393),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_221),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_121),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_317),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_261),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_171),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_194),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_436),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_379),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_237),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_472),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_302),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_155),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_242),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_433),
.Y(n_530)
);

BUFx8_ASAP7_75t_SL g531 ( 
.A(n_307),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_448),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_66),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_380),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_390),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_101),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_366),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_309),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_381),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_1),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_188),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_229),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_56),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_451),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_288),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_13),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_159),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_185),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_216),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_158),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_188),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_430),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_399),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_214),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_460),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_46),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_462),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_75),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_245),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_332),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_132),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_435),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_441),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_179),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_211),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_43),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_194),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_323),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_453),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_375),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_365),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_438),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_388),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_153),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_71),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_32),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_8),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_117),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_313),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_29),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_345),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_351),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_233),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_410),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_122),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_230),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_91),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_258),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_252),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_220),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_125),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_343),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_200),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_174),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_374),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_306),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_442),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_125),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_214),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_469),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_465),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_251),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_50),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_12),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_383),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_296),
.Y(n_608)
);

BUFx2_ASAP7_75t_R g609 ( 
.A(n_126),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_184),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_109),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_60),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_456),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_445),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_431),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_110),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_262),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_249),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_444),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_275),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_167),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_168),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_75),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_217),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_432),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_81),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_428),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_33),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_147),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_11),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_454),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_387),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_391),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_389),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_429),
.Y(n_635)
);

BUFx5_ASAP7_75t_L g636 ( 
.A(n_35),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_412),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_301),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_210),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_213),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_449),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_363),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_231),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_356),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_473),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_282),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_372),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_206),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_197),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_239),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_45),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_464),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_285),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_43),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_232),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_419),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_175),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_406),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_164),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_335),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_457),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_298),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_463),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_165),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_316),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_293),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_187),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_170),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_159),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_225),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_334),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_423),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_475),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_156),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_48),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_212),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_292),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_455),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_123),
.Y(n_679)
);

BUFx5_ASAP7_75t_L g680 ( 
.A(n_141),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_318),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_269),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_284),
.Y(n_683)
);

CKINVDCx16_ASAP7_75t_R g684 ( 
.A(n_434),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_0),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_196),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_107),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_398),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_458),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_150),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_217),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_344),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_420),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_109),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_341),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_96),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_310),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_349),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_76),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_417),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_218),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_151),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_439),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_17),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_446),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_183),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_26),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_126),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_260),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_468),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_38),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_474),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_40),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_45),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_179),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_466),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_467),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_498),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_531),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_531),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_600),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_502),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_498),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_540),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_540),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_556),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_564),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_497),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_600),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_629),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_542),
.Y(n_732)
);

INVxp33_ASAP7_75t_SL g733 ( 
.A(n_543),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_629),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_514),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_569),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_514),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_514),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_525),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_563),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_553),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_514),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_514),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_514),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_636),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_517),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_636),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_636),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_636),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_636),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_636),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_680),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_680),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_680),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_591),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_680),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_659),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_680),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_680),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_479),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_621),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_487),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_621),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_517),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_706),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_646),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_488),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_517),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_517),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_658),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_478),
.B(n_0),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_528),
.Y(n_772)
);

INVxp33_ASAP7_75t_L g773 ( 
.A(n_536),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_541),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_684),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_550),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_549),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_706),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_549),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_484),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_551),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_549),
.Y(n_782)
);

CKINVDCx14_ASAP7_75t_R g783 ( 
.A(n_656),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_554),
.Y(n_784)
);

INVxp67_ASAP7_75t_SL g785 ( 
.A(n_549),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_640),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_533),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_483),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_476),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_565),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_576),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_588),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_581),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_589),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_477),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_481),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_547),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_485),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_640),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_596),
.Y(n_800)
);

INVxp33_ASAP7_75t_SL g801 ( 
.A(n_496),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_605),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_640),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_561),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_640),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_611),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_649),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_759),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_759),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_735),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_737),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_738),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_718),
.B(n_480),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_722),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_743),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_744),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_764),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_789),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_745),
.A2(n_486),
.B(n_482),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_733),
.A2(n_588),
.B1(n_631),
.B2(n_617),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_747),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_783),
.B(n_489),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_741),
.B(n_490),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_764),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_748),
.Y(n_826)
);

AND2x2_ASAP7_75t_SL g827 ( 
.A(n_771),
.B(n_578),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_777),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_801),
.B(n_491),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_741),
.B(n_746),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_719),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_773),
.B(n_579),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_733),
.A2(n_714),
.B1(n_495),
.B2(n_687),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_777),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_749),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_782),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_750),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_751),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_752),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_753),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_754),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_782),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_799),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_799),
.Y(n_844)
);

BUFx12f_ASAP7_75t_L g845 ( 
.A(n_720),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_768),
.B(n_516),
.Y(n_846)
);

OA21x2_ASAP7_75t_L g847 ( 
.A1(n_756),
.A2(n_758),
.B(n_803),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_803),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_769),
.B(n_508),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_796),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_779),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_795),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_785),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_786),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_728),
.B(n_656),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_805),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_723),
.B(n_523),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_760),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_762),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_767),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_SL g861 ( 
.A1(n_721),
.A2(n_609),
.B1(n_631),
.B2(n_617),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_724),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_725),
.B(n_726),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_772),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_774),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_776),
.Y(n_866)
);

AND2x2_ASAP7_75t_SL g867 ( 
.A(n_798),
.B(n_578),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_729),
.B(n_524),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_781),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_731),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_858),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_858),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_859),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_827),
.B(n_728),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_847),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_847),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_864),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_821),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_864),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_832),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_827),
.B(n_732),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_847),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_847),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_869),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_SL g885 ( 
.A1(n_821),
.A2(n_730),
.B1(n_761),
.B2(n_721),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_869),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_851),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_851),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_808),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_832),
.B(n_732),
.Y(n_890)
);

NOR2x1_ASAP7_75t_L g891 ( 
.A(n_823),
.B(n_784),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_856),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_808),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_815),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_852),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_856),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_808),
.B(n_672),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_852),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_810),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_810),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_859),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_829),
.A2(n_736),
.B1(n_775),
.B2(n_755),
.Y(n_902)
);

INVx8_ASAP7_75t_L g903 ( 
.A(n_845),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_809),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_852),
.B(n_736),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_811),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_809),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_852),
.B(n_755),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_811),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_812),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_859),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_812),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_827),
.B(n_775),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_814),
.Y(n_914)
);

NAND3xp33_ASAP7_75t_L g915 ( 
.A(n_833),
.B(n_727),
.C(n_757),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_814),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_867),
.A2(n_801),
.B1(n_509),
.B2(n_515),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_859),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_819),
.B(n_850),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_SL g920 ( 
.A1(n_861),
.A2(n_761),
.B1(n_763),
.B2(n_730),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_816),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_816),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_817),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_830),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_831),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_SL g926 ( 
.A1(n_861),
.A2(n_765),
.B1(n_778),
.B2(n_763),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_820),
.A2(n_822),
.B(n_817),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_859),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_867),
.A2(n_518),
.B1(n_521),
.B2(n_507),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_867),
.B(n_788),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_822),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_826),
.B(n_526),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_826),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_SL g934 ( 
.A1(n_845),
.A2(n_778),
.B1(n_765),
.B2(n_780),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_854),
.B(n_734),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_835),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_830),
.Y(n_937)
);

OAI22xp33_ASAP7_75t_SL g938 ( 
.A1(n_813),
.A2(n_792),
.B1(n_855),
.B2(n_740),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_831),
.B(n_739),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_835),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_837),
.A2(n_548),
.B1(n_558),
.B2(n_546),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_SL g942 ( 
.A(n_860),
.B(n_679),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_837),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_838),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_838),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_830),
.A2(n_566),
.B1(n_574),
.B2(n_567),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_839),
.A2(n_623),
.B1(n_690),
.B2(n_592),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_830),
.B(n_790),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_824),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_862),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_839),
.Y(n_951)
);

CKINVDCx11_ASAP7_75t_R g952 ( 
.A(n_863),
.Y(n_952)
);

BUFx6f_ASAP7_75t_SL g953 ( 
.A(n_863),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_860),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_889),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_889),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_903),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_916),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_899),
.B(n_840),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_950),
.B(n_895),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_874),
.A2(n_841),
.B1(n_840),
.B2(n_860),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_900),
.B(n_841),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_916),
.B(n_860),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_880),
.B(n_766),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_925),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_903),
.B(n_863),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_917),
.A2(n_792),
.B1(n_770),
.B2(n_512),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_921),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_L g969 ( 
.A(n_919),
.B(n_616),
.C(n_612),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_903),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_874),
.B(n_853),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_948),
.B(n_863),
.Y(n_972)
);

NAND2x1_ASAP7_75t_L g973 ( 
.A(n_911),
.B(n_860),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_893),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_950),
.B(n_865),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_894),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_881),
.B(n_853),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_890),
.B(n_930),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_939),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_949),
.B(n_854),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_906),
.B(n_854),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_893),
.Y(n_982)
);

AO221x1_ASAP7_75t_L g983 ( 
.A1(n_885),
.A2(n_679),
.B1(n_628),
.B2(n_639),
.C(n_626),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_904),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_909),
.B(n_849),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_898),
.B(n_865),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_L g987 ( 
.A(n_902),
.B(n_857),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_910),
.B(n_849),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_912),
.B(n_849),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_904),
.Y(n_990)
);

INVx8_ASAP7_75t_L g991 ( 
.A(n_953),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_907),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_921),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_914),
.B(n_922),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_L g995 ( 
.A(n_881),
.B(n_913),
.C(n_908),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_905),
.B(n_862),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_948),
.B(n_862),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_913),
.B(n_780),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_924),
.A2(n_820),
.B(n_870),
.C(n_846),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_924),
.B(n_787),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_933),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_937),
.B(n_865),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_937),
.B(n_787),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_952),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_929),
.B(n_865),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_934),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_933),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_L g1008 ( 
.A(n_952),
.B(n_667),
.C(n_622),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_946),
.B(n_866),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_938),
.B(n_797),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_953),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_923),
.B(n_849),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_891),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_887),
.B(n_888),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_892),
.B(n_797),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_931),
.B(n_866),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_936),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_907),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_936),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_871),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_872),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_896),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_915),
.B(n_870),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_940),
.B(n_866),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_877),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_941),
.B(n_669),
.C(n_668),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_876),
.A2(n_866),
.B1(n_870),
.B2(n_868),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_943),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_R g1029 ( 
.A(n_878),
.B(n_804),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_879),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_947),
.B(n_945),
.C(n_944),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_935),
.B(n_804),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_884),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_886),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_L g1035 ( 
.A(n_920),
.B(n_676),
.C(n_674),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_951),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_876),
.B(n_866),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_911),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_882),
.B(n_825),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_932),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_882),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_883),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_883),
.B(n_825),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_911),
.B(n_575),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_875),
.B(n_825),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_932),
.B(n_825),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_875),
.B(n_954),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_873),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_911),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_873),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_901),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_875),
.B(n_807),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_901),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_875),
.B(n_848),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_918),
.B(n_586),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_954),
.B(n_848),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_928),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_918),
.Y(n_1058)
);

INVx8_ASAP7_75t_L g1059 ( 
.A(n_897),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_918),
.B(n_593),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_928),
.B(n_601),
.C(n_595),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_SL g1062 ( 
.A(n_926),
.B(n_610),
.C(n_606),
.Y(n_1062)
);

INVxp33_ASAP7_75t_L g1063 ( 
.A(n_878),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_918),
.B(n_807),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_927),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_897),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_942),
.B(n_686),
.C(n_685),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_942),
.B(n_624),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_927),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_897),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_897),
.B(n_848),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_897),
.B(n_848),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_916),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_875),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_903),
.B(n_656),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_889),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_899),
.B(n_828),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_880),
.B(n_648),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_899),
.B(n_828),
.Y(n_1079)
);

BUFx2_ASAP7_75t_R g1080 ( 
.A(n_894),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_950),
.B(n_651),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_899),
.B(n_834),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_916),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_875),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_SL g1085 ( 
.A(n_903),
.B(n_579),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_880),
.B(n_654),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_L g1087 ( 
.A(n_995),
.B(n_657),
.Y(n_1087)
);

AO22x2_ASAP7_75t_L g1088 ( 
.A1(n_1035),
.A2(n_702),
.B1(n_522),
.B2(n_577),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_987),
.B(n_664),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_976),
.Y(n_1090)
);

OA22x2_ASAP7_75t_L g1091 ( 
.A1(n_978),
.A2(n_793),
.B1(n_794),
.B2(n_791),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_964),
.B(n_670),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1022),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1028),
.Y(n_1094)
);

AND2x6_ASAP7_75t_SL g1095 ( 
.A(n_1010),
.B(n_1015),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_979),
.B(n_800),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_1000),
.Y(n_1097)
);

BUFx8_ASAP7_75t_L g1098 ( 
.A(n_957),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_955),
.Y(n_1099)
);

AO22x2_ASAP7_75t_L g1100 ( 
.A1(n_969),
.A2(n_522),
.B1(n_577),
.B2(n_508),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1036),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_970),
.B(n_802),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1003),
.A2(n_539),
.B1(n_545),
.B2(n_534),
.Y(n_1103)
);

AO22x2_ASAP7_75t_L g1104 ( 
.A1(n_1029),
.A2(n_711),
.B1(n_630),
.B2(n_696),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_965),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_972),
.B(n_675),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1016),
.Y(n_1107)
);

AO22x2_ASAP7_75t_L g1108 ( 
.A1(n_1008),
.A2(n_711),
.B1(n_630),
.B2(n_701),
.Y(n_1108)
);

AO22x2_ASAP7_75t_L g1109 ( 
.A1(n_1026),
.A2(n_691),
.B1(n_707),
.B2(n_806),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_956),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1016),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_L g1112 ( 
.A(n_1084),
.B(n_694),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1032),
.B(n_579),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_991),
.Y(n_1114)
);

BUFx8_ASAP7_75t_L g1115 ( 
.A(n_1080),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_966),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1024),
.Y(n_1117)
);

BUFx8_ASAP7_75t_L g1118 ( 
.A(n_972),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1024),
.Y(n_1119)
);

BUFx8_ASAP7_75t_L g1120 ( 
.A(n_1023),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_998),
.B(n_699),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1077),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_974),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1077),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_982),
.Y(n_1125)
);

NAND2xp33_ASAP7_75t_L g1126 ( 
.A(n_1084),
.B(n_704),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_980),
.B(n_708),
.Y(n_1127)
);

AO22x2_ASAP7_75t_L g1128 ( 
.A1(n_1041),
.A2(n_692),
.B1(n_693),
.B2(n_672),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1076),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1079),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_966),
.B(n_834),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1079),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1082),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_996),
.B(n_713),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1082),
.Y(n_1135)
);

OAI221xp5_ASAP7_75t_L g1136 ( 
.A1(n_1078),
.A2(n_715),
.B1(n_679),
.B2(n_587),
.C(n_594),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_991),
.Y(n_1137)
);

AO22x2_ASAP7_75t_L g1138 ( 
.A1(n_1042),
.A2(n_693),
.B1(n_692),
.B2(n_583),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1052),
.B(n_500),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1014),
.B(n_997),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_994),
.A2(n_679),
.B1(n_604),
.B2(n_615),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_991),
.Y(n_1142)
);

AO22x2_ASAP7_75t_L g1143 ( 
.A1(n_983),
.A2(n_618),
.B1(n_637),
.B2(n_572),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_958),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_1011),
.B(n_1086),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_968),
.Y(n_1146)
);

AO22x2_ASAP7_75t_L g1147 ( 
.A1(n_1031),
.A2(n_645),
.B1(n_647),
.B2(n_641),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_993),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1006),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1040),
.B(n_608),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_967),
.A2(n_652),
.B1(n_663),
.B2(n_650),
.Y(n_1151)
);

AO22x2_ASAP7_75t_L g1152 ( 
.A1(n_1009),
.A2(n_688),
.B1(n_689),
.B2(n_671),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1001),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1064),
.B(n_842),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1007),
.Y(n_1155)
);

OAI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_1085),
.A2(n_1075),
.B1(n_1013),
.B2(n_994),
.C(n_966),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_971),
.B(n_842),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1017),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_SL g1159 ( 
.A1(n_960),
.A2(n_700),
.B1(n_703),
.B2(n_697),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1084),
.B(n_818),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1019),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1073),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1083),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_977),
.B(n_985),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_1070),
.B(n_553),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_981),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_981),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1020),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1004),
.B(n_843),
.Y(n_1169)
);

OAI221xp5_ASAP7_75t_L g1170 ( 
.A1(n_1081),
.A2(n_705),
.B1(n_712),
.B2(n_529),
.C(n_501),
.Y(n_1170)
);

AO22x2_ASAP7_75t_L g1171 ( 
.A1(n_1005),
.A2(n_1025),
.B1(n_1030),
.B2(n_1021),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1033),
.Y(n_1172)
);

AO22x2_ASAP7_75t_L g1173 ( 
.A1(n_1034),
.A2(n_571),
.B1(n_661),
.B2(n_660),
.Y(n_1173)
);

AO22x2_ASAP7_75t_L g1174 ( 
.A1(n_1063),
.A2(n_571),
.B1(n_661),
.B2(n_660),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_959),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_959),
.Y(n_1176)
);

AO22x2_ASAP7_75t_L g1177 ( 
.A1(n_985),
.A2(n_843),
.B1(n_506),
.B2(n_3),
.Y(n_1177)
);

AO22x2_ASAP7_75t_L g1178 ( 
.A1(n_988),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_988),
.B(n_989),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_962),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_989),
.B(n_818),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_962),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1012),
.B(n_818),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_1012),
.A2(n_5),
.B1(n_2),
.B2(n_4),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1046),
.Y(n_1185)
);

NAND2x1p5_ASAP7_75t_L g1186 ( 
.A(n_1084),
.B(n_818),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1062),
.B(n_818),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1051),
.B(n_836),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1038),
.B(n_492),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1047),
.A2(n_1074),
.B1(n_1037),
.B2(n_1002),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_984),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1067),
.B(n_836),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_990),
.B(n_836),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1047),
.B(n_836),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_992),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1037),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1196)
);

OAI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_961),
.A2(n_499),
.B1(n_503),
.B2(n_494),
.C(n_493),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1038),
.B(n_504),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1038),
.B(n_505),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1018),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1061),
.Y(n_1201)
);

BUFx8_ASAP7_75t_L g1202 ( 
.A(n_1048),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1056),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1057),
.B(n_836),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1045),
.B(n_844),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1039),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_986),
.B(n_510),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_1045),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1039),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1043),
.Y(n_1210)
);

AO22x2_ASAP7_75t_L g1211 ( 
.A1(n_1054),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1044),
.B(n_844),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1043),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1049),
.B(n_1058),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1054),
.B(n_1027),
.Y(n_1215)
);

AND2x6_ASAP7_75t_L g1216 ( 
.A(n_1049),
.B(n_520),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1050),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1053),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1072),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1071),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1055),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_963),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_973),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_975),
.A2(n_513),
.B1(n_519),
.B2(n_511),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1060),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1049),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1058),
.B(n_844),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1058),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1066),
.A2(n_527),
.B1(n_532),
.B2(n_530),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1068),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1059),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1059),
.B(n_535),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_999),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1069),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_1059),
.B(n_844),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1065),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_976),
.Y(n_1237)
);

AO22x2_ASAP7_75t_L g1238 ( 
.A1(n_1035),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1238)
);

NAND2x1p5_ASAP7_75t_L g1239 ( 
.A(n_957),
.B(n_844),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_957),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_978),
.A2(n_717),
.B1(n_537),
.B2(n_544),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_955),
.Y(n_1242)
);

BUFx8_ASAP7_75t_L g1243 ( 
.A(n_976),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_980),
.B(n_538),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_980),
.B(n_552),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1022),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1022),
.Y(n_1247)
);

AO22x2_ASAP7_75t_L g1248 ( 
.A1(n_1035),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1022),
.Y(n_1249)
);

OAI221xp5_ASAP7_75t_L g1250 ( 
.A1(n_1000),
.A2(n_557),
.B1(n_560),
.B2(n_559),
.C(n_555),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_957),
.Y(n_1251)
);

OAI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_1000),
.A2(n_568),
.B1(n_573),
.B2(n_570),
.C(n_562),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_957),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_987),
.B(n_580),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1022),
.Y(n_1255)
);

OAI221xp5_ASAP7_75t_L g1256 ( 
.A1(n_1000),
.A2(n_584),
.B1(n_590),
.B2(n_585),
.C(n_582),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_976),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_987),
.B(n_597),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_980),
.B(n_598),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1029),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_964),
.B(n_599),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_980),
.B(n_602),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_SL g1263 ( 
.A1(n_998),
.A2(n_603),
.B1(n_613),
.B2(n_607),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_978),
.B(n_14),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_980),
.B(n_614),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_955),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_955),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_957),
.B(n_15),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_955),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1022),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_980),
.B(n_619),
.Y(n_1271)
);

AO22x2_ASAP7_75t_L g1272 ( 
.A1(n_1035),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_980),
.B(n_620),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_980),
.B(n_625),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_976),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_955),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1097),
.A2(n_19),
.B(n_16),
.C(n_18),
.Y(n_1277)
);

OR2x6_ASAP7_75t_L g1278 ( 
.A(n_1114),
.B(n_520),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1175),
.B(n_18),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1176),
.B(n_1180),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1092),
.B(n_627),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1121),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_1282)
);

INVx4_ASAP7_75t_L g1283 ( 
.A(n_1251),
.Y(n_1283)
);

OAI21xp33_ASAP7_75t_L g1284 ( 
.A1(n_1103),
.A2(n_633),
.B(n_632),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1182),
.B(n_20),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1164),
.A2(n_635),
.B(n_634),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1115),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1140),
.A2(n_1179),
.B1(n_1167),
.B2(n_1166),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1206),
.A2(n_642),
.B(n_638),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1209),
.A2(n_644),
.B(n_643),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_1156),
.B(n_653),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1233),
.A2(n_683),
.B(n_520),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1210),
.A2(n_662),
.B(n_655),
.Y(n_1293)
);

CKINVDCx6p67_ASAP7_75t_R g1294 ( 
.A(n_1137),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1213),
.A2(n_666),
.B(n_665),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1205),
.A2(n_677),
.B(n_673),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1105),
.A2(n_678),
.B1(n_682),
.B2(n_681),
.Y(n_1297)
);

AOI21xp33_ASAP7_75t_L g1298 ( 
.A1(n_1139),
.A2(n_698),
.B(n_695),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1090),
.B(n_709),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1122),
.A2(n_716),
.B(n_710),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1124),
.A2(n_683),
.B(n_520),
.Y(n_1301)
);

AOI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1109),
.A2(n_1088),
.B1(n_1096),
.B2(n_1113),
.C(n_1108),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1093),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1130),
.A2(n_683),
.B(n_228),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1087),
.A2(n_1250),
.B(n_1256),
.C(n_1252),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1174),
.A2(n_683),
.B1(n_23),
.B2(n_21),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1149),
.B(n_22),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1132),
.B(n_23),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1142),
.B(n_24),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1260),
.B(n_24),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1237),
.B(n_25),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1275),
.B(n_25),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1094),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1133),
.A2(n_234),
.B(n_227),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1135),
.B(n_26),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1127),
.B(n_1150),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1134),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1116),
.B(n_27),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1234),
.A2(n_236),
.B(n_235),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_L g1320 ( 
.A(n_1257),
.B(n_238),
.Y(n_1320)
);

AO32x2_ASAP7_75t_L g1321 ( 
.A1(n_1141),
.A2(n_31),
.A3(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_1321)
);

AOI221xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1264),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.C(n_34),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1243),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1151),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1101),
.B(n_36),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1236),
.A2(n_241),
.B(n_240),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1136),
.A2(n_40),
.B(n_37),
.C(n_38),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1095),
.B(n_37),
.Y(n_1328)
);

OR2x2_ASAP7_75t_SL g1329 ( 
.A(n_1118),
.B(n_41),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1194),
.A2(n_246),
.B(n_244),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1246),
.B(n_41),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1247),
.B(n_1249),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1255),
.A2(n_47),
.B1(n_42),
.B2(n_44),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1270),
.B(n_44),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1109),
.B(n_47),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1107),
.B(n_48),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1111),
.B(n_49),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1181),
.A2(n_248),
.B(n_247),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_SL g1339 ( 
.A(n_1240),
.B(n_49),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1117),
.B(n_50),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1203),
.A2(n_254),
.B(n_250),
.Y(n_1341)
);

AO32x1_ASAP7_75t_L g1342 ( 
.A1(n_1154),
.A2(n_53),
.A3(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1089),
.B(n_51),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1201),
.A2(n_55),
.B(n_52),
.C(n_54),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1102),
.B(n_55),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1119),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1145),
.B(n_57),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1217),
.A2(n_58),
.B(n_59),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1215),
.A2(n_256),
.B(n_255),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1263),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1350)
);

NOR3xp33_ASAP7_75t_L g1351 ( 
.A(n_1106),
.B(n_1170),
.C(n_1254),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1168),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1172),
.B(n_61),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1261),
.B(n_62),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1185),
.B(n_63),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1268),
.B(n_63),
.Y(n_1356)
);

AO21x1_ASAP7_75t_L g1357 ( 
.A1(n_1219),
.A2(n_259),
.B(n_257),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1244),
.B(n_64),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1245),
.B(n_64),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1258),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1159),
.B(n_65),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1231),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1227),
.A2(n_265),
.B(n_264),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1259),
.B(n_67),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1099),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1262),
.B(n_68),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1131),
.B(n_68),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1241),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1368)
);

CKINVDCx10_ASAP7_75t_R g1369 ( 
.A(n_1098),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1221),
.A2(n_1225),
.B(n_1198),
.C(n_1199),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1253),
.A2(n_72),
.B1(n_69),
.B2(n_70),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1214),
.A2(n_267),
.B(n_266),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1104),
.B(n_72),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1169),
.B(n_73),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1189),
.A2(n_1197),
.B(n_1230),
.C(n_1265),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1216),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1271),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1147),
.A2(n_78),
.B1(n_74),
.B2(n_77),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1112),
.A2(n_270),
.B(n_268),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1202),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1273),
.B(n_78),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1126),
.A2(n_273),
.B(n_272),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1222),
.A2(n_276),
.B(n_274),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1274),
.B(n_79),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1144),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1104),
.B(n_80),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1146),
.B(n_82),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1120),
.B(n_82),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1223),
.A2(n_278),
.B(n_277),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1148),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1153),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1229),
.B(n_83),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1155),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1091),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_1183),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1147),
.B(n_84),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1100),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1160),
.A2(n_280),
.B(n_279),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1108),
.B(n_86),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1216),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1158),
.B(n_87),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_SL g1402 ( 
.A(n_1232),
.B(n_88),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1161),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1162),
.B(n_88),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1226),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1187),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1207),
.B(n_89),
.C(n_90),
.Y(n_1407)
);

NOR3xp33_ASAP7_75t_L g1408 ( 
.A(n_1163),
.B(n_89),
.C(n_90),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1174),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1216),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1218),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1220),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1412)
);

NOR3xp33_ASAP7_75t_L g1413 ( 
.A(n_1238),
.B(n_95),
.C(n_97),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1191),
.A2(n_100),
.B(n_98),
.C(n_99),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1088),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.C(n_101),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1228),
.B(n_1200),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_SL g1417 ( 
.A1(n_1110),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1224),
.B(n_102),
.C(n_103),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_SL g1419 ( 
.A1(n_1123),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1212),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1157),
.A2(n_283),
.B(n_281),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1192),
.B(n_105),
.Y(n_1422)
);

OA22x2_ASAP7_75t_L g1423 ( 
.A1(n_1125),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1239),
.Y(n_1424)
);

OAI21xp33_ASAP7_75t_L g1425 ( 
.A1(n_1178),
.A2(n_108),
.B(n_110),
.Y(n_1425)
);

NOR2xp67_ASAP7_75t_SL g1426 ( 
.A(n_1178),
.B(n_111),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1100),
.B(n_111),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1195),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1186),
.A2(n_287),
.B(n_286),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1235),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1129),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1188),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1242),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1266),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1173),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1276),
.B(n_112),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1204),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1267),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1190),
.A2(n_291),
.B(n_289),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1208),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1440)
);

INVx5_ASAP7_75t_L g1441 ( 
.A(n_1165),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1269),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1208),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1443)
);

INVx11_ASAP7_75t_L g1444 ( 
.A(n_1165),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1138),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1138),
.B(n_115),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1238),
.B(n_116),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1193),
.Y(n_1448)
);

AOI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1171),
.A2(n_295),
.B(n_294),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1128),
.B(n_116),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1128),
.B(n_1173),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1152),
.B(n_117),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1171),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1248),
.Y(n_1454)
);

AOI22x1_ASAP7_75t_L g1455 ( 
.A1(n_1196),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1248),
.A2(n_121),
.B1(n_118),
.B2(n_120),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1190),
.A2(n_299),
.B(n_297),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1152),
.A2(n_303),
.B(n_300),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1177),
.A2(n_305),
.B(n_304),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1165),
.B(n_122),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1177),
.A2(n_1196),
.B(n_1211),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1272),
.B(n_1143),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1211),
.A2(n_127),
.B1(n_123),
.B2(n_124),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1272),
.B(n_124),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1280),
.B(n_1143),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1288),
.B(n_1184),
.Y(n_1466)
);

INVx6_ASAP7_75t_SL g1467 ( 
.A(n_1367),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1369),
.Y(n_1468)
);

BUFx4f_ASAP7_75t_SL g1469 ( 
.A(n_1294),
.Y(n_1469)
);

CKINVDCx8_ASAP7_75t_R g1470 ( 
.A(n_1287),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1307),
.B(n_1184),
.Y(n_1471)
);

BUFx8_ASAP7_75t_L g1472 ( 
.A(n_1318),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1422),
.Y(n_1473)
);

NOR3xp33_ASAP7_75t_L g1474 ( 
.A(n_1281),
.B(n_1328),
.C(n_1413),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1376),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1335),
.B(n_127),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1400),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1367),
.B(n_128),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1329),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1332),
.B(n_129),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1303),
.Y(n_1481)
);

OR2x6_ASAP7_75t_L g1482 ( 
.A(n_1422),
.B(n_130),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1352),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1313),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1390),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1318),
.B(n_131),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1456),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1487)
);

AO22x1_ASAP7_75t_L g1488 ( 
.A1(n_1447),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1393),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1403),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1316),
.B(n_1302),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1373),
.B(n_134),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1365),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_SL g1494 ( 
.A1(n_1371),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1386),
.B(n_137),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1433),
.B(n_138),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1399),
.B(n_138),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1323),
.Y(n_1498)
);

BUFx4f_ASAP7_75t_L g1499 ( 
.A(n_1400),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1428),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1434),
.Y(n_1501)
);

NAND2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1283),
.B(n_308),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1298),
.B(n_139),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_R g1504 ( 
.A(n_1388),
.B(n_311),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1394),
.B(n_139),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1431),
.Y(n_1506)
);

AOI22x1_ASAP7_75t_L g1507 ( 
.A1(n_1286),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1435),
.B(n_140),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1384),
.B(n_142),
.Y(n_1509)
);

BUFx4f_ASAP7_75t_L g1510 ( 
.A(n_1400),
.Y(n_1510)
);

AND3x1_ASAP7_75t_SL g1511 ( 
.A(n_1415),
.B(n_143),
.C(n_144),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1438),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1442),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1362),
.B(n_143),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1387),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1410),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1305),
.A2(n_315),
.B(n_314),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1353),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1299),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1339),
.B(n_144),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1454),
.B(n_145),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1325),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1362),
.B(n_145),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1410),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1425),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1309),
.B(n_146),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1309),
.B(n_1423),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1331),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1448),
.B(n_148),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1334),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1279),
.B(n_149),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1380),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1442),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1401),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_SL g1535 ( 
.A(n_1310),
.B(n_150),
.C(n_151),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1405),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1405),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1404),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1285),
.B(n_152),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1464),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1291),
.B(n_1375),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1308),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1376),
.Y(n_1543)
);

INVxp33_ASAP7_75t_SL g1544 ( 
.A(n_1297),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1416),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1462),
.A2(n_160),
.B1(n_157),
.B2(n_158),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1315),
.B(n_157),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1432),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1410),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1453),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1283),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1336),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1337),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1445),
.B(n_160),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1340),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1355),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1356),
.B(n_161),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1436),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1444),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1351),
.B(n_161),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1432),
.B(n_162),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1450),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1430),
.B(n_320),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1437),
.B(n_1395),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1446),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1452),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1396),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1427),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1345),
.B(n_162),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1343),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1378),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1437),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1420),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1374),
.B(n_166),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1278),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1358),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1295),
.B(n_166),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1359),
.Y(n_1578)
);

AOI221x1_ASAP7_75t_L g1579 ( 
.A1(n_1461),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1409),
.B(n_169),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1364),
.Y(n_1581)
);

NAND2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1441),
.B(n_321),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1366),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1430),
.Y(n_1584)
);

BUFx8_ASAP7_75t_L g1585 ( 
.A(n_1321),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1426),
.B(n_171),
.C(n_172),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1441),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1460),
.B(n_172),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1441),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1420),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1381),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1451),
.Y(n_1592)
);

BUFx4f_ASAP7_75t_L g1593 ( 
.A(n_1278),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1406),
.B(n_173),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1320),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1397),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1377),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1282),
.A2(n_173),
.B(n_175),
.C(n_176),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1407),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1424),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1350),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1346),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1306),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1424),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1317),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1424),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1455),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_1607)
);

CKINVDCx8_ASAP7_75t_R g1608 ( 
.A(n_1370),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1391),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1361),
.B(n_182),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1411),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1398),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1392),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1449),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1354),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1348),
.B(n_183),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1429),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1333),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1440),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_L g1620 ( 
.A(n_1341),
.B(n_322),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1475),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1499),
.B(n_1347),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1482),
.B(n_1439),
.Y(n_1623)
);

OR2x6_ASAP7_75t_SL g1624 ( 
.A(n_1532),
.B(n_1468),
.Y(n_1624)
);

NAND2x1p5_ASAP7_75t_L g1625 ( 
.A(n_1499),
.B(n_1402),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1481),
.Y(n_1626)
);

NAND2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1510),
.B(n_1457),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1484),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1482),
.A2(n_1463),
.B1(n_1443),
.B2(n_1324),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1476),
.B(n_1408),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1485),
.Y(n_1631)
);

A2O1A1Ixp33_ASAP7_75t_SL g1632 ( 
.A1(n_1503),
.A2(n_1277),
.B(n_1344),
.C(n_1412),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1475),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1482),
.A2(n_1418),
.B1(n_1327),
.B2(n_1368),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1473),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1483),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1544),
.B(n_1311),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1493),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1466),
.B(n_1322),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1517),
.A2(n_1382),
.B(n_1379),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1469),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1510),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1506),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1545),
.B(n_1312),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1492),
.B(n_1321),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1491),
.B(n_1360),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1564),
.Y(n_1647)
);

NAND2xp33_ASAP7_75t_L g1648 ( 
.A(n_1474),
.B(n_1551),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1472),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1558),
.B(n_1385),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1509),
.A2(n_1458),
.B(n_1459),
.C(n_1414),
.Y(n_1651)
);

A2O1A1Ixp33_ASAP7_75t_SL g1652 ( 
.A1(n_1605),
.A2(n_1289),
.B(n_1293),
.C(n_1290),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1515),
.B(n_1518),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1495),
.B(n_1321),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1489),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1596),
.A2(n_1300),
.B1(n_1314),
.B2(n_1319),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1466),
.B(n_1417),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1465),
.B(n_1419),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1472),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1585),
.A2(n_1304),
.B1(n_1349),
.B2(n_1342),
.Y(n_1660)
);

INVx5_ASAP7_75t_L g1661 ( 
.A(n_1477),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1467),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1543),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1570),
.B(n_1284),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1498),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1601),
.A2(n_1296),
.B(n_1421),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1478),
.B(n_186),
.Y(n_1667)
);

AOI222xp33_ASAP7_75t_L g1668 ( 
.A1(n_1479),
.A2(n_1342),
.B1(n_189),
.B2(n_190),
.C1(n_191),
.C2(n_192),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1477),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1552),
.B(n_1338),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1512),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1553),
.B(n_1330),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1620),
.A2(n_1342),
.B(n_1383),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1585),
.A2(n_1357),
.B1(n_1301),
.B2(n_1326),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1620),
.A2(n_1363),
.B(n_1389),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1470),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1467),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1541),
.A2(n_1372),
.B(n_1292),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1500),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1560),
.A2(n_1616),
.B(n_1607),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1490),
.Y(n_1681)
);

AND3x2_ASAP7_75t_L g1682 ( 
.A(n_1527),
.B(n_1519),
.C(n_1520),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1555),
.B(n_187),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1548),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1501),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1543),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1617),
.A2(n_189),
.B(n_190),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1497),
.B(n_191),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1477),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1559),
.Y(n_1690)
);

NAND2xp33_ASAP7_75t_L g1691 ( 
.A(n_1616),
.B(n_193),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1604),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1568),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1567),
.B(n_193),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1487),
.A2(n_1494),
.B1(n_1471),
.B2(n_1619),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1608),
.B(n_195),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1486),
.B(n_1526),
.Y(n_1697)
);

NOR2xp67_ASAP7_75t_SL g1698 ( 
.A(n_1586),
.B(n_1613),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1536),
.Y(n_1699)
);

AND2x2_ASAP7_75t_SL g1700 ( 
.A(n_1593),
.B(n_195),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1571),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1505),
.B(n_198),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1607),
.A2(n_199),
.B(n_200),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1566),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1516),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1612),
.A2(n_1614),
.B(n_1589),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1584),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1593),
.B(n_325),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1465),
.B(n_199),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1592),
.B(n_201),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1556),
.B(n_201),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1513),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1537),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1554),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1565),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1575),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1516),
.B(n_202),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1516),
.B(n_1524),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1504),
.Y(n_1719)
);

INVx3_ASAP7_75t_SL g1720 ( 
.A(n_1573),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1524),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1612),
.A2(n_1542),
.B(n_1577),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1521),
.B(n_1569),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1522),
.B(n_202),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1562),
.B(n_203),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1524),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1533),
.Y(n_1727)
);

AO21x2_ASAP7_75t_L g1728 ( 
.A1(n_1611),
.A2(n_327),
.B(n_326),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1529),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1550),
.Y(n_1730)
);

OR2x6_ASAP7_75t_SL g1731 ( 
.A(n_1496),
.B(n_203),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1576),
.A2(n_204),
.B(n_205),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1590),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1557),
.B(n_204),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1529),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1574),
.B(n_205),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1572),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1647),
.B(n_1578),
.Y(n_1738)
);

O2A1O1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1632),
.A2(n_1598),
.B(n_1535),
.C(n_1588),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1723),
.B(n_1581),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1697),
.B(n_1583),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1626),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1628),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1695),
.A2(n_1571),
.B1(n_1525),
.B2(n_1487),
.Y(n_1744)
);

OR2x2_ASAP7_75t_SL g1745 ( 
.A(n_1694),
.B(n_1586),
.Y(n_1745)
);

AND2x2_ASAP7_75t_SL g1746 ( 
.A(n_1700),
.B(n_1691),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1701),
.A2(n_1525),
.B1(n_1494),
.B2(n_1601),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1645),
.B(n_1591),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1631),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1701),
.A2(n_1703),
.B1(n_1540),
.B2(n_1619),
.Y(n_1750)
);

AOI21x1_ASAP7_75t_SL g1751 ( 
.A1(n_1650),
.A2(n_1523),
.B(n_1514),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1654),
.B(n_1508),
.Y(n_1752)
);

O2A1O1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1696),
.A2(n_1597),
.B(n_1599),
.C(n_1531),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1635),
.B(n_1549),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1647),
.B(n_1480),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1703),
.A2(n_1579),
.B(n_1582),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1655),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1630),
.B(n_1488),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1684),
.B(n_1549),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1692),
.B(n_1584),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1688),
.B(n_1528),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1693),
.B(n_1480),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1729),
.B(n_1530),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1667),
.B(n_1702),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1704),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1640),
.A2(n_1539),
.B(n_1531),
.Y(n_1766)
);

NAND2x1p5_ASAP7_75t_L g1767 ( 
.A(n_1661),
.B(n_1587),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1653),
.B(n_1534),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1681),
.B(n_1549),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1679),
.B(n_1538),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1734),
.B(n_1615),
.Y(n_1771)
);

BUFx2_ASAP7_75t_R g1772 ( 
.A(n_1649),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1736),
.B(n_1580),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1735),
.B(n_1602),
.Y(n_1774)
);

A2O1A1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1680),
.A2(n_1539),
.B(n_1547),
.C(n_1609),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1715),
.B(n_1618),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1685),
.Y(n_1777)
);

OR2x6_ASAP7_75t_SL g1778 ( 
.A(n_1665),
.B(n_1547),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1707),
.B(n_1606),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1643),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1710),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1671),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1714),
.B(n_1606),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1680),
.B(n_1595),
.Y(n_1784)
);

OAI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1675),
.A2(n_1563),
.B(n_1502),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1642),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1657),
.B(n_1639),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1634),
.A2(n_1610),
.B(n_1594),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1718),
.B(n_1699),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1629),
.B(n_1540),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1656),
.A2(n_1507),
.B(n_1561),
.Y(n_1791)
);

O2A1O1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1634),
.A2(n_1546),
.B(n_1603),
.C(n_1511),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1657),
.B(n_1600),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1716),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1661),
.B(n_1587),
.Y(n_1795)
);

O2A1O1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1651),
.A2(n_1479),
.B(n_1589),
.C(n_208),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1699),
.B(n_1713),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1730),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1639),
.B(n_1600),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1636),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1676),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1709),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1646),
.A2(n_1600),
.B(n_207),
.C(n_208),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1709),
.B(n_206),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1713),
.B(n_207),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1638),
.Y(n_1806)
);

OAI21xp33_ASAP7_75t_L g1807 ( 
.A1(n_1790),
.A2(n_1668),
.B(n_1637),
.Y(n_1807)
);

OR2x2_ASAP7_75t_SL g1808 ( 
.A(n_1781),
.B(n_1710),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1742),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1750),
.A2(n_1668),
.B1(n_1629),
.B2(n_1623),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1765),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1790),
.A2(n_1623),
.B1(n_1731),
.B2(n_1664),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1750),
.A2(n_1682),
.B(n_1732),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1748),
.B(n_1706),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1806),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1744),
.A2(n_1666),
.B1(n_1660),
.B2(n_1698),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1744),
.A2(n_1666),
.B1(n_1658),
.B2(n_1674),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1762),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1747),
.A2(n_1728),
.B1(n_1719),
.B2(n_1658),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1747),
.A2(n_1648),
.B1(n_1717),
.B2(n_1708),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1746),
.A2(n_1712),
.B1(n_1727),
.B2(n_1737),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_SL g1822 ( 
.A1(n_1758),
.A2(n_1728),
.B1(n_1708),
.B2(n_1725),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1798),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1800),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1759),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1752),
.A2(n_1773),
.B1(n_1771),
.B2(n_1802),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1778),
.A2(n_1711),
.B1(n_1683),
.B2(n_1687),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1801),
.B(n_1624),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1745),
.A2(n_1625),
.B1(n_1724),
.B2(n_1717),
.Y(n_1829)
);

OAI222xp33_ASAP7_75t_L g1830 ( 
.A1(n_1796),
.A2(n_1670),
.B1(n_1672),
.B2(n_1644),
.C1(n_1722),
.C2(n_1673),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1743),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1749),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1757),
.B(n_1621),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1759),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1777),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1741),
.B(n_1621),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1787),
.B(n_1633),
.Y(n_1837)
);

BUFx12f_ASAP7_75t_L g1838 ( 
.A(n_1786),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1804),
.A2(n_1622),
.B1(n_1625),
.B2(n_1627),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1791),
.A2(n_1784),
.B1(n_1787),
.B2(n_1805),
.Y(n_1840)
);

AOI222xp33_ASAP7_75t_L g1841 ( 
.A1(n_1775),
.A2(n_1720),
.B1(n_1733),
.B2(n_1652),
.C1(n_1677),
.C2(n_1662),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1764),
.A2(n_1659),
.B1(n_1627),
.B2(n_1622),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1792),
.A2(n_1633),
.B1(n_1663),
.B2(n_1686),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1809),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1837),
.B(n_1740),
.Y(n_1845)
);

INVxp33_ASAP7_75t_L g1846 ( 
.A(n_1818),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1807),
.A2(n_1784),
.B1(n_1803),
.B2(n_1789),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1837),
.B(n_1779),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1836),
.B(n_1761),
.Y(n_1849)
);

AOI211xp5_ASAP7_75t_L g1850 ( 
.A1(n_1812),
.A2(n_1813),
.B(n_1827),
.C(n_1829),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1815),
.Y(n_1851)
);

INVx5_ASAP7_75t_L g1852 ( 
.A(n_1838),
.Y(n_1852)
);

AOI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1839),
.A2(n_1788),
.B(n_1753),
.C(n_1756),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1810),
.A2(n_1816),
.B1(n_1820),
.B2(n_1817),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1836),
.B(n_1760),
.Y(n_1855)
);

BUFx12f_ASAP7_75t_L g1856 ( 
.A(n_1838),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1819),
.A2(n_1766),
.B(n_1739),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1809),
.Y(n_1858)
);

HB1xp67_ASAP7_75t_L g1859 ( 
.A(n_1811),
.Y(n_1859)
);

OAI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1840),
.A2(n_1799),
.B1(n_1794),
.B2(n_1774),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1811),
.B(n_1755),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1814),
.B(n_1797),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1822),
.A2(n_1799),
.B1(n_1793),
.B2(n_1769),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1830),
.A2(n_1763),
.B1(n_1776),
.B2(n_1738),
.C(n_1783),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1842),
.A2(n_1776),
.B1(n_1663),
.B2(n_1686),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1815),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1831),
.Y(n_1867)
);

O2A1O1Ixp33_ASAP7_75t_L g1868 ( 
.A1(n_1843),
.A2(n_1793),
.B(n_1769),
.C(n_1770),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1844),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1862),
.B(n_1814),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1858),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1845),
.B(n_1825),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1859),
.B(n_1833),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1868),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1857),
.A2(n_1821),
.B1(n_1841),
.B2(n_1826),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1856),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1845),
.B(n_1825),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1867),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1862),
.B(n_1834),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1856),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1861),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1849),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1849),
.Y(n_1883)
);

NAND2x1_ASAP7_75t_L g1884 ( 
.A(n_1848),
.B(n_1832),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1848),
.B(n_1846),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1870),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1885),
.B(n_1855),
.Y(n_1887)
);

CKINVDCx20_ASAP7_75t_R g1888 ( 
.A(n_1880),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1869),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1874),
.A2(n_1853),
.B(n_1850),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1869),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1870),
.Y(n_1892)
);

NAND3xp33_ASAP7_75t_L g1893 ( 
.A(n_1875),
.B(n_1864),
.C(n_1860),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1887),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1886),
.B(n_1885),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1889),
.B(n_1881),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1892),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1891),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1898),
.B(n_1890),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1897),
.A2(n_1893),
.B1(n_1890),
.B2(n_1854),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1895),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1894),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1898),
.A2(n_1863),
.B1(n_1847),
.B2(n_1865),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1896),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1899),
.B(n_1882),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1899),
.B(n_1883),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1904),
.B(n_1878),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1905),
.A2(n_1900),
.B1(n_1903),
.B2(n_1902),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1906),
.Y(n_1909)
);

NAND3xp33_ASAP7_75t_L g1910 ( 
.A(n_1908),
.B(n_1907),
.C(n_1901),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1910),
.B(n_1909),
.Y(n_1911)
);

AOI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1876),
.B1(n_1828),
.B2(n_1888),
.C(n_1880),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1911),
.B(n_1641),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1913),
.B(n_1884),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1912),
.B(n_1876),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1888),
.B1(n_1690),
.B2(n_1878),
.C(n_1846),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_R g1917 ( 
.A(n_1914),
.B(n_209),
.Y(n_1917)
);

A2O1A1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1914),
.A2(n_1772),
.B(n_1884),
.C(n_1870),
.Y(n_1918)
);

XNOR2xp5_ASAP7_75t_L g1919 ( 
.A(n_1916),
.B(n_1808),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1917),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1918),
.B(n_1871),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1920),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1919),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1921),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1920),
.A2(n_1879),
.B1(n_1871),
.B2(n_1877),
.Y(n_1925)
);

AND3x4_ASAP7_75t_L g1926 ( 
.A(n_1919),
.B(n_1879),
.C(n_1852),
.Y(n_1926)
);

AND3x4_ASAP7_75t_L g1927 ( 
.A(n_1919),
.B(n_1879),
.C(n_1852),
.Y(n_1927)
);

AND3x1_ASAP7_75t_L g1928 ( 
.A(n_1920),
.B(n_1873),
.C(n_1872),
.Y(n_1928)
);

NOR3xp33_ASAP7_75t_L g1929 ( 
.A(n_1922),
.B(n_209),
.C(n_210),
.Y(n_1929)
);

OAI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1924),
.A2(n_1877),
.B(n_1872),
.Y(n_1930)
);

AOI221xp5_ASAP7_75t_L g1931 ( 
.A1(n_1923),
.A2(n_1835),
.B1(n_1751),
.B2(n_213),
.C(n_215),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1926),
.A2(n_211),
.B(n_212),
.Y(n_1932)
);

AOI322xp5_ASAP7_75t_L g1933 ( 
.A1(n_1927),
.A2(n_1808),
.A3(n_1754),
.B1(n_1852),
.B2(n_1782),
.C1(n_1780),
.C2(n_1855),
.Y(n_1933)
);

NAND4xp25_ASAP7_75t_L g1934 ( 
.A(n_1925),
.B(n_215),
.C(n_216),
.D(n_218),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1928),
.B(n_219),
.Y(n_1935)
);

NAND4xp75_ASAP7_75t_L g1936 ( 
.A(n_1924),
.B(n_219),
.C(n_220),
.D(n_221),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1922),
.A2(n_222),
.B(n_223),
.Y(n_1937)
);

AND3x4_ASAP7_75t_L g1938 ( 
.A(n_1929),
.B(n_222),
.C(n_224),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1936),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1935),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1934),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1931),
.A2(n_1932),
.B1(n_1937),
.B2(n_1930),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1933),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1935),
.A2(n_1852),
.B1(n_1642),
.B2(n_1786),
.Y(n_1944)
);

AO22x2_ASAP7_75t_L g1945 ( 
.A1(n_1936),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1936),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1936),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1935),
.A2(n_1642),
.B1(n_1786),
.B2(n_1833),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1936),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_1935),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1936),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1936),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1935),
.A2(n_1768),
.B1(n_1689),
.B2(n_1726),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1936),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1936),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1936),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1936),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1930),
.B(n_226),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1936),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1935),
.A2(n_1726),
.B1(n_1721),
.B2(n_1689),
.Y(n_1960)
);

AOI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1941),
.A2(n_1940),
.B(n_1959),
.C(n_1951),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1950),
.B(n_1721),
.Y(n_1962)
);

NAND4xp75_ASAP7_75t_L g1963 ( 
.A(n_1947),
.B(n_1678),
.C(n_329),
.D(n_330),
.Y(n_1963)
);

NOR2x1_ASAP7_75t_L g1964 ( 
.A(n_1949),
.B(n_1669),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1945),
.Y(n_1965)
);

OAI211xp5_ASAP7_75t_L g1966 ( 
.A1(n_1946),
.A2(n_1661),
.B(n_1705),
.C(n_1669),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1958),
.Y(n_1967)
);

AOI221xp5_ASAP7_75t_L g1968 ( 
.A1(n_1943),
.A2(n_1669),
.B1(n_1705),
.B2(n_1823),
.C(n_1824),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1945),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1954),
.Y(n_1970)
);

AOI222xp33_ASAP7_75t_L g1971 ( 
.A1(n_1952),
.A2(n_1705),
.B1(n_1823),
.B2(n_1824),
.C1(n_1718),
.C2(n_1866),
.Y(n_1971)
);

XOR2x2_ASAP7_75t_L g1972 ( 
.A(n_1938),
.B(n_1767),
.Y(n_1972)
);

A2O1A1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1942),
.A2(n_1785),
.B(n_1851),
.C(n_1866),
.Y(n_1973)
);

OAI211xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1955),
.A2(n_328),
.B(n_331),
.C(n_333),
.Y(n_1974)
);

AOI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1956),
.A2(n_336),
.B(n_337),
.C(n_338),
.Y(n_1975)
);

NOR3xp33_ASAP7_75t_L g1976 ( 
.A(n_1939),
.B(n_339),
.C(n_340),
.Y(n_1976)
);

OAI211xp5_ASAP7_75t_L g1977 ( 
.A1(n_1957),
.A2(n_342),
.B(n_346),
.C(n_347),
.Y(n_1977)
);

NAND4xp75_ASAP7_75t_L g1978 ( 
.A(n_1948),
.B(n_348),
.C(n_350),
.D(n_352),
.Y(n_1978)
);

NAND4xp25_ASAP7_75t_L g1979 ( 
.A(n_1960),
.B(n_1834),
.C(n_355),
.D(n_357),
.Y(n_1979)
);

XNOR2xp5_ASAP7_75t_L g1980 ( 
.A(n_1961),
.B(n_1944),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1965),
.Y(n_1981)
);

NAND4xp25_ASAP7_75t_L g1982 ( 
.A(n_1970),
.B(n_1953),
.C(n_358),
.D(n_359),
.Y(n_1982)
);

AOI21xp33_ASAP7_75t_L g1983 ( 
.A1(n_1969),
.A2(n_354),
.B(n_360),
.Y(n_1983)
);

NOR4xp25_ASAP7_75t_L g1984 ( 
.A(n_1967),
.B(n_361),
.C(n_362),
.D(n_364),
.Y(n_1984)
);

NAND4xp25_ASAP7_75t_L g1985 ( 
.A(n_1964),
.B(n_368),
.C(n_369),
.D(n_370),
.Y(n_1985)
);

NOR4xp75_ASAP7_75t_L g1986 ( 
.A(n_1978),
.B(n_371),
.C(n_373),
.D(n_377),
.Y(n_1986)
);

NAND5xp2_ASAP7_75t_L g1987 ( 
.A(n_1966),
.B(n_1795),
.C(n_1767),
.D(n_385),
.E(n_386),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1962),
.B(n_1979),
.Y(n_1988)
);

NAND4xp25_ASAP7_75t_L g1989 ( 
.A(n_1976),
.B(n_1974),
.C(n_1975),
.D(n_1968),
.Y(n_1989)
);

AND4x1_ASAP7_75t_L g1990 ( 
.A(n_1972),
.B(n_382),
.C(n_384),
.D(n_392),
.Y(n_1990)
);

XOR2x2_ASAP7_75t_L g1991 ( 
.A(n_1980),
.B(n_1963),
.Y(n_1991)
);

AND4x1_ASAP7_75t_L g1992 ( 
.A(n_1981),
.B(n_1971),
.C(n_1977),
.D(n_1973),
.Y(n_1992)
);

NAND3x1_ASAP7_75t_L g1993 ( 
.A(n_1988),
.B(n_394),
.C(n_395),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1990),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_1987),
.B1(n_1989),
.B2(n_1982),
.Y(n_1995)
);

XNOR2xp5_ASAP7_75t_L g1996 ( 
.A(n_1991),
.B(n_1986),
.Y(n_1996)
);

OAI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1992),
.A2(n_1985),
.B1(n_1983),
.B2(n_1984),
.Y(n_1997)
);

AOI221x1_ASAP7_75t_L g1998 ( 
.A1(n_1993),
.A2(n_396),
.B1(n_397),
.B2(n_400),
.C(n_402),
.Y(n_1998)
);

OAI322xp33_ASAP7_75t_L g1999 ( 
.A1(n_1997),
.A2(n_1795),
.A3(n_404),
.B1(n_405),
.B2(n_407),
.C1(n_408),
.C2(n_409),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1996),
.Y(n_2000)
);

AOI22xp33_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1995),
.B1(n_1999),
.B2(n_1998),
.Y(n_2001)
);

XNOR2xp5_ASAP7_75t_L g2002 ( 
.A(n_2001),
.B(n_403),
.Y(n_2002)
);

OAI321xp33_ASAP7_75t_L g2003 ( 
.A1(n_2002),
.A2(n_411),
.A3(n_413),
.B1(n_414),
.B2(n_415),
.C(n_416),
.Y(n_2003)
);

AOI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_2003),
.A2(n_418),
.B1(n_421),
.B2(n_422),
.C(n_424),
.Y(n_2004)
);

AOI211xp5_ASAP7_75t_L g2005 ( 
.A1(n_2004),
.A2(n_425),
.B(n_426),
.C(n_427),
.Y(n_2005)
);


endmodule