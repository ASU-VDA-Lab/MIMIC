module fake_jpeg_10924_n_379 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_60),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_58),
.Y(n_135)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_59),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_61),
.B(n_81),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_62),
.Y(n_128)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_82),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_31),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g83 ( 
.A(n_23),
.B(n_3),
.CON(n_83),
.SN(n_83)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_52),
.Y(n_125)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_4),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_4),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_25),
.B(n_7),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_90),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_25),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_7),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_96),
.Y(n_119)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_35),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_35),
.B(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_38),
.Y(n_129)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_103),
.Y(n_161)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_105),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_63),
.A2(n_52),
.B1(n_51),
.B2(n_44),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_142),
.B1(n_143),
.B2(n_148),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_125),
.B(n_100),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_38),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_126),
.B(n_138),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_129),
.B(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_82),
.B(n_37),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_66),
.A2(n_51),
.B1(n_44),
.B2(n_43),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_145),
.B1(n_71),
.B2(n_104),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_43),
.B1(n_34),
.B2(n_32),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_95),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_37),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_68),
.A2(n_39),
.B1(n_45),
.B2(n_42),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_36),
.B1(n_42),
.B2(n_41),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_146),
.A2(n_73),
.B(n_83),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_62),
.A2(n_39),
.B1(n_45),
.B2(n_41),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_72),
.A2(n_47),
.B1(n_12),
.B2(n_13),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_148),
.B1(n_125),
.B2(n_143),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_70),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_47),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_87),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_58),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_56),
.B(n_10),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_163),
.B(n_67),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_166),
.A2(n_170),
.B1(n_207),
.B2(n_176),
.Y(n_241)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_99),
.B1(n_101),
.B2(n_69),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_128),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_175),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_77),
.B1(n_78),
.B2(n_94),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_172),
.A2(n_191),
.B1(n_215),
.B2(n_195),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_64),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_173),
.B(n_178),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_187),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_124),
.B(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_110),
.B(n_13),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_177),
.B(n_180),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_117),
.B(n_102),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_113),
.B(n_13),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_119),
.B(n_14),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_189),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_114),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_116),
.B(n_92),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_54),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_190),
.B(n_197),
.C(n_200),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_133),
.A2(n_62),
.B1(n_55),
.B2(n_75),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_192),
.B(n_198),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_216),
.B1(n_120),
.B2(n_151),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_89),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_115),
.B(n_89),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_80),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

BUFx24_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_115),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_108),
.B(n_84),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_205),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_156),
.B(n_59),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g206 ( 
.A(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_121),
.B(n_142),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_189),
.Y(n_256)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_210),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_212),
.Y(n_253)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_164),
.A2(n_159),
.B(n_109),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_106),
.B(n_111),
.C(n_149),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_151),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_214),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_118),
.A2(n_120),
.B1(n_136),
.B2(n_158),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_220),
.A2(n_206),
.B1(n_171),
.B2(n_174),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_227),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_202),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_132),
.B1(n_157),
.B2(n_134),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_236),
.B1(n_238),
.B2(n_244),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_175),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_165),
.A2(n_157),
.B1(n_141),
.B2(n_149),
.Y(n_236)
);

HB1xp67_ASAP7_75t_SL g269 ( 
.A(n_237),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_141),
.B1(n_106),
.B2(n_111),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_256),
.B1(n_235),
.B2(n_250),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_SL g242 ( 
.A1(n_166),
.A2(n_197),
.B(n_207),
.C(n_199),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_242),
.A2(n_256),
.B(n_181),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_177),
.B1(n_180),
.B2(n_175),
.Y(n_244)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_168),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_210),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_170),
.A2(n_213),
.B1(n_216),
.B2(n_186),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_183),
.B1(n_244),
.B2(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_169),
.C(n_185),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_260),
.C(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_167),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_278),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_184),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_268),
.B1(n_273),
.B2(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_271),
.B(n_276),
.Y(n_289)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_267),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_250),
.B1(n_235),
.B2(n_239),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_272),
.B(n_277),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_242),
.A2(n_212),
.B1(n_182),
.B2(n_215),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_209),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_252),
.B(n_179),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_286),
.C(n_260),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_219),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_219),
.B(n_252),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_218),
.C(n_225),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_282),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_248),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_218),
.B(n_234),
.C(n_221),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_246),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_255),
.Y(n_299)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_218),
.B(n_238),
.C(n_243),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_249),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_283),
.Y(n_306)
);

OAI32xp33_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_257),
.A3(n_254),
.B1(n_237),
.B2(n_245),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_302),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_251),
.B(n_240),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_293),
.B(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_305),
.B1(n_270),
.B2(n_264),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_240),
.B(n_227),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_297),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_259),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_299),
.B(n_306),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_276),
.A2(n_229),
.B1(n_245),
.B2(n_231),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_255),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_273),
.A2(n_217),
.B1(n_232),
.B2(n_226),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_308),
.A2(n_280),
.B(n_270),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_275),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_317),
.C(n_292),
.Y(n_329)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_295),
.B(n_279),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_315),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_307),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_326),
.B1(n_302),
.B2(n_304),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_282),
.C(n_274),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_318),
.A2(n_290),
.B(n_293),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g340 ( 
.A1(n_319),
.A2(n_299),
.B(n_288),
.Y(n_340)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_303),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_323),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_294),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_330),
.C(n_332),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_296),
.C(n_291),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_301),
.C(n_294),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_333),
.A2(n_266),
.B(n_325),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_327),
.A2(n_297),
.B1(n_289),
.B2(n_266),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_342),
.B1(n_305),
.B2(n_321),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_289),
.C(n_304),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_326),
.C(n_312),
.Y(n_347)
);

NAND4xp25_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_318),
.C(n_328),
.D(n_323),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_348),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_327),
.B(n_322),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_353),
.B(n_342),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_352),
.C(n_338),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_322),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_349),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_336),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_312),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_332),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_298),
.C(n_324),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_354),
.A2(n_353),
.B(n_346),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_357),
.Y(n_367)
);

XOR2x2_ASAP7_75t_SL g357 ( 
.A(n_347),
.B(n_337),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_345),
.C(n_352),
.Y(n_365)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_361),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_355),
.B(n_351),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_365),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_366),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_341),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_365),
.B(n_358),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_369),
.B(n_371),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_361),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_368),
.A2(n_345),
.B(n_362),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_372),
.A2(n_374),
.B(n_217),
.Y(n_376)
);

AOI32xp33_ASAP7_75t_L g374 ( 
.A1(n_370),
.A2(n_367),
.A3(n_331),
.B1(n_320),
.B2(n_313),
.Y(n_374)
);

AOI322xp5_ASAP7_75t_L g375 ( 
.A1(n_373),
.A2(n_331),
.A3(n_232),
.B1(n_262),
.B2(n_267),
.C1(n_285),
.C2(n_300),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_335),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_226),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_378),
.Y(n_379)
);


endmodule