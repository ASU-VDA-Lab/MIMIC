module fake_jpeg_13442_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_1),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_21),
.B1(n_38),
.B2(n_37),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_67),
.B1(n_40),
.B2(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_41),
.Y(n_68)
);

NAND2x1_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_0),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_18),
.B1(n_36),
.B2(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_79),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_60),
.B1(n_55),
.B2(n_58),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_70),
.B1(n_78),
.B2(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_57),
.B1(n_50),
.B2(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_75),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_81),
.B(n_41),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_50),
.B1(n_42),
.B2(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_75),
.B1(n_74),
.B2(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_90),
.B1(n_11),
.B2(n_12),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_66),
.C(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_46),
.B1(n_52),
.B2(n_48),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_89),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_10),
.Y(n_112)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_45),
.B1(n_44),
.B2(n_63),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_52),
.B1(n_48),
.B2(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_46),
.C(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_22),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_39),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_107),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_105),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_2),
.A3(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_14),
.B(n_16),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_8),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_109),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_9),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_10),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_100),
.B(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_33),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_14),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_97),
.B1(n_87),
.B2(n_26),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_121),
.B1(n_113),
.B2(n_108),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g121 ( 
.A1(n_115),
.A2(n_23),
.B(n_29),
.C(n_28),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_104),
.B1(n_103),
.B2(n_114),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.C(n_130),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_24),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

OAI322xp33_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_122),
.A3(n_116),
.B1(n_127),
.B2(n_119),
.C1(n_126),
.C2(n_121),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_119),
.B1(n_133),
.B2(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_124),
.B(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_118),
.Y(n_141)
);


endmodule