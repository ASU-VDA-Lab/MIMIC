module real_jpeg_32369_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_0),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_0),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_1),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_1),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_1),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_1),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_1),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_2),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_2),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_2),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_2),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_2),
.B(n_109),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_2),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_2),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_3),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_3),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_3),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_3),
.B(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_6),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_6),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_6),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_6),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g326 ( 
.A(n_6),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_6),
.B(n_341),
.Y(n_340)
);

NAND2x1_ASAP7_75t_L g57 ( 
.A(n_7),
.B(n_58),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_7),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_7),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_9),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_11),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_12),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_12),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_12),
.B(n_218),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_12),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_12),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_12),
.B(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_13),
.Y(n_189)
);

AND2x4_ASAP7_75t_SL g46 ( 
.A(n_14),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_14),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_14),
.B(n_86),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_14),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_14),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_14),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_15),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_15),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_15),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_15),
.B(n_141),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_15),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_15),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_15),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_221),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_220),
.Y(n_17)
);

INVxp67_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_173),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_21),
.B(n_173),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_103),
.C(n_146),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_24),
.A2(n_25),
.B1(n_105),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_77),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_54),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_27),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_41),
.B(n_53),
.Y(n_27)
);

NOR2xp67_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_35),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_29),
.B(n_35),
.Y(n_170)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_33),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_34),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_34),
.Y(n_355)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_40),
.Y(n_256)
);

XNOR2x2_ASAP7_75t_L g169 ( 
.A(n_41),
.B(n_170),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.C(n_49),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_42),
.A2(n_43),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_42),
.A2(n_43),
.B1(n_49),
.B2(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_45),
.B(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_47),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_48),
.Y(n_332)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_49),
.Y(n_262)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_52),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_76),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_57),
.Y(n_64)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_61),
.B(n_64),
.C(n_76),
.Y(n_193)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_63),
.Y(n_244)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.C(n_73),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_73),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_70),
.B(n_202),
.Y(n_269)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.C(n_87),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_78),
.B(n_80),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_80),
.A2(n_81),
.B(n_85),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_87),
.B(n_382),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.C(n_99),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_88),
.A2(n_89),
.B1(n_99),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_94),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_95),
.B(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_98),
.Y(n_219)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_102),
.Y(n_305)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_105),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_122),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_181),
.C(n_182),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_108),
.B(n_116),
.C(n_120),
.Y(n_192)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_113),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_115),
.Y(n_240)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_135),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_123),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_131),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_128),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_135),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_136),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_136),
.A2(n_137),
.B1(n_274),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_198),
.B(n_205),
.Y(n_197)
);

OAI221xp5_ASAP7_75t_L g205 ( 
.A1(n_137),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_137),
.B(n_142),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_137),
.B(n_142),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_145),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_139),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_142),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_142),
.A2(n_145),
.B1(n_155),
.B2(n_156),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_143),
.Y(n_341)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_147),
.B(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_169),
.C(n_171),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_148),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_159),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_149),
.A2(n_150),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_153),
.A2(n_154),
.B1(n_159),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_167),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_160),
.B(n_167),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_162),
.B(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_163),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_168),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_169),
.B(n_171),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_196),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_187),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_193),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_206),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_198)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_209),
.A2(n_250),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_385),
.B(n_391),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_374),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_283),
.B(n_373),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_263),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_225),
.B(n_263),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_227),
.B(n_246),
.C(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.Y(n_231)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_232),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_245),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_245),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.C(n_242),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_237),
.B(n_243),
.Y(n_316)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_241),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_260),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_248),
.B(n_260),
.C(n_384),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_249),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.C(n_257),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_258),
.Y(n_266)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_268),
.B(n_277),
.C(n_280),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_264),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_265),
.A2(n_268),
.B1(n_281),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_265),
.Y(n_371)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.C(n_273),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_277),
.A2(n_278),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_365),
.B(n_372),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_322),
.B(n_364),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_312),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_286),
.B(n_312),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_302),
.C(n_309),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_287),
.A2(n_288),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_295),
.C(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_302),
.A2(n_309),
.B1(n_310),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_306),
.Y(n_325)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx4f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_319),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_315),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_317),
.C(n_367),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_337),
.B(n_363),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_333),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_333),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.C(n_329),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_326),
.A2(n_329),
.B1(n_330),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_326),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_350),
.B(n_362),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_347),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_339),
.B(n_347),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_342),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_340),
.B(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_357),
.B(n_361),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_356),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_356),
.Y(n_361)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_368),
.Y(n_372)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_377),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_381),
.C(n_383),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21x1_ASAP7_75t_L g392 ( 
.A1(n_386),
.A2(n_393),
.B(n_394),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_388),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);


endmodule