module fake_jpeg_1896_n_98 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_41),
.B1(n_39),
.B2(n_35),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_49),
.Y(n_53)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_28),
.B1(n_32),
.B2(n_30),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_1),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_50),
.B1(n_49),
.B2(n_34),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_65),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_50),
.B1(n_34),
.B2(n_43),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_58),
.B1(n_43),
.B2(n_5),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_43),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_75),
.B(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_74),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_13),
.B1(n_23),
.B2(n_22),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_3),
.B(n_4),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_5),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_14),
.C(n_21),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_65),
.C(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_87),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_12),
.C(n_20),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_75),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_6),
.B(n_7),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_81),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_88),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_90),
.Y(n_93)
);

OAI221xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_89),
.B1(n_84),
.B2(n_83),
.C(n_11),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_9),
.C(n_15),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_17),
.C(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_24),
.B1(n_7),
.B2(n_8),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_8),
.Y(n_98)
);


endmodule