module fake_jpeg_10281_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_34),
.Y(n_43)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_0),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_20),
.B2(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_21),
.B1(n_20),
.B2(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_50),
.B1(n_37),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_31),
.B1(n_37),
.B2(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_24),
.B1(n_22),
.B2(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_63),
.B1(n_66),
.B2(n_17),
.Y(n_81)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_34),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_27),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_14),
.B(n_15),
.C(n_23),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_33),
.B1(n_32),
.B2(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_13),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_81),
.B1(n_56),
.B2(n_66),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_14),
.B(n_23),
.C(n_15),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_29),
.B1(n_36),
.B2(n_28),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_22),
.B1(n_53),
.B2(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_29),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_90),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_44),
.B(n_17),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_70),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_75),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_71),
.B1(n_73),
.B2(n_6),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_6),
.C(n_2),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_12),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_83),
.B(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_82),
.B1(n_75),
.B2(n_73),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_87),
.C(n_90),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_116),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_107),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_117),
.Y(n_119)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_99),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_100),
.B1(n_111),
.B2(n_112),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_101),
.B1(n_95),
.B2(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_110),
.C(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.C(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_119),
.B1(n_121),
.B2(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_131),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_7),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_91),
.B1(n_97),
.B2(n_102),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_3),
.B(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_9),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_132),
.B(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_137),
.B(n_135),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_10),
.Y(n_139)
);


endmodule