module fake_jpeg_24704_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_225;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_23),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_56),
.Y(n_103)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_23),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_5),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_73),
.Y(n_99)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_16),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_25),
.B1(n_29),
.B2(n_19),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_79),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_30),
.B1(n_33),
.B2(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_28),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_69),
.B1(n_77),
.B2(n_12),
.Y(n_113)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_109),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_22),
.B(n_21),
.C(n_19),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_104),
.B(n_73),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_34),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_70),
.B(n_55),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_15),
.B(n_13),
.C(n_76),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_6),
.B(n_7),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_107),
.B1(n_63),
.B2(n_71),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_54),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_105),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_123),
.B(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_121),
.B1(n_82),
.B2(n_100),
.Y(n_147)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_129),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_65),
.B1(n_79),
.B2(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_130),
.B1(n_97),
.B2(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_125),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_92),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_65),
.B1(n_78),
.B2(n_60),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g154 ( 
.A(n_122),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_76),
.B(n_57),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_57),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_15),
.B1(n_103),
.B2(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_134),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_87),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_145),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_99),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_115),
.B1(n_128),
.B2(n_123),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_151),
.B(n_158),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_R g151 ( 
.A(n_120),
.B(n_93),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_117),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_87),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_127),
.B(n_104),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_116),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_82),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_82),
.B(n_88),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_113),
.B(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_98),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_173),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_171),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_174),
.B(n_176),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_177),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_132),
.B(n_113),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_114),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_95),
.C(n_112),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_176),
.C(n_172),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_191),
.C(n_164),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_180),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_186),
.B(n_139),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_194),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_164),
.A3(n_156),
.B1(n_174),
.B2(n_158),
.C1(n_168),
.C2(n_145),
.Y(n_190)
);

OA21x2_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_140),
.B(n_141),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_181),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_155),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g196 ( 
.A(n_169),
.B(n_163),
.C(n_150),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_147),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_142),
.B1(n_158),
.B2(n_160),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_141),
.B1(n_162),
.B2(n_148),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_175),
.B1(n_153),
.B2(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_208),
.C(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_201),
.B(n_148),
.Y(n_216)
);

NAND2xp67_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_157),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_188),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_197),
.B1(n_192),
.B2(n_154),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_193),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_178),
.B1(n_171),
.B2(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_194),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_180),
.C(n_161),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_183),
.C(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_192),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_214),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_220),
.B(n_202),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_205),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_185),
.C(n_193),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_203),
.B(n_211),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_202),
.B(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_215),
.C(n_220),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_182),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_209),
.B1(n_204),
.B2(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_233),
.A2(n_204),
.B1(n_227),
.B2(n_144),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_204),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_228),
.C(n_154),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_234),
.C(n_144),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_182),
.B(n_129),
.Y(n_240)
);


endmodule