module real_jpeg_105_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_6),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_18),
.C(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_29),
.B1(n_67),
.B2(n_68),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_6),
.B(n_20),
.C(n_46),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_35),
.C(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_39),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_6),
.B(n_54),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_82),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_80),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_60),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_12),
.B(n_60),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_48),
.C(n_52),
.Y(n_12)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_13),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_15),
.B1(n_30),
.B2(n_31),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_15),
.B1(n_52),
.B2(n_53),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_14),
.A2(n_53),
.B(n_110),
.C(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_32),
.C(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_15),
.B(n_52),
.Y(n_114)
);

AO21x2_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_24),
.B(n_28),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_24),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_17)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

OA22x2_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_19),
.A2(n_20),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_51),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_25),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_25),
.B(n_89),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_31)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_32),
.A2(n_47),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_32),
.A2(n_47),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_32),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_32),
.B(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_32),
.B(n_52),
.C(n_94),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_32),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_39),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_35),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_35),
.B(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AO21x2_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_65),
.B(n_70),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_46),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_53),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_53),
.B1(n_87),
.B2(n_88),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_87),
.Y(n_86)
);

OA21x2_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B(n_59),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_58),
.Y(n_57)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_73),
.B2(n_74),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_71),
.B2(n_72),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_79),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_72),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_112),
.B(n_118),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_106),
.B(n_111),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_96),
.B(n_105),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_115),
.Y(n_118)
);


endmodule