module fake_jpeg_23164_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_0),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_33),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_65),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_30),
.B(n_28),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_49),
.B(n_50),
.Y(n_99)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_71),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_26),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_38),
.B1(n_17),
.B2(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_19),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_9),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_94),
.Y(n_137)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_83),
.B(n_91),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_90),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_93),
.A2(n_46),
.B1(n_37),
.B2(n_44),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_114),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_102),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_18),
.B(n_22),
.C(n_34),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_19),
.B(n_21),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_20),
.B(n_31),
.Y(n_123)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_19),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_77),
.B1(n_25),
.B2(n_32),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_44),
.C(n_40),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_44),
.C(n_46),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_20),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_46),
.B(n_45),
.C(n_43),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_32),
.B1(n_37),
.B2(n_43),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_126),
.Y(n_155)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_148),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_25),
.B(n_24),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_127),
.A2(n_130),
.B(n_134),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_23),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_26),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_112),
.C(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_145),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_110),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_17),
.B1(n_45),
.B2(n_43),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_106),
.B1(n_102),
.B2(n_84),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_103),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_161),
.B1(n_167),
.B2(n_175),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_99),
.B1(n_89),
.B2(n_98),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_92),
.C(n_97),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_164),
.C(n_22),
.Y(n_211)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_156),
.B(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_84),
.Y(n_158)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_103),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_177),
.B(n_120),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_109),
.B1(n_106),
.B2(n_91),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_165),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_133),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_163),
.A2(n_176),
.B1(n_1),
.B2(n_3),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_92),
.C(n_104),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_109),
.B1(n_116),
.B2(n_111),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_109),
.B(n_37),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_120),
.B(n_140),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_170),
.Y(n_190)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_184),
.B1(n_128),
.B2(n_34),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_27),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_179),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_32),
.B1(n_108),
.B2(n_81),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_133),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_34),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_83),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_183),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_27),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_141),
.A2(n_86),
.B1(n_31),
.B2(n_28),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_168),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_123),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_12),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_121),
.B(n_143),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_198),
.B(n_208),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_121),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_192),
.B(n_11),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_201),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_197),
.B(n_175),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_196),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_149),
.B(n_138),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_182),
.A2(n_124),
.B1(n_122),
.B2(n_128),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_207),
.B1(n_216),
.B2(n_184),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_108),
.B1(n_124),
.B2(n_32),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_202),
.B1(n_152),
.B2(n_170),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_11),
.C(n_15),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_23),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_211),
.C(n_218),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_34),
.B1(n_22),
.B2(n_4),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_160),
.B(n_151),
.Y(n_208)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_176),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_22),
.B1(n_9),
.B2(n_10),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_1),
.C(n_3),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_222),
.A2(n_240),
.B1(n_241),
.B2(n_204),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_193),
.A2(n_157),
.B(n_153),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_155),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_155),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_227),
.B(n_208),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_244),
.B1(n_210),
.B2(n_196),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_232),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_154),
.Y(n_233)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_193),
.B1(n_172),
.B2(n_189),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_243),
.B1(n_202),
.B2(n_200),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_156),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_159),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_192),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_180),
.B1(n_4),
.B2(n_5),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_195),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_1),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_245),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_218),
.C(n_205),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_262),
.B(n_232),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_266),
.B1(n_270),
.B2(n_220),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_252),
.B(n_259),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_185),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_226),
.B(n_230),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_203),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_211),
.B1(n_188),
.B2(n_191),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_264),
.B1(n_267),
.B2(n_220),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_194),
.B1(n_215),
.B2(n_187),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_234),
.A2(n_214),
.B1(n_6),
.B2(n_5),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_214),
.B1(n_6),
.B2(n_8),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_6),
.C(n_7),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_245),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_221),
.B(n_7),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_223),
.Y(n_280)
);

OAI31xp33_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_221),
.A3(n_222),
.B(n_224),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_277),
.B(n_279),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_238),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_261),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_224),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_288),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_244),
.B1(n_235),
.B2(n_239),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_264),
.C(n_247),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_219),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_256),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_263),
.C(n_255),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_304),
.C(n_295),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_257),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_305),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

OR2x6_ASAP7_75t_SL g323 ( 
.A(n_308),
.B(n_248),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_309),
.B(n_313),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_276),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_312),
.B(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_273),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_283),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_302),
.Y(n_327)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_318),
.B(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_229),
.Y(n_319)
);

XOR2x1_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_272),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_324),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_326),
.B(n_315),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_303),
.Y(n_324)
);

AOI21x1_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_255),
.B(n_299),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_325),
.A2(n_286),
.B(n_268),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_305),
.C(n_298),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_307),
.A2(n_282),
.B1(n_271),
.B2(n_275),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_316),
.C(n_289),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_243),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_335),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_329),
.B(n_321),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_337),
.A2(n_340),
.B(n_339),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_291),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_336),
.B1(n_329),
.B2(n_333),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_342),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_313),
.C(n_291),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_246),
.C(n_225),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_286),
.B(n_280),
.C(n_15),
.D(n_13),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_12),
.Y(n_347)
);


endmodule