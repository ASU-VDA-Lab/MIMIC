module fake_jpeg_30699_n_287 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_287);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_15),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_49),
.A2(n_51),
.B1(n_93),
.B2(n_17),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_26),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_36),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_32),
.B(n_35),
.C(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_61),
.Y(n_101)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_65),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_78),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_33),
.B1(n_26),
.B2(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_104)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_76),
.Y(n_119)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_27),
.Y(n_80)
);

NAND2x1_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_30),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_95),
.C(n_28),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_85),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_89),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_39),
.A2(n_33),
.B1(n_28),
.B2(n_23),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_88),
.B1(n_1),
.B2(n_3),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_39),
.A2(n_28),
.B1(n_17),
.B2(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_37),
.A2(n_31),
.B(n_35),
.C(n_22),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_94),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_40),
.B(n_22),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_37),
.B(n_34),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_37),
.A2(n_30),
.B(n_8),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_98),
.B(n_105),
.CI(n_115),
.CON(n_145),
.SN(n_145)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_107),
.B1(n_114),
.B2(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_30),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_69),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_55),
.B(n_77),
.C(n_82),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_96),
.B1(n_117),
.B2(n_78),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_7),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_115),
.B1(n_14),
.B2(n_1),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_49),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_88),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_103),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_129),
.A2(n_141),
.B1(n_149),
.B2(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_131),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_69),
.C(n_53),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_73),
.B1(n_79),
.B2(n_52),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_69),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_13),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_71),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_116),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_146),
.A2(n_104),
.B1(n_119),
.B2(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_52),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_62),
.B1(n_82),
.B2(n_68),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_99),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_155),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_62),
.B(n_55),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_156),
.B(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_63),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_158),
.Y(n_172)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_112),
.A2(n_63),
.B1(n_77),
.B2(n_76),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_113),
.B(n_14),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_174),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_178),
.B(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_126),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_142),
.B1(n_132),
.B2(n_146),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_145),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_112),
.B(n_110),
.C(n_120),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_124),
.B(n_97),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_189),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_134),
.B(n_116),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_188),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_136),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_121),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_190),
.B(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_206),
.B1(n_208),
.B2(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_187),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_196),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_130),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_164),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_149),
.B1(n_131),
.B2(n_158),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_141),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_209),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_129),
.B1(n_131),
.B2(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_143),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_210),
.A2(n_211),
.B1(n_183),
.B2(n_133),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_171),
.B(n_161),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_166),
.B(n_174),
.Y(n_213)
);

OAI321xp33_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_172),
.A3(n_177),
.B1(n_187),
.B2(n_160),
.C(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_231),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_171),
.B1(n_161),
.B2(n_176),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_212),
.B1(n_211),
.B2(n_210),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_228),
.B1(n_196),
.B2(n_191),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_188),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_165),
.B1(n_176),
.B2(n_168),
.Y(n_228)
);

OAI321xp33_ASAP7_75t_L g230 ( 
.A1(n_197),
.A2(n_178),
.A3(n_186),
.B1(n_170),
.B2(n_182),
.C(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_169),
.C(n_152),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_203),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_234),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_222),
.B(n_209),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_243),
.C(n_231),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_228),
.Y(n_248)
);

FAx1_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_199),
.CI(n_213),
.CON(n_239),
.SN(n_239)
);

NOR3xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_221),
.C(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_208),
.B1(n_196),
.B2(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_241),
.B1(n_245),
.B2(n_230),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_204),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_207),
.B1(n_199),
.B2(n_198),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_217),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_240),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_220),
.C(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_251),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_232),
.B(n_216),
.C(n_219),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_256),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_244),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_221),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_215),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_237),
.B(n_236),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_241),
.B(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_264),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_237),
.B1(n_238),
.B2(n_242),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_246),
.B(n_245),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_265),
.Y(n_273)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_192),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_251),
.B(n_249),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_271),
.B(n_272),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_169),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_247),
.B(n_194),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_265),
.Y(n_279)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_278),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_264),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_279),
.A2(n_266),
.B(n_270),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_281),
.B(n_195),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_276),
.A2(n_277),
.B(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_260),
.C(n_184),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.C(n_205),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_285),
.A2(n_184),
.B(n_154),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_121),
.Y(n_287)
);


endmodule