module fake_jpeg_10142_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_18),
.B1(n_29),
.B2(n_27),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_27),
.C(n_18),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_21),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_22),
.B1(n_21),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_17),
.B1(n_23),
.B2(n_32),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_66),
.B1(n_23),
.B2(n_32),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_0),
.Y(n_62)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_51),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_32),
.B1(n_23),
.B2(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_68),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_64),
.B1(n_51),
.B2(n_60),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_85),
.B(n_86),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_78),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_33),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_62),
.C(n_47),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_25),
.Y(n_130)
);

CKINVDCx11_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_103),
.Y(n_114)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_53),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_105),
.B(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_56),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_69),
.A2(n_49),
.B(n_60),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_51),
.B1(n_64),
.B2(n_89),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_15),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_14),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_62),
.Y(n_108)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_84),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_74),
.B1(n_67),
.B2(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_131),
.B(n_63),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_78),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_107),
.C(n_28),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_64),
.B1(n_82),
.B2(n_87),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_63),
.B1(n_48),
.B2(n_58),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_99),
.B1(n_28),
.B2(n_95),
.Y(n_154)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_90),
.B1(n_109),
.B2(n_63),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_102),
.C(n_93),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_135),
.C(n_138),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_100),
.C(n_91),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_91),
.B1(n_100),
.B2(n_108),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_131),
.B1(n_120),
.B2(n_112),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_108),
.C(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_153),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_152),
.B(n_153),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_95),
.B(n_28),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_125),
.B1(n_131),
.B2(n_132),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_154),
.B1(n_126),
.B2(n_95),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_33),
.B(n_28),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_43),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_33),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_38),
.C(n_43),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_163),
.B1(n_167),
.B2(n_166),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_162),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_157),
.B(n_170),
.Y(n_178)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_164),
.Y(n_188)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_133),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_158),
.C(n_160),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_171),
.A2(n_172),
.B1(n_111),
.B2(n_6),
.Y(n_187)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_172),
.A2(n_136),
.B1(n_138),
.B2(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_187),
.B1(n_182),
.B2(n_185),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_179),
.B1(n_183),
.B2(n_155),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_134),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_177),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_151),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_180),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_150),
.B(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_126),
.C(n_111),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_3),
.B(n_4),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_5),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_166),
.B1(n_165),
.B2(n_171),
.Y(n_183)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_199),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_196),
.B(n_177),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_164),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_176),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_204),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_178),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_179),
.CI(n_174),
.CON(n_205),
.SN(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_200),
.B(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_207),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_206),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_190),
.B(n_194),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_215),
.A2(n_181),
.B(n_155),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_193),
.B(n_194),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_205),
.B1(n_209),
.B2(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_219),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_211),
.A2(n_215),
.B1(n_213),
.B2(n_111),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_220),
.A2(n_11),
.B(n_13),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

AO221x1_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_224),
.B(n_6),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_225),
.C(n_221),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_229),
.C(n_8),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_226),
.A2(n_223),
.B(n_218),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_230),
.B(n_9),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_10),
.Y(n_232)
);


endmodule