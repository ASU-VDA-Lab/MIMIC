module fake_jpeg_28479_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_5),
.Y(n_8)
);

HAxp5_ASAP7_75t_SL g9 ( 
.A(n_0),
.B(n_3),
.CON(n_9),
.SN(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_2),
.Y(n_12)
);

A2O1A1Ixp33_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_16),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_10),
.A2(n_11),
.B1(n_6),
.B2(n_7),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_23)
);

CKINVDCx12_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_6),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

XOR2x2_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_18),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_25),
.C(n_22),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_20),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_31),
.C(n_32),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_23),
.Y(n_31)
);

AOI31xp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_28),
.A3(n_29),
.B(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_33),
.B(n_28),
.Y(n_36)
);

AOI321xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_29),
.A3(n_21),
.B1(n_8),
.B2(n_24),
.C(n_19),
.Y(n_37)
);


endmodule