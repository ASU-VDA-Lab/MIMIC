module fake_jpeg_25586_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_31),
.Y(n_52)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_56),
.C(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_30),
.B1(n_17),
.B2(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_42),
.B1(n_35),
.B2(n_30),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_33),
.C(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_62),
.B1(n_85),
.B2(n_88),
.Y(n_94)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_30),
.B1(n_17),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_42),
.B1(n_38),
.B2(n_35),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_89),
.B1(n_57),
.B2(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_67),
.Y(n_90)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_75),
.Y(n_95)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_79),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_29),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_40),
.B1(n_35),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_16),
.B1(n_24),
.B2(n_19),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_17),
.B1(n_20),
.B2(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_45),
.A2(n_20),
.B1(n_27),
.B2(n_41),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_20),
.B1(n_27),
.B2(n_41),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_92),
.A2(n_98),
.B1(n_83),
.B2(n_79),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_32),
.B1(n_29),
.B2(n_22),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_56),
.B1(n_57),
.B2(n_39),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_32),
.B1(n_29),
.B2(n_21),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_105),
.B1(n_24),
.B2(n_19),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_39),
.C(n_37),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_104),
.C(n_81),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_58),
.B1(n_66),
.B2(n_21),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_61),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_144),
.C(n_36),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_134),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_124),
.B1(n_145),
.B2(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_65),
.B1(n_71),
.B2(n_83),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_65),
.B(n_1),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_142),
.B(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_132),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_95),
.B1(n_117),
.B2(n_115),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_33),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_28),
.Y(n_134)
);

XOR2x2_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_33),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_16),
.B(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_109),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_82),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_19),
.B(n_24),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_22),
.B(n_25),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_103),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_39),
.B1(n_37),
.B2(n_36),
.Y(n_145)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_155),
.B1(n_160),
.B2(n_113),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_153),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_110),
.B(n_108),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_167),
.B(n_169),
.Y(n_188)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_109),
.B(n_95),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_156),
.A2(n_175),
.B1(n_26),
.B2(n_1),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_129),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_166),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_95),
.B1(n_111),
.B2(n_102),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_174),
.B1(n_119),
.B2(n_121),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_93),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_165),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_127),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_172),
.B(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_37),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_123),
.A2(n_111),
.B1(n_102),
.B2(n_110),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_93),
.B1(n_113),
.B2(n_108),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_186),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_179),
.A2(n_183),
.B1(n_192),
.B2(n_195),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_157),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_142),
.B(n_143),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_0),
.B(n_3),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_75),
.B1(n_37),
.B2(n_25),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_18),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_185),
.C(n_187),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_172),
.C(n_151),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_146),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_18),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_26),
.C(n_18),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_194),
.C(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_193),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_26),
.B1(n_9),
.B2(n_10),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_26),
.C(n_9),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_26),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_26),
.C(n_9),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_168),
.C(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_152),
.A2(n_8),
.B1(n_14),
.B2(n_12),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_150),
.B1(n_162),
.B2(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_171),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_155),
.B1(n_158),
.B2(n_156),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_205),
.A2(n_217),
.B1(n_192),
.B2(n_193),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_220),
.Y(n_234)
);

OA21x2_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_155),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_155),
.C(n_173),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_0),
.C(n_3),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_194),
.B1(n_198),
.B2(n_12),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_179),
.A2(n_150),
.B1(n_1),
.B2(n_2),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_10),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_178),
.B(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_8),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_182),
.B(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_226),
.A2(n_221),
.B(n_217),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_197),
.B1(n_182),
.B2(n_181),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_223),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_196),
.B1(n_185),
.B2(n_183),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_190),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_240),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_15),
.B1(n_5),
.B2(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_5),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_208),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_209),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_245),
.Y(n_257)
);

AND2x4_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_206),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_252),
.Y(n_263)
);

XOR2x2_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_205),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_248),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_222),
.B(n_205),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_204),
.C(n_207),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_255),
.C(n_213),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_207),
.C(n_208),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_262),
.C(n_265),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_225),
.C(n_231),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_231),
.C(n_235),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_219),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_259),
.A2(n_247),
.B1(n_250),
.B2(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_248),
.B1(n_243),
.B2(n_224),
.Y(n_268)
);

OAI321xp33_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_271),
.A3(n_269),
.B1(n_263),
.B2(n_258),
.C(n_239),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_246),
.B(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_257),
.A2(n_246),
.B(n_233),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_274),
.C(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_264),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_251),
.C(n_255),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_254),
.B1(n_232),
.B2(n_216),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_261),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_264),
.B(n_272),
.C(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_282),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_260),
.C(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_283),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_15),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_287),
.A2(n_278),
.B(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_290),
.Y(n_291)
);

OAI21x1_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_286),
.B(n_285),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_0),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_291),
.B(n_4),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_4),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_4),
.B(n_209),
.Y(n_297)
);


endmodule