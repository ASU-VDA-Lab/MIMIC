module fake_jpeg_29652_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_34),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_38),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_54),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_43),
.C(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_45),
.Y(n_66)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_16),
.B1(n_32),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_57),
.B1(n_0),
.B2(n_1),
.Y(n_61)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_56),
.B1(n_47),
.B2(n_4),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_58),
.Y(n_77)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_6),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_40),
.B(n_41),
.C(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_75),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_7),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_18),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_19),
.B1(n_29),
.B2(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_8),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_91),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_6),
.C(n_7),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_76),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_62),
.C(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_95),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_97),
.B1(n_83),
.B2(n_94),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_73),
.C(n_95),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_94),
.B1(n_90),
.B2(n_80),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_86),
.B1(n_10),
.B2(n_9),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_105),
.C(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_11),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_15),
.B(n_17),
.C(n_21),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_23),
.A3(n_25),
.B1(n_26),
.B2(n_27),
.C1(n_33),
.C2(n_100),
.Y(n_115)
);


endmodule