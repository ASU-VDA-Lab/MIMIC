module real_aes_8669_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g444 ( .A(n_0), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_1), .A2(n_149), .B(n_152), .C(n_232), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_2), .A2(n_178), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g510 ( .A(n_3), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_4), .B(n_208), .Y(n_207) );
AOI21xp33_ASAP7_75t_L g493 ( .A1(n_5), .A2(n_178), .B(n_494), .Y(n_493) );
AND2x6_ASAP7_75t_L g149 ( .A(n_6), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g245 ( .A(n_7), .Y(n_245) );
INVx1_ASAP7_75t_L g108 ( .A(n_8), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_8), .B(n_43), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_9), .A2(n_177), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_10), .B(n_161), .Y(n_234) );
INVx1_ASAP7_75t_L g498 ( .A(n_11), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_12), .B(n_202), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_13), .A2(n_453), .B1(n_454), .B2(n_460), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_13), .Y(n_460) );
INVx1_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
INVx1_ASAP7_75t_L g545 ( .A(n_15), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_16), .A2(n_81), .B1(n_458), .B2(n_459), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_16), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_17), .A2(n_186), .B(n_267), .C(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_18), .B(n_208), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_19), .B(n_476), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_20), .B(n_178), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_21), .B(n_192), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_22), .A2(n_202), .B(n_253), .C(n_255), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_23), .B(n_208), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_24), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_25), .A2(n_188), .B(n_269), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_26), .B(n_161), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g143 ( .A(n_27), .Y(n_143) );
INVx1_ASAP7_75t_L g215 ( .A(n_28), .Y(n_215) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_29), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_30), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_31), .B(n_161), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_32), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g184 ( .A(n_33), .Y(n_184) );
INVx1_ASAP7_75t_L g488 ( .A(n_34), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_35), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_35), .Y(n_455) );
INVx2_ASAP7_75t_L g147 ( .A(n_36), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_37), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_38), .A2(n_202), .B(n_203), .C(n_205), .Y(n_201) );
INVxp67_ASAP7_75t_L g187 ( .A(n_39), .Y(n_187) );
CKINVDCx14_ASAP7_75t_R g200 ( .A(n_40), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_41), .A2(n_152), .B(n_214), .C(n_218), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_42), .A2(n_149), .B(n_152), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_43), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g487 ( .A(n_44), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_45), .A2(n_163), .B(n_243), .C(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_46), .B(n_161), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_47), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_48), .Y(n_180) );
INVx1_ASAP7_75t_L g251 ( .A(n_49), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_50), .Y(n_489) );
AOI222xp33_ASAP7_75t_SL g450 ( .A1(n_51), .A2(n_451), .B1(n_452), .B2(n_461), .C1(n_747), .C2(n_750), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g432 ( .A1(n_52), .A2(n_61), .B1(n_433), .B2(n_434), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_52), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_53), .B(n_178), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_54), .A2(n_152), .B1(n_255), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_55), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_56), .Y(n_507) );
CKINVDCx14_ASAP7_75t_R g241 ( .A(n_57), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_58), .A2(n_205), .B(n_243), .C(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_59), .A2(n_123), .B1(n_124), .B2(n_437), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_59), .Y(n_437) );
INVx1_ASAP7_75t_L g495 ( .A(n_60), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_61), .Y(n_434) );
INVx1_ASAP7_75t_L g150 ( .A(n_62), .Y(n_150) );
INVx1_ASAP7_75t_L g140 ( .A(n_63), .Y(n_140) );
INVx1_ASAP7_75t_SL g204 ( .A(n_64), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_66), .A2(n_432), .B1(n_435), .B2(n_436), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_66), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_67), .B(n_208), .Y(n_257) );
INVx1_ASAP7_75t_L g156 ( .A(n_68), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_SL g475 ( .A1(n_69), .A2(n_205), .B(n_476), .C(n_477), .Y(n_475) );
INVxp67_ASAP7_75t_L g478 ( .A(n_70), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_71), .A2(n_105), .B1(n_115), .B2(n_754), .Y(n_104) );
INVx1_ASAP7_75t_L g114 ( .A(n_72), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_73), .A2(n_178), .B(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_74), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_75), .A2(n_178), .B(n_264), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_76), .Y(n_491) );
INVx1_ASAP7_75t_L g551 ( .A(n_77), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_78), .A2(n_177), .B(n_179), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g212 ( .A(n_79), .Y(n_212) );
INVx1_ASAP7_75t_L g265 ( .A(n_80), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_81), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_82), .A2(n_149), .B(n_152), .C(n_553), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_83), .A2(n_178), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g268 ( .A(n_84), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_85), .B(n_185), .Y(n_522) );
INVx2_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
INVx1_ASAP7_75t_L g233 ( .A(n_87), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_88), .B(n_476), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_89), .A2(n_149), .B(n_152), .C(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g111 ( .A(n_90), .Y(n_111) );
OR2x2_ASAP7_75t_L g441 ( .A(n_90), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g462 ( .A(n_90), .B(n_443), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_91), .A2(n_152), .B(n_155), .C(n_165), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_92), .B(n_170), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_93), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_94), .A2(n_149), .B(n_152), .C(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_95), .Y(n_537) );
INVx1_ASAP7_75t_L g474 ( .A(n_96), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_97), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_98), .B(n_185), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_99), .B(n_136), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_100), .B(n_136), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_101), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g254 ( .A(n_102), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_103), .A2(n_178), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g754 ( .A(n_105), .Y(n_754) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g746 ( .A(n_111), .B(n_443), .Y(n_746) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_111), .B(n_442), .Y(n_749) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_449), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g753 ( .A(n_119), .Y(n_753) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_438), .B(n_446), .Y(n_121) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_431), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_125), .A2(n_462), .B1(n_463), .B2(n_744), .Y(n_461) );
INVx2_ASAP7_75t_L g751 ( .A(n_125), .Y(n_751) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_365), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_294), .C(n_324), .D(n_345), .E(n_351), .Y(n_126) );
AOI221xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_224), .B1(n_258), .B2(n_260), .C(n_271), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_221), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_193), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_SL g345 ( .A1(n_132), .A2(n_209), .B(n_346), .C(n_349), .Y(n_345) );
AND2x2_ASAP7_75t_L g415 ( .A(n_132), .B(n_210), .Y(n_415) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_171), .Y(n_132) );
AND2x2_ASAP7_75t_L g273 ( .A(n_133), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g277 ( .A(n_133), .B(n_274), .Y(n_277) );
OR2x2_ASAP7_75t_L g303 ( .A(n_133), .B(n_210), .Y(n_303) );
AND2x2_ASAP7_75t_L g305 ( .A(n_133), .B(n_196), .Y(n_305) );
AND2x2_ASAP7_75t_L g323 ( .A(n_133), .B(n_195), .Y(n_323) );
INVx1_ASAP7_75t_L g356 ( .A(n_133), .Y(n_356) );
INVx2_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_L g223 ( .A(n_134), .Y(n_223) );
AND2x2_ASAP7_75t_L g259 ( .A(n_134), .B(n_196), .Y(n_259) );
AND2x2_ASAP7_75t_L g412 ( .A(n_134), .B(n_210), .Y(n_412) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_167), .Y(n_134) );
INVx3_ASAP7_75t_L g208 ( .A(n_135), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_135), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_135), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_SL g524 ( .A(n_135), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_136), .A2(n_472), .B(n_479), .Y(n_471) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_138), .B(n_139), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_151), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_144), .A2(n_170), .B(n_212), .C(n_213), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_144), .A2(n_230), .B(n_231), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_144), .A2(n_166), .B1(n_485), .B2(n_489), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_144), .A2(n_507), .B(n_508), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_144), .A2(n_551), .B(n_552), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
AND2x4_ASAP7_75t_L g178 ( .A(n_145), .B(n_149), .Y(n_178) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g256 ( .A(n_147), .Y(n_256) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
INVx3_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g476 ( .A(n_148), .Y(n_476) );
INVx4_ASAP7_75t_SL g166 ( .A(n_149), .Y(n_166) );
BUFx3_ASAP7_75t_L g218 ( .A(n_149), .Y(n_218) );
INVx5_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx3_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_153), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_160), .C(n_162), .Y(n_155) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_157), .A2(n_162), .B(n_233), .C(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g486 ( .A1(n_158), .A2(n_159), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
INVx4_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g243 ( .A(n_161), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_162), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_162), .A2(n_554), .B(n_555), .Y(n_553) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g269 ( .A(n_164), .Y(n_269) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g179 ( .A1(n_166), .A2(n_180), .B(n_181), .C(n_182), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_181), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_SL g240 ( .A1(n_166), .A2(n_181), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_166), .A2(n_181), .B(n_251), .C(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_166), .A2(n_181), .B(n_265), .C(n_266), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_166), .A2(n_181), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_166), .A2(n_181), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_166), .A2(n_181), .B(n_542), .C(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_169), .A2(n_529), .B(n_536), .Y(n_528) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_170), .A2(n_239), .B(n_246), .Y(n_238) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_170), .A2(n_540), .B(n_546), .Y(n_539) );
AND2x2_ASAP7_75t_L g293 ( .A(n_171), .B(n_194), .Y(n_293) );
OR2x2_ASAP7_75t_L g297 ( .A(n_171), .B(n_210), .Y(n_297) );
AND2x2_ASAP7_75t_L g322 ( .A(n_171), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g369 ( .A(n_171), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_171), .B(n_331), .Y(n_417) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_190), .Y(n_171) );
INVx1_ASAP7_75t_L g275 ( .A(n_172), .Y(n_275) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_172), .A2(n_550), .B(n_556), .Y(n_549) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_SL g518 ( .A1(n_173), .A2(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_174), .A2(n_484), .B(n_490), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_174), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_174), .A2(n_506), .B(n_513), .Y(n_505) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_176), .A2(n_191), .B(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_183), .B(n_189), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B1(n_187), .B2(n_188), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_185), .A2(n_215), .B(n_216), .C(n_217), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_185), .A2(n_510), .B(n_511), .C(n_512), .Y(n_509) );
INVx5_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_186), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_186), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_186), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_188), .B(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_188), .B(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_188), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g217 ( .A(n_189), .Y(n_217) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI322xp33_ASAP7_75t_L g418 ( .A1(n_193), .A2(n_354), .A3(n_377), .B1(n_398), .B2(n_419), .C1(n_421), .C2(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_194), .B(n_274), .Y(n_421) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_209), .Y(n_194) );
AND2x2_ASAP7_75t_L g222 ( .A(n_195), .B(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g290 ( .A(n_195), .B(n_210), .Y(n_290) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g331 ( .A(n_196), .B(n_210), .Y(n_331) );
AND2x2_ASAP7_75t_L g375 ( .A(n_196), .B(n_209), .Y(n_375) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_207), .Y(n_196) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_197), .A2(n_249), .B(n_257), .Y(n_248) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_197), .A2(n_263), .B(n_270), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_202), .B(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_206), .Y(n_534) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_208), .A2(n_493), .B(n_499), .Y(n_492) );
AND2x2_ASAP7_75t_L g258 ( .A(n_209), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g276 ( .A(n_209), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_209), .B(n_305), .Y(n_429) );
INVx3_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g221 ( .A(n_210), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_210), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g343 ( .A(n_210), .B(n_274), .Y(n_343) );
AND2x2_ASAP7_75t_L g370 ( .A(n_210), .B(n_305), .Y(n_370) );
OR2x2_ASAP7_75t_L g426 ( .A(n_210), .B(n_277), .Y(n_426) );
OR2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_219), .Y(n_210) );
INVx1_ASAP7_75t_SL g312 ( .A(n_221), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_222), .B(n_343), .Y(n_344) );
AND2x2_ASAP7_75t_L g378 ( .A(n_222), .B(n_368), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_222), .B(n_301), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_222), .B(n_423), .Y(n_422) );
OAI31xp33_ASAP7_75t_L g396 ( .A1(n_224), .A2(n_258), .A3(n_397), .B(n_399), .Y(n_396) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_237), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_225), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g379 ( .A(n_225), .B(n_314), .Y(n_379) );
OR2x2_ASAP7_75t_L g386 ( .A(n_225), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g398 ( .A(n_225), .B(n_287), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g332 ( .A(n_226), .B(n_333), .Y(n_332) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g260 ( .A(n_227), .B(n_261), .Y(n_260) );
INVx4_ASAP7_75t_L g281 ( .A(n_227), .Y(n_281) );
AND2x2_ASAP7_75t_L g318 ( .A(n_227), .B(n_262), .Y(n_318) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_228), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_228), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_228), .B(n_437), .Y(n_556) );
AND2x2_ASAP7_75t_L g317 ( .A(n_237), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g387 ( .A(n_237), .Y(n_387) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_247), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_238), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g287 ( .A(n_238), .B(n_248), .Y(n_287) );
INVx2_ASAP7_75t_L g307 ( .A(n_238), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_238), .B(n_248), .Y(n_321) );
AND2x2_ASAP7_75t_L g328 ( .A(n_238), .B(n_284), .Y(n_328) );
BUFx3_ASAP7_75t_L g338 ( .A(n_238), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_238), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g283 ( .A(n_247), .Y(n_283) );
AND2x2_ASAP7_75t_L g291 ( .A(n_247), .B(n_281), .Y(n_291) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g261 ( .A(n_248), .B(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
INVx2_ASAP7_75t_L g512 ( .A(n_255), .Y(n_512) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_SL g298 ( .A(n_259), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_259), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_259), .B(n_368), .Y(n_389) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_260), .B(n_338), .Y(n_391) );
INVx1_ASAP7_75t_SL g425 ( .A(n_260), .Y(n_425) );
INVx1_ASAP7_75t_SL g333 ( .A(n_261), .Y(n_333) );
INVx1_ASAP7_75t_SL g284 ( .A(n_262), .Y(n_284) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
OR2x2_ASAP7_75t_L g306 ( .A(n_262), .B(n_281), .Y(n_306) );
AND2x2_ASAP7_75t_L g320 ( .A(n_262), .B(n_281), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_262), .B(n_310), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_276), .B(n_278), .C(n_289), .Y(n_271) );
AOI31xp33_ASAP7_75t_L g388 ( .A1(n_272), .A2(n_389), .A3(n_390), .B(n_391), .Y(n_388) );
AND2x2_ASAP7_75t_L g361 ( .A(n_273), .B(n_290), .Y(n_361) );
BUFx3_ASAP7_75t_L g301 ( .A(n_274), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_274), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g337 ( .A(n_274), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_274), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g292 ( .A(n_277), .Y(n_292) );
OAI222xp33_ASAP7_75t_L g401 ( .A1(n_277), .A2(n_402), .B1(n_405), .B2(n_406), .C1(n_407), .C2(n_408), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_285), .Y(n_278) );
INVx1_ASAP7_75t_L g407 ( .A(n_279), .Y(n_407) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_281), .B(n_284), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_281), .B(n_307), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_281), .B(n_282), .Y(n_377) );
INVx1_ASAP7_75t_L g428 ( .A(n_281), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_282), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g430 ( .A(n_282), .Y(n_430) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx2_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
AOI32xp33_ASAP7_75t_L g289 ( .A1(n_285), .A2(n_290), .A3(n_291), .B1(n_292), .B2(n_293), .Y(n_289) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_287), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g364 ( .A(n_287), .Y(n_364) );
OR2x2_ASAP7_75t_L g405 ( .A(n_287), .B(n_306), .Y(n_405) );
INVx1_ASAP7_75t_L g341 ( .A(n_288), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_290), .B(n_301), .Y(n_326) );
INVx3_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
AOI322xp5_ASAP7_75t_L g351 ( .A1(n_290), .A2(n_335), .A3(n_352), .B1(n_354), .B2(n_357), .C1(n_361), .C2(n_362), .Y(n_351) );
AND2x2_ASAP7_75t_L g327 ( .A(n_291), .B(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g404 ( .A(n_291), .Y(n_404) );
A2O1A1O1Ixp25_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_299), .C(n_307), .D(n_308), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_295), .B(n_338), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_297), .A2(n_309), .B1(n_312), .B2(n_313), .C(n_316), .Y(n_308) );
INVx1_ASAP7_75t_SL g423 ( .A(n_297), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_304), .B(n_306), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_301), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_303), .A2(n_387), .B1(n_394), .B2(n_395), .C(n_396), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g424 ( .A1(n_304), .A2(n_425), .B1(n_426), .B2(n_427), .C1(n_429), .C2(n_430), .Y(n_424) );
AND2x2_ASAP7_75t_L g382 ( .A(n_305), .B(n_368), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_305), .A2(n_320), .B(n_367), .Y(n_394) );
INVx1_ASAP7_75t_L g408 ( .A(n_305), .Y(n_408) );
INVx2_ASAP7_75t_SL g311 ( .A(n_306), .Y(n_311) );
AND2x2_ASAP7_75t_L g314 ( .A(n_307), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_SL g348 ( .A(n_310), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_310), .B(n_320), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_311), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_311), .B(n_321), .Y(n_350) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI21xp5_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_319), .B(n_322), .Y(n_316) );
INVx1_ASAP7_75t_SL g334 ( .A(n_318), .Y(n_334) );
AND2x2_ASAP7_75t_L g381 ( .A(n_318), .B(n_364), .Y(n_381) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g420 ( .A(n_320), .B(n_338), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_321), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g406 ( .A(n_322), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_329), .B2(n_336), .C(n_339), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B1(n_334), .B2(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_333), .A2(n_340), .B1(n_342), .B2(n_344), .Y(n_339) );
OR2x2_ASAP7_75t_L g410 ( .A(n_334), .B(n_338), .Y(n_410) );
OR2x2_ASAP7_75t_L g413 ( .A(n_334), .B(n_348), .Y(n_413) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_355), .A2(n_410), .B1(n_411), .B2(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g365 ( .A(n_366), .B(n_380), .C(n_392), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_373), .B2(n_376), .C1(n_378), .C2(n_379), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_368), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g390 ( .A(n_370), .Y(n_390) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_383), .B2(n_385), .C(n_388), .Y(n_380) );
INVx1_ASAP7_75t_L g395 ( .A(n_381), .Y(n_395) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NOR5xp2_ASAP7_75t_L g392 ( .A(n_393), .B(n_401), .C(n_409), .D(n_418), .E(n_424), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_432), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g448 ( .A(n_441), .Y(n_448) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_446), .B(n_450), .C(n_752), .Y(n_449) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_462), .A2(n_464), .B1(n_744), .B2(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_465), .B(n_681), .Y(n_464) );
NOR4xp25_ASAP7_75t_L g465 ( .A(n_466), .B(n_611), .C(n_642), .D(n_661), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_569), .C(n_584), .D(n_602), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_515), .B1(n_547), .B2(n_557), .C1(n_562), .C2(n_564), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_500), .Y(n_468) );
INVx1_ASAP7_75t_L g625 ( .A(n_469), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_480), .Y(n_469) );
AND2x2_ASAP7_75t_L g501 ( .A(n_470), .B(n_492), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_470), .B(n_504), .Y(n_654) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g561 ( .A(n_471), .B(n_482), .Y(n_561) );
AND2x2_ASAP7_75t_L g570 ( .A(n_471), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g596 ( .A(n_471), .Y(n_596) );
AND2x2_ASAP7_75t_L g617 ( .A(n_471), .B(n_482), .Y(n_617) );
BUFx2_ASAP7_75t_L g640 ( .A(n_471), .Y(n_640) );
AND2x2_ASAP7_75t_L g664 ( .A(n_471), .B(n_483), .Y(n_664) );
AND2x2_ASAP7_75t_L g728 ( .A(n_471), .B(n_492), .Y(n_728) );
AND2x2_ASAP7_75t_L g629 ( .A(n_480), .B(n_560), .Y(n_629) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_481), .B(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .Y(n_481) );
OR2x2_ASAP7_75t_L g589 ( .A(n_482), .B(n_505), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_482), .B(n_560), .Y(n_601) );
BUFx2_ASAP7_75t_L g733 ( .A(n_482), .Y(n_733) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g503 ( .A(n_483), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g583 ( .A(n_483), .B(n_505), .Y(n_583) );
AND2x2_ASAP7_75t_L g636 ( .A(n_483), .B(n_492), .Y(n_636) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_483), .Y(n_672) );
AND2x2_ASAP7_75t_L g559 ( .A(n_492), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_SL g571 ( .A(n_492), .Y(n_571) );
INVx2_ASAP7_75t_L g582 ( .A(n_492), .Y(n_582) );
BUFx2_ASAP7_75t_L g606 ( .A(n_492), .Y(n_606) );
AND2x2_ASAP7_75t_SL g663 ( .A(n_492), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AOI332xp33_ASAP7_75t_L g584 ( .A1(n_501), .A2(n_585), .A3(n_589), .B1(n_590), .B2(n_594), .B3(n_597), .C1(n_598), .C2(n_600), .Y(n_584) );
NAND2x1_ASAP7_75t_L g669 ( .A(n_501), .B(n_560), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_501), .B(n_574), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_SL g602 ( .A1(n_502), .A2(n_603), .B(n_606), .C(n_607), .Y(n_602) );
AND2x2_ASAP7_75t_L g741 ( .A(n_502), .B(n_582), .Y(n_741) );
INVx3_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g638 ( .A(n_503), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g643 ( .A(n_503), .B(n_640), .Y(n_643) );
INVx1_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
AND2x2_ASAP7_75t_L g677 ( .A(n_504), .B(n_636), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_504), .B(n_617), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_504), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_504), .B(n_595), .Y(n_703) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g560 ( .A(n_505), .Y(n_560) );
OAI31xp33_ASAP7_75t_L g742 ( .A1(n_515), .A2(n_663), .A3(n_670), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .Y(n_515) );
AND2x2_ASAP7_75t_L g547 ( .A(n_516), .B(n_548), .Y(n_547) );
NAND2x1_ASAP7_75t_SL g565 ( .A(n_516), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_516), .Y(n_652) );
AND2x2_ASAP7_75t_L g657 ( .A(n_516), .B(n_568), .Y(n_657) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_517), .A2(n_570), .B(n_572), .C(n_575), .Y(n_569) );
OR2x2_ASAP7_75t_L g586 ( .A(n_517), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g599 ( .A(n_517), .Y(n_599) );
AND2x2_ASAP7_75t_L g605 ( .A(n_517), .B(n_549), .Y(n_605) );
INVx2_ASAP7_75t_L g623 ( .A(n_517), .Y(n_623) );
AND2x2_ASAP7_75t_L g634 ( .A(n_517), .B(n_588), .Y(n_634) );
AND2x2_ASAP7_75t_L g666 ( .A(n_517), .B(n_624), .Y(n_666) );
AND2x2_ASAP7_75t_L g670 ( .A(n_517), .B(n_593), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_517), .B(n_526), .Y(n_675) );
AND2x2_ASAP7_75t_L g709 ( .A(n_517), .B(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_517), .B(n_612), .Y(n_743) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_524), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_526), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g651 ( .A(n_526), .Y(n_651) );
AND2x2_ASAP7_75t_L g713 ( .A(n_526), .B(n_634), .Y(n_713) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .Y(n_526) );
OR2x2_ASAP7_75t_L g567 ( .A(n_527), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g577 ( .A(n_527), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_527), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g685 ( .A(n_527), .Y(n_685) );
AND2x2_ASAP7_75t_L g702 ( .A(n_527), .B(n_549), .Y(n_702) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g593 ( .A(n_528), .B(n_538), .Y(n_593) );
AND2x2_ASAP7_75t_L g622 ( .A(n_528), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g633 ( .A(n_528), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_528), .B(n_588), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g548 ( .A(n_539), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g568 ( .A(n_539), .Y(n_568) );
AND2x2_ASAP7_75t_L g624 ( .A(n_539), .B(n_588), .Y(n_624) );
INVx1_ASAP7_75t_L g726 ( .A(n_547), .Y(n_726) );
INVx1_ASAP7_75t_L g730 ( .A(n_548), .Y(n_730) );
INVx2_ASAP7_75t_L g588 ( .A(n_549), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_559), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_559), .B(n_664), .Y(n_722) );
OR2x2_ASAP7_75t_L g563 ( .A(n_560), .B(n_561), .Y(n_563) );
INVx1_ASAP7_75t_SL g615 ( .A(n_560), .Y(n_615) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_566), .A2(n_619), .B1(n_621), .B2(n_625), .C(n_626), .Y(n_618) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g646 ( .A(n_567), .B(n_610), .Y(n_646) );
INVx2_ASAP7_75t_L g578 ( .A(n_568), .Y(n_578) );
INVx1_ASAP7_75t_L g604 ( .A(n_568), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_568), .B(n_588), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_568), .B(n_591), .Y(n_698) );
INVx1_ASAP7_75t_L g706 ( .A(n_568), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_570), .B(n_574), .Y(n_620) );
AND2x4_ASAP7_75t_L g595 ( .A(n_571), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g708 ( .A(n_574), .B(n_664), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_577), .B(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_L g716 ( .A(n_578), .Y(n_716) );
INVxp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g616 ( .A(n_582), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g688 ( .A(n_582), .B(n_664), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_582), .B(n_601), .Y(n_694) );
AOI322xp5_ASAP7_75t_L g648 ( .A1(n_583), .A2(n_617), .A3(n_624), .B1(n_649), .B2(n_652), .C1(n_653), .C2(n_655), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_583), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g714 ( .A(n_586), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g660 ( .A(n_587), .Y(n_660) );
INVx2_ASAP7_75t_L g591 ( .A(n_588), .Y(n_591) );
INVx1_ASAP7_75t_L g650 ( .A(n_588), .Y(n_650) );
CKINVDCx16_ASAP7_75t_R g597 ( .A(n_589), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g686 ( .A(n_591), .B(n_599), .Y(n_686) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_593), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g641 ( .A(n_593), .B(n_634), .Y(n_641) );
AND2x2_ASAP7_75t_L g645 ( .A(n_593), .B(n_605), .Y(n_645) );
OAI21xp33_ASAP7_75t_SL g655 ( .A1(n_594), .A2(n_656), .B(n_658), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_594), .A2(n_726), .B1(n_727), .B2(n_729), .Y(n_725) );
INVx3_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_595), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_595), .B(n_615), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_597), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g737 ( .A(n_604), .Y(n_737) );
INVx4_ASAP7_75t_L g610 ( .A(n_605), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_605), .B(n_632), .Y(n_680) );
INVx1_ASAP7_75t_SL g692 ( .A(n_606), .Y(n_692) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp67_ASAP7_75t_L g705 ( .A(n_610), .B(n_706), .Y(n_705) );
OAI211xp5_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_613), .B(n_618), .C(n_635), .Y(n_611) );
OAI221xp5_ASAP7_75t_SL g731 ( .A1(n_613), .A2(n_651), .B1(n_730), .B2(n_732), .C(n_734), .Y(n_731) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_615), .B(n_728), .Y(n_727) );
OAI31xp33_ASAP7_75t_L g707 ( .A1(n_616), .A2(n_693), .A3(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g647 ( .A(n_617), .Y(n_647) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g697 ( .A(n_622), .Y(n_697) );
AND2x2_ASAP7_75t_L g710 ( .A(n_624), .B(n_633), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_634), .B(n_737), .Y(n_736) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_641), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI221xp5_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_644), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_643), .A2(n_712), .B(n_714), .C(n_717), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_646), .B(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g673 ( .A(n_654), .Y(n_673) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g659 ( .A(n_657), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g701 ( .A(n_657), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_667), .C(n_676), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g738 ( .A1(n_665), .A2(n_675), .B1(n_739), .B2(n_740), .C(n_742), .Y(n_738) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B1(n_671), .B2(n_674), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI21xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B(n_679), .Y(n_676) );
INVx1_ASAP7_75t_SL g739 ( .A(n_678), .Y(n_739) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR4xp25_ASAP7_75t_L g681 ( .A(n_682), .B(n_711), .C(n_731), .D(n_738), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B(n_689), .C(n_707), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B(n_695), .C(n_699), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g718 ( .A(n_696), .Y(n_718) );
OR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
OR2x2_ASAP7_75t_L g729 ( .A(n_697), .B(n_730), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B(n_704), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_721), .B2(n_723), .C(n_725), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_728), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule