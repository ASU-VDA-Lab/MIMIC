module real_jpeg_27250_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_342, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_342;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_0),
.B(n_56),
.Y(n_96)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_29),
.B1(n_56),
.B2(n_58),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_4),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_4),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_122),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_122),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_56),
.B1(n_58),
.B2(n_122),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_6),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_6),
.A2(n_31),
.B(n_35),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_126),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_33),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_6),
.A2(n_62),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_6),
.B(n_62),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_6),
.B(n_78),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_6),
.A2(n_95),
.B1(n_250),
.B2(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_6),
.A2(n_34),
.B(n_266),
.Y(n_265)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_8),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_116),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_116),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_8),
.A2(n_56),
.B1(n_58),
.B2(n_116),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_9),
.A2(n_53),
.B1(n_56),
.B2(n_58),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_9),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_53),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_10),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_111),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_111),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_10),
.A2(n_56),
.B1(n_58),
.B2(n_111),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_12),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_113),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_12),
.A2(n_56),
.B1(n_58),
.B2(n_113),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_113),
.Y(n_270)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_15),
.A2(n_39),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_15),
.A2(n_39),
.B1(n_56),
.B2(n_58),
.Y(n_135)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_16),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_17),
.A2(n_62),
.B1(n_63),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_17),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_17),
.A2(n_34),
.B1(n_35),
.B2(n_106),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_17),
.A2(n_26),
.B1(n_27),
.B2(n_106),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_17),
.A2(n_56),
.B1(n_58),
.B2(n_106),
.Y(n_201)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_43),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_41),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_23),
.B(n_45),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_25),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_31),
.Y(n_32)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_27),
.A2(n_37),
.B(n_126),
.C(n_127),
.Y(n_125)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_33),
.B(n_38),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_33),
.B1(n_49),
.B2(n_52),
.Y(n_48)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_30),
.A2(n_33),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_30),
.A2(n_33),
.B1(n_112),
.B2(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_30),
.A2(n_33),
.B1(n_121),
.B2(n_193),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_33),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_34),
.A2(n_70),
.B(n_72),
.C(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_70),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_34),
.A2(n_63),
.A3(n_74),
.B1(n_267),
.B2(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_35),
.B(n_126),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_86),
.B(n_338),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_79),
.C(n_81),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_46),
.A2(n_47),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.C(n_67),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_48),
.B(n_323),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_50),
.A2(n_83),
.B1(n_85),
.B2(n_173),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_52),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_54),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_54),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_54),
.A2(n_67),
.B1(n_317),
.B2(n_324),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B(n_66),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_60),
.B1(n_104),
.B2(n_107),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_55),
.A2(n_60),
.B1(n_107),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_55),
.A2(n_60),
.B1(n_66),
.B2(n_146),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_55),
.A2(n_60),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_55),
.A2(n_60),
.B1(n_224),
.B2(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_55),
.B(n_126),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_55),
.A2(n_60),
.B1(n_191),
.B2(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_56),
.B(n_59),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_56),
.B(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_58),
.A2(n_62),
.A3(n_65),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_63),
.B1(n_71),
.B2(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_62),
.B(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_67),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_78),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_68),
.A2(n_78),
.B1(n_117),
.B2(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_68),
.A2(n_78),
.B1(n_187),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_68),
.A2(n_76),
.B1(n_78),
.B2(n_315),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_73),
.B(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_73),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_69),
.A2(n_73),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_69),
.A2(n_73),
.B1(n_131),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_69),
.A2(n_73),
.B1(n_199),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_74),
.Y(n_276)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_77),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_79),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_85),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_83),
.A2(n_85),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_331),
.B(n_337),
.Y(n_86)
);

OAI321xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_308),
.A3(n_327),
.B1(n_329),
.B2(n_330),
.C(n_341),
.Y(n_87)
);

AOI321xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_157),
.A3(n_179),
.B1(n_302),
.B2(n_307),
.C(n_342),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_90),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_138),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_91),
.B(n_138),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_118),
.C(n_133),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_92),
.B(n_133),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_108),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_109),
.C(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_94),
.B(n_103),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_99),
.B2(n_102),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_99),
.B1(n_102),
.B2(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_95),
.A2(n_99),
.B(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_95),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_95),
.A2(n_101),
.B1(n_244),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_95),
.A2(n_238),
.B1(n_239),
.B2(n_278),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_96),
.A2(n_100),
.B1(n_129),
.B2(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_96),
.A2(n_100),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_SL g239 ( 
.A(n_100),
.Y(n_239)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_101),
.B(n_126),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_105),
.A2(n_144),
.B1(n_147),
.B2(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.C(n_130),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_119),
.B(n_130),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_124),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_128),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_137),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_156),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_150),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_150),
.C(n_156),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_148),
.B2(n_149),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_144),
.A2(n_147),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_149),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_148),
.A2(n_171),
.B(n_174),
.Y(n_319)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_150),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.CI(n_155),
.CON(n_150),
.SN(n_150)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_158),
.B(n_159),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_177),
.B2(n_178),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_162),
.B(n_168),
.C(n_178),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_166),
.B(n_167),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_166),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_165),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_167),
.B(n_310),
.CI(n_319),
.CON(n_309),
.SN(n_309)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_209),
.C(n_214),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_203),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_181),
.B(n_203),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_194),
.C(n_195),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_182),
.B(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_192),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_189),
.C(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_300),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_194),
.Y(n_300)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_197),
.B(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_200),
.B(n_202),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_201),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.C(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_210),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_211),
.B(n_212),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_296),
.B(n_301),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_282),
.B(n_295),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_260),
.B(n_281),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_240),
.B(n_259),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_229),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_219),
.B(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_235),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_258),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_246),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_252),
.B(n_257),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_262),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_273),
.B1(n_279),
.B2(n_280),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_272),
.C(n_280),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_283),
.B(n_284),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_291),
.C(n_293),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_320),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_309),
.B(n_328),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_320),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_318),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_312),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_314),
.C(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_325),
.C(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);


endmodule