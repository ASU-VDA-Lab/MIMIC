module fake_netlist_1_8243_n_35 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_6), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_6), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_2), .B(n_7), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_10), .B(n_1), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_11), .B(n_3), .Y(n_20) );
NOR2x1p5_ASAP7_75t_L g21 ( .A(n_19), .B(n_12), .Y(n_21) );
CKINVDCx16_ASAP7_75t_R g22 ( .A(n_19), .Y(n_22) );
OR2x6_ASAP7_75t_L g23 ( .A(n_18), .B(n_15), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_19), .A2(n_15), .B1(n_14), .B2(n_13), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_22), .B(n_16), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_21), .B(n_16), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_23), .B(n_20), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_25), .B(n_24), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_25), .B1(n_27), .B2(n_23), .Y(n_30) );
AOI21xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_24), .B(n_23), .Y(n_31) );
OA21x2_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_17), .B(n_28), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_30), .Y(n_33) );
OAI22xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_9), .B1(n_29), .B2(n_17), .Y(n_34) );
AOI22xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_32), .B1(n_8), .B2(n_4), .Y(n_35) );
endmodule