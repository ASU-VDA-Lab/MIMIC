module real_aes_1624_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
AOI221xp5_ASAP7_75t_L g8 ( .A1(n_1), .A2(n_9), .B1(n_18), .B2(n_19), .C(n_21), .Y(n_8) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_1), .B(n_4), .Y(n_18) );
CKINVDCx16_ASAP7_75t_R g28 ( .A(n_2), .Y(n_28) );
INVx3_ASAP7_75t_L g31 ( .A(n_3), .Y(n_31) );
INVx1_ASAP7_75t_SL g20 ( .A(n_4), .Y(n_20) );
AND2x4_ASAP7_75t_L g16 ( .A(n_5), .B(n_17), .Y(n_16) );
INVx1_ASAP7_75t_L g33 ( .A(n_5), .Y(n_33) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVxp67_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_9), .B(n_20), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
OR2x2_ASAP7_75t_L g10 ( .A(n_11), .B(n_15), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_13), .B(n_14), .Y(n_12) );
INVxp67_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g24 ( .A(n_17), .Y(n_24) );
CKINVDCx14_ASAP7_75t_R g21 ( .A(n_22), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_23), .B(n_25), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_26), .B(n_32), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
NOR2xp33_ASAP7_75t_L g27 ( .A(n_28), .B(n_29), .Y(n_27) );
INVx2_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
CKINVDCx14_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
endmodule