module fake_jpeg_3270_n_573 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_573);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_573;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_65),
.Y(n_108)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g156 ( 
.A(n_56),
.Y(n_156)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_49),
.Y(n_61)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_66),
.Y(n_162)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_67),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_15),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_0),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_86),
.B(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_45),
.B(n_13),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_40),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_24),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_98),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_24),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_13),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_13),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_34),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_113),
.B(n_139),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_115),
.B(n_124),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_85),
.Y(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_61),
.A2(n_39),
.B1(n_33),
.B2(n_20),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_130),
.A2(n_169),
.B1(n_49),
.B2(n_74),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_157),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_58),
.A2(n_26),
.B1(n_24),
.B2(n_41),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_160),
.B1(n_170),
.B2(n_21),
.Y(n_177)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_148),
.Y(n_197)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_150),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_91),
.Y(n_157)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_59),
.A2(n_41),
.B1(n_26),
.B2(n_34),
.Y(n_160)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_71),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_60),
.A2(n_26),
.B1(n_41),
.B2(n_50),
.Y(n_170)
);

BUFx16f_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

CKINVDCx12_ASAP7_75t_R g172 ( 
.A(n_114),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_172),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_173),
.B(n_200),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_132),
.A2(n_93),
.B1(n_73),
.B2(n_75),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_174),
.B(n_179),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_113),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_175),
.B(n_176),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_30),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_177),
.A2(n_189),
.B1(n_145),
.B2(n_123),
.Y(n_254)
);

CKINVDCx12_ASAP7_75t_R g178 ( 
.A(n_134),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_178),
.Y(n_256)
);

OR2x2_ASAP7_75t_SL g179 ( 
.A(n_112),
.B(n_104),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_37),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_181),
.B(n_176),
.Y(n_267)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_122),
.B(n_62),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_184),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_21),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_193),
.Y(n_234)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_187),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_112),
.A2(n_80),
.B1(n_82),
.B2(n_68),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_92),
.B(n_84),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_191),
.A2(n_110),
.B(n_116),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_126),
.B(n_21),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_194),
.A2(n_199),
.B1(n_207),
.B2(n_210),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_46),
.B1(n_37),
.B2(n_30),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_198),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_120),
.A2(n_46),
.B1(n_36),
.B2(n_52),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_108),
.B(n_21),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_216),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_158),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_205),
.B(n_213),
.Y(n_266)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_140),
.A2(n_48),
.B1(n_36),
.B2(n_52),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_107),
.B(n_56),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_214),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_162),
.A2(n_42),
.B1(n_48),
.B2(n_33),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_158),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_56),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_146),
.Y(n_215)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_139),
.B(n_42),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_108),
.A2(n_49),
.B(n_77),
.C(n_76),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_222),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_49),
.B(n_12),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_220),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_118),
.A2(n_35),
.B1(n_95),
.B2(n_103),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_138),
.A2(n_33),
.B1(n_35),
.B2(n_51),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_223),
.A2(n_224),
.B1(n_131),
.B2(n_144),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_111),
.A2(n_33),
.B1(n_35),
.B2(n_2),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_119),
.Y(n_225)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_L g230 ( 
.A(n_121),
.B(n_0),
.C(n_1),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_3),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_119),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_143),
.B1(n_147),
.B2(n_123),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_169),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_3),
.Y(n_285)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_233),
.Y(n_273)
);

OR2x6_ASAP7_75t_L g238 ( 
.A(n_179),
.B(n_166),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_238),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_243),
.A2(n_184),
.B(n_194),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_261),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_211),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_254),
.A2(n_258),
.B1(n_225),
.B2(n_209),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_191),
.A2(n_166),
.B1(n_145),
.B2(n_164),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_171),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g323 ( 
.A1(n_264),
.A2(n_228),
.B1(n_196),
.B2(n_229),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_171),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_197),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_267),
.B(n_185),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_175),
.A2(n_161),
.B1(n_147),
.B2(n_143),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_181),
.B(n_161),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_174),
.A2(n_194),
.B1(n_222),
.B2(n_208),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_283),
.Y(n_313)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_180),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_183),
.B(n_156),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_203),
.B(n_156),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_180),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_208),
.B(n_133),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_4),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_214),
.A2(n_133),
.B1(n_131),
.B2(n_6),
.Y(n_286)
);

INVx3_ASAP7_75t_SL g326 ( 
.A(n_286),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_217),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_285),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_203),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_293),
.B(n_299),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_214),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_337),
.C(n_274),
.Y(n_338)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_194),
.B1(n_187),
.B2(n_232),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_297),
.A2(n_310),
.B1(n_283),
.B2(n_260),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_298),
.A2(n_260),
.B(n_262),
.Y(n_342)
);

OAI21xp33_ASAP7_75t_L g368 ( 
.A1(n_300),
.A2(n_317),
.B(n_336),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_234),
.B(n_182),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_301),
.B(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_197),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_267),
.B(n_204),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_309),
.Y(n_344)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_305),
.Y(n_359)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_239),
.Y(n_306)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

INVx11_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_308),
.A2(n_270),
.B1(n_248),
.B2(n_246),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_244),
.B(n_206),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_250),
.A2(n_192),
.B1(n_190),
.B2(n_188),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_235),
.B(n_185),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_312),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_249),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_240),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_314),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_266),
.B(n_190),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_316),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_252),
.B(n_188),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_237),
.B(n_192),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_324),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_240),
.Y(n_320)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_320),
.Y(n_380)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_321),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_238),
.B(n_209),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_245),
.B(n_209),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_327),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_273),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_195),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

CKINVDCx12_ASAP7_75t_R g330 ( 
.A(n_265),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_330),
.Y(n_370)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_255),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_333),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_237),
.B(n_202),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_257),
.Y(n_333)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_335),
.Y(n_354)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_270),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_259),
.B(n_227),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_237),
.B(n_226),
.C(n_219),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_302),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_296),
.A2(n_262),
.B1(n_250),
.B2(n_258),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_341),
.B1(n_360),
.B2(n_363),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_296),
.A2(n_262),
.B1(n_241),
.B2(n_243),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_342),
.A2(n_372),
.B(n_375),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_346),
.A2(n_350),
.B1(n_356),
.B2(n_292),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_294),
.B(n_278),
.C(n_238),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_376),
.C(n_377),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_297),
.A2(n_278),
.B1(n_268),
.B2(n_238),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g357 ( 
.A1(n_324),
.A2(n_287),
.B1(n_238),
.B2(n_269),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_357),
.A2(n_290),
.B1(n_307),
.B2(n_326),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_322),
.A2(n_269),
.B1(n_272),
.B2(n_246),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_322),
.A2(n_285),
.B(n_248),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_361),
.A2(n_365),
.B(n_381),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_298),
.A2(n_272),
.B1(n_284),
.B2(n_242),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_313),
.A2(n_242),
.B(n_284),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_313),
.A2(n_247),
.B1(n_215),
.B2(n_263),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_366),
.A2(n_335),
.B1(n_310),
.B2(n_306),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_259),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_378),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_300),
.A2(n_253),
.B(n_263),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_290),
.A2(n_253),
.B(n_282),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_299),
.B(n_5),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_7),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_311),
.B(n_315),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_316),
.A2(n_7),
.B(n_8),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_289),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_383),
.B(n_385),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_356),
.A2(n_346),
.B1(n_362),
.B2(n_345),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_384),
.A2(n_389),
.B1(n_343),
.B2(n_367),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_348),
.B(n_291),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_337),
.C(n_318),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_387),
.B(n_393),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_412),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_362),
.A2(n_326),
.B1(n_308),
.B2(n_317),
.Y(n_389)
);

INVx13_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

BUFx24_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_395),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_333),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_397),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_398),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_344),
.B(n_305),
.Y(n_399)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_319),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_401),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_342),
.A2(n_361),
.B(n_341),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_402),
.A2(n_404),
.B(n_416),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_321),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_403),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_345),
.A2(n_332),
.B(n_326),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_349),
.B(n_368),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_407),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_295),
.Y(n_408)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_339),
.A2(n_336),
.B1(n_323),
.B2(n_288),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_409),
.A2(n_410),
.B1(n_349),
.B2(n_375),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_366),
.A2(n_323),
.B1(n_288),
.B2(n_292),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_353),
.Y(n_411)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_411),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_330),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_418),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_365),
.A2(n_323),
.B(n_334),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_371),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_420),
.A2(n_425),
.B1(n_446),
.B2(n_353),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_402),
.A2(n_343),
.B1(n_378),
.B2(n_372),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_408),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_435),
.B(n_406),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_438),
.A2(n_448),
.B1(n_394),
.B2(n_395),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_396),
.B(n_354),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_354),
.Y(n_441)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_441),
.Y(n_460)
);

BUFx24_ASAP7_75t_SL g444 ( 
.A(n_385),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_386),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_409),
.A2(n_340),
.B1(n_358),
.B2(n_374),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_373),
.Y(n_447)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_384),
.A2(n_394),
.B1(n_382),
.B2(n_392),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_418),
.B(n_373),
.Y(n_451)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_451),
.Y(n_468)
);

BUFx4f_ASAP7_75t_SL g452 ( 
.A(n_449),
.Y(n_452)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_461),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_439),
.A2(n_416),
.B(n_413),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_454),
.A2(n_476),
.B(n_424),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_451),
.B(n_390),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_455),
.Y(n_490)
);

XOR2x2_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_405),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_478),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_448),
.A2(n_438),
.B1(n_421),
.B2(n_424),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_458),
.A2(n_450),
.B1(n_442),
.B2(n_445),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_459),
.B(n_474),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_462),
.A2(n_475),
.B1(n_467),
.B2(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_417),
.Y(n_463)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_463),
.Y(n_494)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_464),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_465),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_SL g466 ( 
.A(n_425),
.B(n_414),
.C(n_387),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_469),
.C(n_473),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_386),
.C(n_428),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_376),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_470),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_423),
.B(n_404),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_480),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_413),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_420),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_390),
.C(n_389),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_427),
.B(n_377),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_432),
.A2(n_410),
.B1(n_381),
.B2(n_340),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_391),
.B(n_353),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_441),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_479),
.A2(n_421),
.B1(n_443),
.B2(n_446),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_433),
.B(n_415),
.Y(n_480)
);

MAJx2_ASAP7_75t_L g509 ( 
.A(n_481),
.B(n_487),
.C(n_457),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_455),
.A2(n_454),
.B(n_476),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_483),
.A2(n_501),
.B(n_437),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_486),
.A2(n_437),
.B(n_352),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_424),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_491),
.A2(n_458),
.B1(n_461),
.B2(n_463),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_479),
.A2(n_443),
.B1(n_419),
.B2(n_442),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_492),
.A2(n_502),
.B1(n_473),
.B2(n_460),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_493),
.A2(n_352),
.B1(n_320),
.B2(n_314),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_445),
.C(n_434),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_498),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_456),
.B(n_449),
.C(n_450),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_472),
.B(n_471),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_453),
.A2(n_426),
.B1(n_436),
.B2(n_358),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_488),
.Y(n_505)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_505),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_506),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_507),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_480),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_509),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_323),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_510),
.B(n_518),
.C(n_519),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_492),
.A2(n_452),
.B1(n_464),
.B2(n_400),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_512),
.A2(n_520),
.B1(n_521),
.B2(n_522),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_374),
.C(n_398),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_513),
.B(n_517),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_452),
.Y(n_515)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_515),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_489),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_320),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_484),
.B(n_329),
.C(n_437),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_484),
.B(n_498),
.C(n_501),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_494),
.A2(n_352),
.B1(n_437),
.B2(n_314),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_7),
.Y(n_522)
);

O2A1O1Ixp5_ASAP7_75t_L g524 ( 
.A1(n_519),
.A2(n_494),
.B(n_488),
.C(n_500),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_524),
.A2(n_532),
.B1(n_525),
.B2(n_531),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_493),
.C(n_495),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_527),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_495),
.C(n_486),
.Y(n_527)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_508),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_534),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_531),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_490),
.C(n_483),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_523),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_536),
.A2(n_490),
.B1(n_485),
.B2(n_491),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_541),
.A2(n_534),
.B1(n_497),
.B2(n_11),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_507),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_542),
.B(n_544),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_537),
.A2(n_523),
.B1(n_512),
.B2(n_506),
.Y(n_543)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_543),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_533),
.A2(n_516),
.B(n_500),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_509),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_545),
.B(n_546),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_535),
.B(n_489),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_510),
.C(n_520),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_550),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_539),
.B(n_497),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_551),
.A2(n_8),
.B(n_9),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_545),
.B(n_538),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_552),
.B(n_554),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_556),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_8),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_557),
.B(n_8),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_562),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_553),
.B(n_540),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_558),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_565),
.B(n_566),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_560),
.A2(n_559),
.B(n_547),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_564),
.A2(n_555),
.B1(n_548),
.B2(n_552),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_541),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_567),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_556),
.B(n_557),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_9),
.C(n_536),
.Y(n_572)
);

BUFx24_ASAP7_75t_SL g573 ( 
.A(n_572),
.Y(n_573)
);


endmodule