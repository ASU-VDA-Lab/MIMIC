module fake_jpeg_4981_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_8),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_47),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_26),
.B(n_29),
.C(n_21),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_64),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_28),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_67),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_80),
.B1(n_88),
.B2(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_59),
.B1(n_52),
.B2(n_61),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_30),
.B1(n_23),
.B2(n_18),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_80)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_39),
.B1(n_24),
.B2(n_55),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_60),
.B1(n_17),
.B2(n_25),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_96),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_56),
.B1(n_45),
.B2(n_69),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_121),
.B1(n_70),
.B2(n_90),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_60),
.B(n_63),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_17),
.B(n_25),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_68),
.B(n_49),
.C(n_19),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_111),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_118),
.B1(n_88),
.B2(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_108),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_29),
.C(n_21),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_30),
.B1(n_18),
.B2(n_23),
.Y(n_145)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_18),
.B1(n_30),
.B2(n_23),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_63),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_46),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_89),
.A2(n_53),
.B1(n_68),
.B2(n_20),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_46),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_124),
.B(n_144),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_129),
.Y(n_163)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_136),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_146),
.B1(n_114),
.B2(n_100),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_142),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_145),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_90),
.B1(n_76),
.B2(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_151),
.B(n_155),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_102),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_111),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_112),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_32),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_141),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_46),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_122),
.B(n_137),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_134),
.B(n_107),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_117),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_100),
.B1(n_116),
.B2(n_107),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_127),
.B1(n_98),
.B2(n_79),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_119),
.C(n_104),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_118),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_84),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_84),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_147),
.B1(n_145),
.B2(n_144),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_177),
.A2(n_180),
.B(n_155),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

XNOR2x2_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_134),
.Y(n_180)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_191),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_153),
.B(n_149),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_98),
.B1(n_128),
.B2(n_104),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_194),
.B1(n_203),
.B2(n_127),
.Y(n_223)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_169),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_200),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_199),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_156),
.A2(n_32),
.B1(n_83),
.B2(n_27),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_222),
.B(n_202),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_200),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_153),
.B1(n_163),
.B2(n_151),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_217),
.B1(n_219),
.B2(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_154),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_216),
.C(n_218),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_150),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_176),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_163),
.B(n_152),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_170),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_164),
.B(n_159),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_196),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_169),
.B(n_150),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_223),
.A2(n_224),
.B1(n_177),
.B2(n_198),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_138),
.B1(n_32),
.B2(n_25),
.Y(n_224)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_181),
.C(n_187),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_28),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_180),
.A2(n_27),
.B(n_28),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_142),
.C(n_140),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_218),
.C(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_28),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_8),
.B(n_14),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_179),
.B1(n_203),
.B2(n_192),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_238),
.B1(n_246),
.B2(n_208),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_227),
.C(n_205),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_183),
.B1(n_184),
.B2(n_191),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_182),
.C(n_186),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_228),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_184),
.C(n_194),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_244),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_212),
.B(n_47),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_142),
.C(n_140),
.Y(n_244)
);

INVxp33_ASAP7_75t_SL g245 ( 
.A(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_250),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_27),
.B1(n_93),
.B2(n_83),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_28),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_28),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_222),
.A2(n_93),
.B1(n_31),
.B2(n_19),
.Y(n_250)
);

AOI21x1_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_226),
.B(n_206),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_254),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_260),
.B1(n_240),
.B2(n_244),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_257),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_215),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_232),
.A2(n_224),
.B1(n_19),
.B2(n_31),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_19),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_0),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_92),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_265),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_9),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_7),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_229),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_270),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_233),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_277),
.B(n_9),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_239),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_279),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_237),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_276),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_235),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_263),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_265),
.B1(n_10),
.B2(n_11),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_262),
.B1(n_252),
.B2(n_266),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_284),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_258),
.C(n_264),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_287),
.B(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_258),
.C(n_256),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_279),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_292),
.B(n_296),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_0),
.C(n_2),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_10),
.B(n_14),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_304),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_293),
.A2(n_282),
.B1(n_269),
.B2(n_2),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_300),
.C(n_5),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_290),
.B1(n_295),
.B2(n_294),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_3),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_11),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_15),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_10),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_12),
.B(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_285),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_310),
.B(n_313),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_311),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_314),
.B(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_6),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_15),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_299),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_308),
.B(n_12),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_308),
.B(n_315),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_13),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_13),
.B1(n_14),
.B2(n_3),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_13),
.C(n_3),
.Y(n_326)
);


endmodule