module fake_jpeg_5757_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_28),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_31),
.B1(n_19),
.B2(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_36),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_41),
.B(n_46),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_16),
.B(n_25),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_61),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_13),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_27),
.A2(n_19),
.B1(n_21),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_17),
.B1(n_18),
.B2(n_13),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_1),
.Y(n_78)
);

OR2x4_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_68),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_30),
.B(n_40),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_59),
.B(n_44),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_76),
.B1(n_45),
.B2(n_52),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_37),
.B1(n_21),
.B2(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_11),
.Y(n_91)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_87),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_41),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_64),
.C(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_58),
.B1(n_50),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_49),
.B1(n_46),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_47),
.B1(n_32),
.B2(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_85),
.C(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_92),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_64),
.B1(n_79),
.B2(n_78),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_83),
.B1(n_90),
.B2(n_87),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_81),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_106),
.C(n_107),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_67),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_100),
.B1(n_5),
.B2(n_7),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_102),
.B(n_97),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_114),
.B(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_103),
.C(n_67),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_115),
.A2(n_100),
.B1(n_110),
.B2(n_11),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_107),
.C(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_106),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_92),
.C(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_122),
.C(n_2),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_8),
.Y(n_125)
);


endmodule