module fake_jpeg_21082_n_159 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_79),
.Y(n_82)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_51),
.B1(n_71),
.B2(n_76),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_88),
.B1(n_49),
.B2(n_70),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_63),
.B1(n_65),
.B2(n_59),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_73),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_93),
.B(n_54),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_46),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_62),
.B1(n_64),
.B2(n_69),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_103),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_72),
.C(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_66),
.Y(n_105)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_88),
.B1(n_50),
.B2(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_56),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_55),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_117),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_58),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_57),
.B1(n_61),
.B2(n_60),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_116),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_25),
.C(n_44),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_125),
.A2(n_108),
.B1(n_120),
.B2(n_2),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_139),
.B1(n_0),
.B2(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_108),
.B(n_26),
.C(n_29),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_141),
.B1(n_0),
.B2(n_2),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

FAx1_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_124),
.CI(n_126),
.CON(n_143),
.SN(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_146),
.B(n_135),
.C(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_147),
.B1(n_134),
.B2(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_136),
.C(n_30),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_24),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_31),
.B(n_42),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_22),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_18),
.C(n_37),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_17),
.C(n_36),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_9),
.B(n_14),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_33),
.B(n_34),
.Y(n_159)
);


endmodule