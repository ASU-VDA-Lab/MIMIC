module fake_jpeg_28241_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_12),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_1),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_48),
.B1(n_53),
.B2(n_47),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_92),
.B1(n_83),
.B2(n_82),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_48),
.B1(n_70),
.B2(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_89),
.B1(n_67),
.B2(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_70),
.B1(n_62),
.B2(n_65),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_99),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_105),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_46),
.B1(n_55),
.B2(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_103),
.A2(n_91),
.B1(n_85),
.B2(n_50),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_59),
.B1(n_57),
.B2(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_88),
.B1(n_60),
.B2(n_63),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_115),
.B1(n_116),
.B2(n_104),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_69),
.B(n_3),
.C(n_4),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_5),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_59),
.B1(n_57),
.B2(n_51),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_52),
.B1(n_19),
.B2(n_43),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_121),
.B1(n_115),
.B2(n_10),
.Y(n_138)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_125),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_105),
.B1(n_52),
.B2(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_2),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_95),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_90),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_126),
.C(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_131),
.C(n_139),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_133),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_116),
.C(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_126),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_138),
.B1(n_140),
.B2(n_8),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_24),
.C(n_40),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_144),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_128),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_14),
.C(n_15),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_149),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_146),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_143),
.C(n_147),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_156),
.A2(n_143),
.B1(n_141),
.B2(n_137),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_150),
.C(n_136),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_16),
.CI(n_18),
.CON(n_159),
.SN(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_21),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_159),
.B(n_29),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_25),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_31),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_32),
.Y(n_164)
);


endmodule