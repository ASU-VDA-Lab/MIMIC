module real_aes_17963_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_51;
wire n_35;
wire n_42;
wire n_45;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
INVx2_ASAP7_75t_L g36 ( .A(n_0), .Y(n_36) );
INVx2_ASAP7_75t_L g39 ( .A(n_1), .Y(n_39) );
INVx1_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_3), .B(n_9), .Y(n_18) );
BUFx6f_ASAP7_75t_L g25 ( .A(n_4), .Y(n_25) );
AND2x2_ASAP7_75t_L g16 ( .A(n_5), .B(n_17), .Y(n_16) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_5), .Y(n_29) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_6), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_7), .B(n_34), .Y(n_33) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_11), .A2(n_19), .B1(n_26), .B2(n_37), .C(n_40), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g11 ( .A(n_12), .B(n_14), .Y(n_11) );
INVx1_ASAP7_75t_L g41 ( .A(n_12), .Y(n_41) );
INVx1_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
INVxp67_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_16), .B(n_18), .Y(n_15) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_17), .Y(n_31) );
INVx1_ASAP7_75t_L g47 ( .A(n_18), .Y(n_47) );
INVx1_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_22), .B(n_24), .Y(n_21) );
HB1xp67_ASAP7_75t_L g44 ( .A(n_22), .Y(n_44) );
INVx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
BUFx2_ASAP7_75t_L g51 ( .A(n_25), .Y(n_51) );
INVx1_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_28), .B(n_32), .Y(n_27) );
NOR2xp33_ASAP7_75t_L g28 ( .A(n_29), .B(n_30), .Y(n_28) );
INVx1_ASAP7_75t_L g45 ( .A(n_29), .Y(n_45) );
AOI221xp5_ASAP7_75t_SL g46 ( .A1(n_29), .A2(n_30), .B1(n_33), .B2(n_45), .C(n_47), .Y(n_46) );
INVx1_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
INVxp67_ASAP7_75t_SL g32 ( .A(n_33), .Y(n_32) );
INVx2_ASAP7_75t_SL g34 ( .A(n_35), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
BUFx3_ASAP7_75t_L g37 ( .A(n_38), .Y(n_37) );
INVx3_ASAP7_75t_L g38 ( .A(n_39), .Y(n_38) );
A2O1A1O1Ixp25_ASAP7_75t_L g40 ( .A1(n_41), .A2(n_42), .B(n_45), .C(n_46), .D(n_48), .Y(n_40) );
INVx1_ASAP7_75t_L g42 ( .A(n_43), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
INVx1_ASAP7_75t_L g48 ( .A(n_49), .Y(n_48) );
INVx1_ASAP7_75t_L g49 ( .A(n_50), .Y(n_49) );
INVx1_ASAP7_75t_L g50 ( .A(n_51), .Y(n_50) );
endmodule