module real_aes_4591_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_1083, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_1083;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_370;
wire n_1078;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_1053;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_973;
wire n_1081;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_769;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_1041;
wire n_488;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_1079;
wire n_843;
wire n_810;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1014;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1056;
wire n_358;
wire n_385;
wire n_397;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_354;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_756;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_307;
wire n_500;
wire n_601;
wire n_1076;
wire n_463;
wire n_661;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_877;
wire n_868;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_1061;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_0), .A2(n_115), .B1(n_650), .B2(n_777), .Y(n_776) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_1), .Y(n_309) );
AND2x4_ASAP7_75t_L g812 ( .A(n_1), .B(n_813), .Y(n_812) );
AND2x4_ASAP7_75t_L g821 ( .A(n_1), .B(n_287), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_2), .A2(n_245), .B1(n_531), .B2(n_772), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_3), .A2(n_45), .B1(n_818), .B2(n_822), .Y(n_817) );
XNOR2xp5_ASAP7_75t_L g1056 ( .A(n_4), .B(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_5), .A2(n_125), .B1(n_702), .B2(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g749 ( .A(n_6), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_7), .A2(n_58), .B1(n_387), .B2(n_437), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_8), .A2(n_113), .B1(n_836), .B2(n_837), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_9), .A2(n_17), .B1(n_449), .B2(n_468), .Y(n_467) );
AOI21xp33_ASAP7_75t_SL g1074 ( .A1(n_10), .A2(n_437), .B(n_1075), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_11), .A2(n_111), .B1(n_443), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_12), .A2(n_127), .B1(n_416), .B2(n_775), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_13), .A2(n_385), .B(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_14), .A2(n_294), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_15), .A2(n_172), .B1(n_504), .B2(n_505), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_16), .A2(n_150), .B1(n_443), .B2(n_675), .Y(n_674) );
XNOR2x2_ASAP7_75t_L g743 ( .A(n_18), .B(n_744), .Y(n_743) );
AO22x1_ASAP7_75t_L g692 ( .A1(n_19), .A2(n_21), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_20), .A2(n_146), .B1(n_416), .B2(n_418), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_22), .A2(n_80), .B1(n_501), .B2(n_502), .Y(n_599) );
INVx1_ASAP7_75t_L g700 ( .A(n_23), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_24), .A2(n_66), .B1(n_468), .B2(n_650), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_25), .A2(n_229), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_26), .A2(n_49), .B1(n_557), .B2(n_780), .C(n_781), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_27), .A2(n_74), .B1(n_371), .B2(n_374), .Y(n_370) );
INVx1_ASAP7_75t_SL g622 ( .A(n_28), .Y(n_622) );
INVx1_ASAP7_75t_L g519 ( .A(n_29), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g810 ( .A1(n_29), .A2(n_101), .B1(n_811), .B2(n_815), .Y(n_810) );
INVx1_ASAP7_75t_L g713 ( .A(n_30), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_31), .A2(n_194), .B1(n_446), .B2(n_449), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_32), .A2(n_40), .B1(n_451), .B2(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g782 ( .A(n_33), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_34), .B(n_224), .Y(n_307) );
INVx1_ASAP7_75t_L g345 ( .A(n_34), .Y(n_345) );
INVxp67_ASAP7_75t_L g396 ( .A(n_34), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_35), .A2(n_137), .B1(n_385), .B2(n_387), .Y(n_384) );
OA22x2_ASAP7_75t_L g726 ( .A1(n_36), .A2(n_727), .B1(n_739), .B2(n_740), .Y(n_726) );
INVx1_ASAP7_75t_L g740 ( .A(n_36), .Y(n_740) );
INVx1_ASAP7_75t_L g1039 ( .A(n_37), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_38), .A2(n_52), .B1(n_452), .B2(n_465), .Y(n_671) );
INVx1_ASAP7_75t_L g609 ( .A(n_39), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_41), .A2(n_212), .B1(n_818), .B2(n_822), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_42), .A2(n_151), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_43), .A2(n_272), .B1(n_826), .B2(n_847), .Y(n_891) );
INVx1_ASAP7_75t_L g595 ( .A(n_44), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_46), .B(n_331), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_47), .A2(n_109), .B1(n_678), .B2(n_680), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_48), .A2(n_124), .B1(n_374), .B2(n_676), .Y(n_1035) );
INVx1_ASAP7_75t_SL g613 ( .A(n_50), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_51), .A2(n_286), .B1(n_434), .B2(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g1076 ( .A(n_53), .Y(n_1076) );
INVx1_ASAP7_75t_L g711 ( .A(n_54), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_55), .A2(n_234), .B1(n_510), .B2(n_512), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_56), .A2(n_123), .B1(n_836), .B2(n_837), .Y(n_896) );
XNOR2x1_ASAP7_75t_L g1032 ( .A(n_56), .B(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_56), .A2(n_1054), .B1(n_1056), .B2(n_1077), .Y(n_1053) );
AOI21xp33_ASAP7_75t_L g593 ( .A1(n_57), .A2(n_517), .B(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_59), .A2(n_275), .B1(n_349), .B2(n_650), .Y(n_758) );
INVx1_ASAP7_75t_SL g619 ( .A(n_60), .Y(n_619) );
INVx2_ASAP7_75t_L g304 ( .A(n_61), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_62), .A2(n_184), .B1(n_509), .B2(n_518), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_63), .A2(n_130), .B1(n_540), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_64), .A2(n_143), .B1(n_324), .B2(n_454), .Y(n_747) );
INVx1_ASAP7_75t_SL g814 ( .A(n_65), .Y(n_814) );
AND2x4_ASAP7_75t_L g816 ( .A(n_65), .B(n_304), .Y(n_816) );
INVx1_ASAP7_75t_L g820 ( .A(n_65), .Y(n_820) );
INVx1_ASAP7_75t_SL g617 ( .A(n_67), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_68), .A2(n_77), .B1(n_632), .B2(n_635), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_69), .A2(n_97), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_70), .A2(n_216), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_71), .A2(n_187), .B1(n_535), .B2(n_537), .Y(n_1046) );
INVx1_ASAP7_75t_L g715 ( .A(n_72), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_73), .A2(n_185), .B1(n_534), .B2(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g578 ( .A(n_75), .Y(n_578) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_76), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_78), .A2(n_84), .B1(n_416), .B2(n_531), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_79), .A2(n_177), .B1(n_818), .B2(n_822), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_81), .A2(n_292), .B1(n_324), .B2(n_542), .Y(n_581) );
INVx1_ASAP7_75t_L g707 ( .A(n_82), .Y(n_707) );
INVx1_ASAP7_75t_L g844 ( .A(n_83), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_85), .A2(n_293), .B1(n_811), .B2(n_815), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_86), .A2(n_147), .B1(n_457), .B2(n_459), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_87), .A2(n_284), .B1(n_454), .B2(n_455), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_88), .A2(n_119), .B1(n_501), .B2(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g334 ( .A(n_89), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_89), .B(n_223), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_90), .A2(n_257), .B1(n_495), .B2(n_501), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_91), .A2(n_195), .B1(n_556), .B2(n_558), .Y(n_555) );
OAI22x1_ASAP7_75t_L g461 ( .A1(n_92), .A2(n_462), .B1(n_469), .B2(n_486), .Y(n_461) );
NAND5xp2_ASAP7_75t_SL g462 ( .A(n_92), .B(n_463), .C(n_464), .D(n_466), .E(n_467), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_92), .A2(n_102), .B1(n_811), .B2(n_815), .Y(n_827) );
INVx1_ASAP7_75t_L g754 ( .A(n_93), .Y(n_754) );
AO22x1_ASAP7_75t_L g433 ( .A1(n_94), .A2(n_117), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_95), .A2(n_259), .B1(n_764), .B2(n_1073), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_96), .A2(n_193), .B1(n_434), .B2(n_574), .Y(n_1036) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_98), .A2(n_430), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_99), .B(n_557), .Y(n_572) );
INVx1_ASAP7_75t_SL g641 ( .A(n_100), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_103), .A2(n_256), .B1(n_452), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_104), .A2(n_219), .B1(n_454), .B2(n_455), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_105), .A2(n_288), .B1(n_498), .B2(n_499), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_106), .A2(n_242), .B1(n_349), .B2(n_650), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_107), .B(n_432), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_108), .A2(n_141), .B1(n_374), .B2(n_561), .Y(n_575) );
AOI221xp5_ASAP7_75t_SL g733 ( .A1(n_110), .A2(n_262), .B1(n_512), .B2(n_676), .C(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_112), .A2(n_255), .B1(n_452), .B2(n_540), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_114), .A2(n_204), .B1(n_452), .B2(n_465), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_116), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_118), .A2(n_197), .B1(n_509), .B2(n_510), .C(n_737), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_120), .A2(n_432), .B(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_121), .A2(n_228), .B1(n_818), .B2(n_826), .Y(n_825) );
INVxp33_ASAP7_75t_SL g850 ( .A(n_122), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_126), .A2(n_165), .B1(n_387), .B2(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_128), .B(n_398), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_129), .B(n_1041), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_131), .A2(n_203), .B1(n_574), .B2(n_1069), .Y(n_1068) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_132), .A2(n_198), .B1(n_398), .B2(n_401), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_133), .A2(n_181), .B1(n_833), .B2(n_834), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_134), .A2(n_158), .B1(n_349), .B2(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_135), .A2(n_173), .B1(n_496), .B2(n_502), .Y(n_732) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_136), .B(n_324), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_138), .A2(n_209), .B1(n_504), .B2(n_505), .Y(n_600) );
INVx1_ASAP7_75t_L g788 ( .A(n_139), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_140), .A2(n_265), .B1(n_454), .B2(n_455), .Y(n_463) );
INVx1_ASAP7_75t_L g685 ( .A(n_142), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_144), .A2(n_246), .B1(n_457), .B2(n_459), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_145), .A2(n_160), .B1(n_535), .B2(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_148), .A2(n_217), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_149), .A2(n_190), .B1(n_537), .B2(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_152), .A2(n_235), .B1(n_410), .B2(n_446), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_153), .A2(n_183), .B1(n_387), .B2(n_561), .Y(n_762) );
INVx1_ASAP7_75t_L g474 ( .A(n_154), .Y(n_474) );
INVx1_ASAP7_75t_L g706 ( .A(n_155), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g1037 ( .A1(n_156), .A2(n_561), .B(n_1038), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_157), .A2(n_168), .B1(n_324), .B2(n_362), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1045 ( .A1(n_159), .A2(n_231), .B1(n_349), .B2(n_650), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_161), .A2(n_227), .B1(n_498), .B2(n_499), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_162), .A2(n_163), .B1(n_455), .B2(n_459), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_164), .A2(n_202), .B1(n_560), .B2(n_562), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_166), .A2(n_281), .B1(n_349), .B2(n_410), .Y(n_585) );
INVx1_ASAP7_75t_L g611 ( .A(n_167), .Y(n_611) );
INVx1_ASAP7_75t_L g848 ( .A(n_169), .Y(n_848) );
AO22x1_ASAP7_75t_L g737 ( .A1(n_170), .A2(n_253), .B1(n_518), .B2(n_738), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_171), .A2(n_258), .B1(n_495), .B2(n_496), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_174), .A2(n_280), .B1(n_531), .B2(n_535), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_175), .A2(n_191), .B1(n_434), .B2(n_720), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_176), .A2(n_261), .B1(n_495), .B2(n_496), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_178), .A2(n_282), .B1(n_362), .B2(n_535), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_179), .A2(n_218), .B1(n_530), .B2(n_532), .Y(n_529) );
XNOR2x1_ASAP7_75t_L g569 ( .A(n_180), .B(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_182), .Y(n_661) );
XOR2x2_ASAP7_75t_L g689 ( .A(n_186), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_188), .B(n_401), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g1060 ( .A1(n_189), .A2(n_237), .B1(n_459), .B2(n_1061), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_192), .A2(n_274), .B1(n_457), .B2(n_459), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_196), .A2(n_260), .B1(n_437), .B2(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g799 ( .A(n_199), .Y(n_799) );
INVx1_ASAP7_75t_L g333 ( .A(n_200), .Y(n_333) );
OA22x2_ASAP7_75t_L g359 ( .A1(n_200), .A2(n_224), .B1(n_331), .B2(n_357), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_201), .A2(n_221), .B1(n_410), .B2(n_412), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_205), .A2(n_239), .B1(n_574), .B2(n_764), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_206), .A2(n_248), .B1(n_717), .B2(n_797), .C(n_798), .Y(n_796) );
INVx1_ASAP7_75t_L g514 ( .A(n_207), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_208), .A2(n_545), .B(n_548), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_210), .A2(n_268), .B1(n_459), .B2(n_540), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_211), .A2(n_283), .B1(n_833), .B2(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g554 ( .A(n_213), .Y(n_554) );
AOI221x1_ASAP7_75t_L g348 ( .A1(n_214), .A2(n_266), .B1(n_349), .B2(n_362), .C(n_364), .Y(n_348) );
INVx1_ASAP7_75t_L g551 ( .A(n_215), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_220), .A2(n_264), .B1(n_468), .B2(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_222), .Y(n_426) );
INVx1_ASAP7_75t_L g347 ( .A(n_223), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_223), .B(n_329), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g335 ( .A1(n_224), .A2(n_240), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g364 ( .A(n_225), .B(n_365), .Y(n_364) );
AO22x2_ASAP7_75t_L g524 ( .A1(n_226), .A2(n_525), .B1(n_564), .B2(n_565), .Y(n_524) );
INVx1_ASAP7_75t_L g565 ( .A(n_226), .Y(n_565) );
INVx1_ASAP7_75t_L g890 ( .A(n_230), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_232), .A2(n_247), .B1(n_441), .B2(n_443), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_233), .A2(n_252), .B1(n_811), .B2(n_815), .Y(n_861) );
INVx1_ASAP7_75t_SL g648 ( .A(n_236), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_238), .A2(n_254), .B1(n_479), .B2(n_802), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_240), .B(n_277), .Y(n_308) );
INVx1_ASAP7_75t_L g356 ( .A(n_240), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_241), .A2(n_273), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g752 ( .A1(n_243), .A2(n_676), .B(n_753), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_244), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_249), .B(n_717), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_250), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g587 ( .A(n_251), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_263), .A2(n_267), .B1(n_539), .B2(n_541), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g321 ( .A(n_269), .B(n_322), .C(n_369), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_269), .A2(n_369), .B1(n_383), .B2(n_1083), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_269), .A2(n_322), .B(n_408), .Y(n_423) );
INVx1_ASAP7_75t_SL g640 ( .A(n_270), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_271), .A2(n_291), .B1(n_437), .B2(n_443), .Y(n_803) );
INVx1_ASAP7_75t_L g703 ( .A(n_276), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_277), .B(n_330), .Y(n_340) );
AOI21xp33_ASAP7_75t_L g511 ( .A1(n_278), .A2(n_512), .B(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_279), .A2(n_290), .B1(n_540), .B2(n_542), .Y(n_746) );
INVxp33_ASAP7_75t_L g842 ( .A(n_285), .Y(n_842) );
INVx1_ASAP7_75t_L g813 ( .A(n_287), .Y(n_813) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_287), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_289), .B(n_481), .Y(n_480) );
XNOR2x1_ASAP7_75t_L g768 ( .A(n_295), .B(n_769), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_296), .A2(n_430), .B(n_433), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_310), .B(n_805), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .C(n_309), .Y(n_301) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_302), .B(n_1051), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_302), .B(n_1052), .Y(n_1055) );
AOI21xp5_ASAP7_75t_L g1081 ( .A1(n_302), .A2(n_309), .B(n_814), .Y(n_1081) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AO21x1_ASAP7_75t_L g1078 ( .A1(n_303), .A2(n_1079), .B(n_1081), .Y(n_1078) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND3x4_ASAP7_75t_L g811 ( .A(n_304), .B(n_812), .C(n_814), .Y(n_811) );
AND2x2_ASAP7_75t_L g819 ( .A(n_304), .B(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g1051 ( .A(n_305), .B(n_1052), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_306), .A2(n_405), .B(n_406), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g1052 ( .A(n_309), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_723), .B2(n_804), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
XNOR2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_522), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_460), .B1(n_520), .B2(n_521), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g520 ( .A(n_315), .Y(n_520) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_424), .B2(n_425), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_382), .B(n_421), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_348), .Y(n_322) );
INVx5_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g637 ( .A(n_325), .Y(n_637) );
INVx3_ASAP7_75t_L g772 ( .A(n_325), .Y(n_772) );
INVx1_ASAP7_75t_L g1061 ( .A(n_325), .Y(n_1061) );
INVx6_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx12f_ASAP7_75t_L g455 ( .A(n_326), .Y(n_455) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_337), .Y(n_326) );
AND2x4_ASAP7_75t_L g375 ( .A(n_327), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g414 ( .A(n_327), .B(n_367), .Y(n_414) );
AND2x4_ASAP7_75t_L g496 ( .A(n_327), .B(n_337), .Y(n_496) );
AND2x4_ASAP7_75t_L g502 ( .A(n_327), .B(n_367), .Y(n_502) );
AND2x4_ASAP7_75t_L g518 ( .A(n_327), .B(n_376), .Y(n_518) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_335), .Y(n_327) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_328), .B(n_341), .C(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_330), .B(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g336 ( .A(n_331), .Y(n_336) );
NAND2xp33_ASAP7_75t_L g346 ( .A(n_331), .B(n_347), .Y(n_346) );
NAND2xp33_ASAP7_75t_L g354 ( .A(n_331), .B(n_334), .Y(n_354) );
INVx2_ASAP7_75t_L g357 ( .A(n_331), .Y(n_357) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_331), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_336), .A2(n_356), .B(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g363 ( .A(n_337), .B(n_351), .Y(n_363) );
AND2x4_ASAP7_75t_L g499 ( .A(n_337), .B(n_366), .Y(n_499) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g420 ( .A(n_338), .Y(n_420) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_342), .Y(n_338) );
AND2x4_ASAP7_75t_L g360 ( .A(n_339), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g367 ( .A(n_339), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g377 ( .A(n_339), .Y(n_377) );
AND2x2_ASAP7_75t_L g390 ( .A(n_339), .B(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g361 ( .A(n_343), .Y(n_361) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_349), .Y(n_647) );
BUFx12f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g448 ( .A(n_350), .Y(n_448) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_350), .Y(n_468) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_360), .Y(n_350) );
AND2x2_ASAP7_75t_L g411 ( .A(n_351), .B(n_376), .Y(n_411) );
AND2x4_ASAP7_75t_L g417 ( .A(n_351), .B(n_367), .Y(n_417) );
AND2x4_ASAP7_75t_L g495 ( .A(n_351), .B(n_420), .Y(n_495) );
AND2x4_ASAP7_75t_L g501 ( .A(n_351), .B(n_367), .Y(n_501) );
AND2x4_ASAP7_75t_L g504 ( .A(n_351), .B(n_360), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_351), .B(n_376), .Y(n_505) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_358), .Y(n_351) );
AND2x2_ASAP7_75t_L g381 ( .A(n_352), .B(n_359), .Y(n_381) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g366 ( .A(n_353), .B(n_359), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g394 ( .A(n_359), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g373 ( .A(n_360), .B(n_366), .Y(n_373) );
AND2x4_ASAP7_75t_L g386 ( .A(n_360), .B(n_381), .Y(n_386) );
AND2x4_ASAP7_75t_L g509 ( .A(n_360), .B(n_366), .Y(n_509) );
AND2x4_ASAP7_75t_L g512 ( .A(n_360), .B(n_381), .Y(n_512) );
AND2x4_ASAP7_75t_L g376 ( .A(n_361), .B(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g693 ( .A(n_362), .Y(n_693) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_363), .Y(n_454) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_363), .Y(n_531) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_363), .Y(n_634) );
BUFx4f_ASAP7_75t_L g583 ( .A(n_365), .Y(n_583) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_365), .Y(n_702) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g400 ( .A(n_366), .B(n_376), .Y(n_400) );
AND2x4_ASAP7_75t_L g419 ( .A(n_366), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g458 ( .A(n_366), .B(n_367), .Y(n_458) );
AND2x4_ASAP7_75t_L g498 ( .A(n_366), .B(n_367), .Y(n_498) );
AND2x2_ASAP7_75t_L g738 ( .A(n_366), .B(n_376), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_378), .Y(n_369) );
BUFx3_ASAP7_75t_L g680 ( .A(n_371), .Y(n_680) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_372), .Y(n_439) );
INVx1_ASAP7_75t_L g802 ( .A(n_372), .Y(n_802) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g478 ( .A(n_373), .Y(n_478) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_373), .Y(n_574) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_375), .Y(n_443) );
INVx3_ASAP7_75t_L g765 ( .A(n_375), .Y(n_765) );
AND2x4_ASAP7_75t_L g380 ( .A(n_376), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g517 ( .A(n_376), .B(n_381), .Y(n_517) );
BUFx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g442 ( .A(n_380), .Y(n_442) );
INVx2_ASAP7_75t_L g485 ( .A(n_380), .Y(n_485) );
BUFx8_ASAP7_75t_SL g557 ( .A(n_380), .Y(n_557) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_380), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_408), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_397), .Y(n_383) );
INVx2_ASAP7_75t_L g679 ( .A(n_385), .Y(n_679) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_386), .Y(n_437) );
BUFx3_ASAP7_75t_L g561 ( .A(n_386), .Y(n_561) );
INVx4_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g479 ( .A(n_388), .Y(n_479) );
INVx2_ASAP7_75t_L g550 ( .A(n_388), .Y(n_550) );
INVx2_ASAP7_75t_L g1069 ( .A(n_388), .Y(n_1069) );
INVx5_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g434 ( .A(n_389), .Y(n_434) );
BUFx2_ASAP7_75t_L g684 ( .A(n_389), .Y(n_684) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_394), .Y(n_389) );
AND2x2_ASAP7_75t_L g510 ( .A(n_390), .B(n_394), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g405 ( .A(n_392), .Y(n_405) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_399), .Y(n_482) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g432 ( .A(n_400), .Y(n_432) );
INVx3_ASAP7_75t_L g718 ( .A(n_400), .Y(n_718) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g1075 ( .A(n_402), .B(n_1076), .Y(n_1075) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_403), .Y(n_579) );
INVx2_ASAP7_75t_SL g625 ( .A(n_403), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_403), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g756 ( .A(n_403), .Y(n_756) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g476 ( .A(n_404), .Y(n_476) );
NAND2x1_ASAP7_75t_SL g408 ( .A(n_409), .B(n_415), .Y(n_408) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx5_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_411), .Y(n_650) );
INVx1_ASAP7_75t_L g670 ( .A(n_411), .Y(n_670) );
INVx4_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx4_ASAP7_75t_L g452 ( .A(n_413), .Y(n_452) );
INVx2_ASAP7_75t_L g537 ( .A(n_413), .Y(n_537) );
INVx1_ASAP7_75t_L g698 ( .A(n_413), .Y(n_698) );
INVx4_ASAP7_75t_L g760 ( .A(n_413), .Y(n_760) );
INVx2_ASAP7_75t_SL g775 ( .A(n_413), .Y(n_775) );
INVx1_ASAP7_75t_L g1065 ( .A(n_413), .Y(n_1065) );
INVx8_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx12f_ASAP7_75t_L g451 ( .A(n_416), .Y(n_451) );
INVx1_ASAP7_75t_L g630 ( .A(n_416), .Y(n_630) );
BUFx12f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_417), .Y(n_535) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
BUFx12f_ASAP7_75t_L g542 ( .A(n_419), .Y(n_542) );
BUFx3_ASAP7_75t_L g643 ( .A(n_419), .Y(n_643) );
BUFx6f_ASAP7_75t_L g1044 ( .A(n_419), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
XNOR2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_428), .B(n_444), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_436), .C(n_440), .Y(n_428) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx4_ASAP7_75t_L g612 ( .A(n_437), .Y(n_612) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g615 ( .A(n_439), .Y(n_615) );
INVx2_ASAP7_75t_L g709 ( .A(n_439), .Y(n_709) );
INVx2_ASAP7_75t_L g785 ( .A(n_439), .Y(n_785) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g797 ( .A(n_442), .Y(n_797) );
BUFx3_ASAP7_75t_L g558 ( .A(n_443), .Y(n_558) );
INVx4_ASAP7_75t_L g620 ( .A(n_443), .Y(n_620) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_450), .C(n_453), .D(n_456), .Y(n_444) );
BUFx4f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g777 ( .A(n_448), .Y(n_777) );
BUFx3_ASAP7_75t_L g528 ( .A(n_449), .Y(n_528) );
BUFx3_ASAP7_75t_L g532 ( .A(n_455), .Y(n_532) );
BUFx8_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_458), .Y(n_540) );
INVx2_ASAP7_75t_L g521 ( .A(n_460), .Y(n_521) );
XNOR2x1_ASAP7_75t_L g460 ( .A(n_461), .B(n_490), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g487 ( .A(n_463), .B(n_464), .C(n_467), .D(n_480), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_466), .B(n_483), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_480), .C(n_483), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g488 ( .A(n_471), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_477), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_475), .B(n_595), .Y(n_594) );
INVx4_ASAP7_75t_L g720 ( .A(n_475), .Y(n_720) );
INVx4_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
INVx2_ASAP7_75t_L g563 ( .A(n_478), .Y(n_563) );
INVx1_ASAP7_75t_L g623 ( .A(n_481), .Y(n_623) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g547 ( .A(n_482), .Y(n_547) );
INVx2_ASAP7_75t_L g751 ( .A(n_482), .Y(n_751) );
INVx2_ASAP7_75t_L g618 ( .A(n_484), .Y(n_618) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g1073 ( .A(n_485), .Y(n_1073) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_491), .Y(n_653) );
INVx2_ASAP7_75t_L g656 ( .A(n_491), .Y(n_656) );
XOR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_519), .Y(n_491) );
NOR2xp67_ASAP7_75t_L g492 ( .A(n_493), .B(n_506), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .C(n_500), .D(n_503), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .C(n_511), .D(n_516), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx4_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g1038 ( .A(n_515), .B(n_1039), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_604), .B1(n_721), .B2(n_722), .Y(n_522) );
INVx1_ASAP7_75t_L g722 ( .A(n_523), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_566), .B1(n_567), .B2(n_603), .Y(n_523) );
INVx4_ASAP7_75t_L g603 ( .A(n_524), .Y(n_603) );
INVx1_ASAP7_75t_L g564 ( .A(n_525), .Y(n_564) );
NOR2x1_ASAP7_75t_L g525 ( .A(n_526), .B(n_543), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .C(n_533), .D(n_538), .Y(n_526) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g639 ( .A(n_539), .Y(n_639) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .C(n_559), .Y(n_543) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_551), .B1(n_552), .B2(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_565), .A2(n_841), .B1(n_843), .B2(n_890), .C(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OA22x2_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_586), .B2(n_602), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_580), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .C(n_575), .D(n_576), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .C(n_584), .D(n_585), .Y(n_580) );
INVx2_ASAP7_75t_L g602 ( .A(n_586), .Y(n_602) );
AO21x2_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_601), .Y(n_586) );
NOR3xp33_ASAP7_75t_SL g601 ( .A(n_587), .B(n_589), .C(n_596), .Y(n_601) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_596), .Y(n_588) );
NAND4xp75_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .C(n_592), .D(n_593), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .C(n_599), .D(n_600), .Y(n_596) );
INVx1_ASAP7_75t_L g721 ( .A(n_604), .Y(n_721) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_658), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_653), .B1(n_654), .B2(n_657), .Y(n_605) );
INVx4_ASAP7_75t_L g657 ( .A(n_606), .Y(n_657) );
AO22x2_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_626), .B2(n_651), .Y(n_606) );
NOR4xp25_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .C(n_616), .D(n_621), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_609), .Y(n_608) );
NOR3xp33_ASAP7_75t_SL g652 ( .A(n_610), .B(n_616), .C(n_621), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_612), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_620), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_710) );
OAI21xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B(n_624), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_626), .B(n_652), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_638), .C(n_644), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_637), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_642), .A2(n_700), .B1(n_701), .B2(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI22x1_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_646), .B1(n_648), .B2(n_649), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVxp33_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_688), .B2(n_689), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AO21x2_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B(n_687), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_661), .B(n_664), .C(n_673), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_672), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND4xp25_ASAP7_75t_SL g664 ( .A(n_665), .B(n_666), .C(n_667), .D(n_671), .Y(n_664) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .C(n_681), .Y(n_673) );
INVx1_ASAP7_75t_L g712 ( .A(n_675), .Y(n_712) );
BUFx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_685), .B(n_686), .Y(n_682) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_704), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_695), .C(n_699), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_710), .C(n_714), .Y(n_704) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g780 ( .A(n_718), .Y(n_780) );
INVx2_ASAP7_75t_L g1041 ( .A(n_718), .Y(n_1041) );
INVx2_ASAP7_75t_L g800 ( .A(n_720), .Y(n_800) );
INVx1_ASAP7_75t_L g804 ( .A(n_723), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_741), .Y(n_723) );
BUFx4_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g739 ( .A(n_727), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_733), .C(n_736), .Y(n_727) );
AND4x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .C(n_731), .D(n_732), .Y(n_728) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_766), .Y(n_742) );
NAND4xp75_ASAP7_75t_L g744 ( .A(n_745), .B(n_748), .C(n_757), .D(n_761), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
OA21x2_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_755), .B(n_782), .Y(n_781) );
INVx3_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx3_ASAP7_75t_L g786 ( .A(n_765), .Y(n_786) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
XNOR2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_787), .Y(n_767) );
NOR2x1_ASAP7_75t_L g769 ( .A(n_770), .B(n_778), .Y(n_769) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .C(n_774), .D(n_776), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_783), .C(n_784), .Y(n_778) );
XNOR2x1_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_795), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .C(n_793), .D(n_794), .Y(n_790) );
NAND3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_801), .C(n_803), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_1028), .B1(n_1030), .B2(n_1048), .C(n_1053), .Y(n_805) );
AOI211x1_ASAP7_75t_SL g806 ( .A1(n_807), .A2(n_885), .B(n_898), .C(n_1006), .Y(n_806) );
OAI211xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_828), .B(n_854), .C(n_874), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_823), .Y(n_808) );
INVx1_ASAP7_75t_L g859 ( .A(n_809), .Y(n_859) );
OR2x2_ASAP7_75t_L g877 ( .A(n_809), .B(n_860), .Y(n_877) );
AND2x2_ASAP7_75t_L g915 ( .A(n_809), .B(n_860), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_809), .B(n_824), .Y(n_934) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_817), .Y(n_809) );
AND2x4_ASAP7_75t_L g815 ( .A(n_812), .B(n_816), .Y(n_815) );
AND2x4_ASAP7_75t_L g833 ( .A(n_812), .B(n_819), .Y(n_833) );
AND2x4_ASAP7_75t_L g834 ( .A(n_812), .B(n_816), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_812), .B(n_816), .Y(n_843) );
AND2x2_ASAP7_75t_L g822 ( .A(n_816), .B(n_821), .Y(n_822) );
AND2x4_ASAP7_75t_L g826 ( .A(n_816), .B(n_821), .Y(n_826) );
AND2x2_ASAP7_75t_L g837 ( .A(n_816), .B(n_821), .Y(n_837) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_821), .Y(n_818) );
AND2x2_ASAP7_75t_L g836 ( .A(n_819), .B(n_821), .Y(n_836) );
AND2x4_ASAP7_75t_L g847 ( .A(n_819), .B(n_821), .Y(n_847) );
NOR2x1_ASAP7_75t_R g871 ( .A(n_823), .B(n_872), .Y(n_871) );
AND2x2_ASAP7_75t_L g911 ( .A(n_823), .B(n_858), .Y(n_911) );
AND2x2_ASAP7_75t_L g929 ( .A(n_823), .B(n_859), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_823), .B(n_963), .Y(n_962) );
AND2x2_ASAP7_75t_L g976 ( .A(n_823), .B(n_915), .Y(n_976) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_823), .B(n_967), .Y(n_1003) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_SL g857 ( .A(n_824), .Y(n_857) );
AND2x2_ASAP7_75t_L g868 ( .A(n_824), .B(n_869), .Y(n_868) );
OR2x2_ASAP7_75t_L g904 ( .A(n_824), .B(n_870), .Y(n_904) );
AND2x2_ASAP7_75t_L g966 ( .A(n_824), .B(n_967), .Y(n_966) );
OR2x2_ASAP7_75t_L g996 ( .A(n_824), .B(n_877), .Y(n_996) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_824), .B(n_859), .Y(n_1008) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
INVx2_ASAP7_75t_L g849 ( .A(n_826), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_838), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_829), .B(n_929), .Y(n_928) );
NAND2xp67_ASAP7_75t_L g1026 ( .A(n_829), .B(n_855), .Y(n_1026) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NOR2x1_ASAP7_75t_L g869 ( .A(n_830), .B(n_870), .Y(n_869) );
NAND2xp5_ASAP7_75t_SL g872 ( .A(n_830), .B(n_873), .Y(n_872) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_830), .Y(n_883) );
INVx2_ASAP7_75t_L g903 ( .A(n_830), .Y(n_903) );
INVx1_ASAP7_75t_L g917 ( .A(n_830), .Y(n_917) );
AND2x2_ASAP7_75t_L g959 ( .A(n_830), .B(n_839), .Y(n_959) );
AND2x2_ASAP7_75t_L g965 ( .A(n_830), .B(n_966), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_830), .B(n_908), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_830), .B(n_929), .Y(n_986) );
AND2x2_ASAP7_75t_L g994 ( .A(n_830), .B(n_906), .Y(n_994) );
INVx4_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_831), .B(n_866), .Y(n_935) );
OR2x2_ASAP7_75t_L g939 ( .A(n_831), .B(n_856), .Y(n_939) );
AND2x2_ASAP7_75t_L g954 ( .A(n_831), .B(n_839), .Y(n_954) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_835), .Y(n_831) );
INVx3_ASAP7_75t_L g841 ( .A(n_833), .Y(n_841) );
INVx1_ASAP7_75t_L g941 ( .A(n_838), .Y(n_941) );
AND2x2_ASAP7_75t_L g838 ( .A(n_839), .B(n_851), .Y(n_838) );
INVx2_ASAP7_75t_L g866 ( .A(n_839), .Y(n_866) );
INVx1_ASAP7_75t_L g906 ( .A(n_839), .Y(n_906) );
OR2x2_ASAP7_75t_L g948 ( .A(n_839), .B(n_851), .Y(n_948) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_839), .B(n_955), .Y(n_1000) );
OR2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_845), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_843), .B2(n_844), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_848), .B1(n_849), .B2(n_850), .Y(n_845) );
INVx3_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_847), .Y(n_1029) );
OR2x2_ASAP7_75t_L g879 ( .A(n_851), .B(n_866), .Y(n_879) );
AND2x2_ASAP7_75t_L g884 ( .A(n_851), .B(n_866), .Y(n_884) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_851), .Y(n_918) );
OR2x2_ASAP7_75t_L g922 ( .A(n_851), .B(n_894), .Y(n_922) );
AND2x2_ASAP7_75t_L g931 ( .A(n_851), .B(n_893), .Y(n_931) );
OR2x2_ASAP7_75t_L g950 ( .A(n_851), .B(n_895), .Y(n_950) );
AND2x2_ASAP7_75t_L g955 ( .A(n_851), .B(n_894), .Y(n_955) );
INVx2_ASAP7_75t_L g982 ( .A(n_851), .Y(n_982) );
AND2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_853), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_863), .B1(n_864), .B2(n_871), .Y(n_854) );
INVx1_ASAP7_75t_L g940 ( .A(n_855), .Y(n_940) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_858), .Y(n_855) );
AOI22xp33_ASAP7_75t_SL g874 ( .A1(n_856), .A2(n_875), .B1(n_878), .B2(n_880), .Y(n_874) );
AND2x4_ASAP7_75t_L g875 ( .A(n_856), .B(n_876), .Y(n_875) );
AND2x2_ASAP7_75t_L g914 ( .A(n_856), .B(n_915), .Y(n_914) );
AND2x2_ASAP7_75t_L g927 ( .A(n_856), .B(n_860), .Y(n_927) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
AOI211xp5_ASAP7_75t_L g923 ( .A1(n_858), .A2(n_924), .B(n_925), .C(n_936), .Y(n_923) );
INVx1_ASAP7_75t_L g991 ( .A(n_858), .Y(n_991) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
OR2x2_ASAP7_75t_L g870 ( .A(n_859), .B(n_860), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_859), .B(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g967 ( .A(n_860), .Y(n_967) );
AOI222xp33_ASAP7_75t_L g1015 ( .A1(n_860), .A2(n_884), .B1(n_1016), .B2(n_1017), .C1(n_1019), .C2(n_1020), .Y(n_1015) );
AND2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_867), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_864), .B(n_910), .Y(n_909) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_865), .B(n_921), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_865), .B(n_927), .Y(n_926) );
A2O1A1Ixp33_ASAP7_75t_L g1023 ( .A1(n_865), .A2(n_1024), .B(n_1025), .C(n_1027), .Y(n_1023) );
NOR2xp67_ASAP7_75t_SL g1025 ( .A(n_865), .B(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g978 ( .A(n_866), .B(n_908), .Y(n_978) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx3_ASAP7_75t_SL g873 ( .A(n_870), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_873), .B(n_938), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_873), .A2(n_924), .B1(n_1008), .B2(n_1009), .C(n_1010), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_875), .B(n_902), .Y(n_901) );
INVx2_ASAP7_75t_SL g921 ( .A(n_875), .Y(n_921) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_875), .B(n_903), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_876), .B(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_877), .B(n_957), .Y(n_963) );
AND2x2_ASAP7_75t_L g924 ( .A(n_878), .B(n_907), .Y(n_924) );
AOI321xp33_ASAP7_75t_L g970 ( .A1(n_878), .A2(n_971), .A3(n_972), .B1(n_973), .B2(n_975), .C(n_977), .Y(n_970) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_884), .Y(n_881) );
AND2x2_ASAP7_75t_L g999 ( .A(n_882), .B(n_976), .Y(n_999) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g943 ( .A1(n_883), .A2(n_944), .B1(n_949), .B2(n_950), .C(n_951), .Y(n_943) );
OAI321xp33_ASAP7_75t_L g961 ( .A1(n_883), .A2(n_950), .A3(n_962), .B1(n_964), .B2(n_968), .C(n_970), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_883), .B(n_884), .Y(n_1021) );
AND2x2_ASAP7_75t_L g975 ( .A(n_884), .B(n_976), .Y(n_975) );
INVxp67_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_892), .Y(n_886) );
OAI31xp33_ASAP7_75t_L g899 ( .A1(n_887), .A2(n_900), .A3(n_909), .B(n_912), .Y(n_899) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
AOI211xp5_ASAP7_75t_L g942 ( .A1(n_888), .A2(n_943), .B(n_961), .C(n_980), .Y(n_942) );
AOI222xp33_ASAP7_75t_L g987 ( .A1(n_888), .A2(n_931), .B1(n_988), .B2(n_989), .C1(n_992), .C2(n_997), .Y(n_987) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g974 ( .A(n_889), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_889), .B(n_907), .Y(n_1022) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g908 ( .A(n_895), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
NAND4xp25_ASAP7_75t_L g898 ( .A(n_899), .B(n_942), .C(n_987), .D(n_998), .Y(n_898) );
AOI21xp33_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_904), .B(n_905), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_902), .B(n_914), .Y(n_984) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_903), .B(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g1024 ( .A(n_904), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
INVx2_ASAP7_75t_L g969 ( .A(n_906), .Y(n_969) );
OAI322xp33_ASAP7_75t_L g1010 ( .A1(n_906), .A2(n_957), .A3(n_967), .B1(n_990), .B2(n_1011), .C1(n_1012), .C2(n_1014), .Y(n_1010) );
INVx1_ASAP7_75t_L g997 ( .A(n_907), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_907), .B(n_994), .Y(n_1014) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
BUFx3_ASAP7_75t_L g946 ( .A(n_908), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_908), .B(n_948), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_911), .B(n_914), .Y(n_913) );
AOI321xp33_ASAP7_75t_L g998 ( .A1(n_911), .A2(n_974), .A3(n_982), .B1(n_999), .B2(n_1000), .C(n_1001), .Y(n_998) );
OAI221xp5_ASAP7_75t_SL g912 ( .A1(n_913), .A2(n_916), .B1(n_919), .B2(n_922), .C(n_923), .Y(n_912) );
INVx1_ASAP7_75t_L g949 ( .A(n_914), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_915), .B(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g957 ( .A(n_915), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g1005 ( .A(n_917), .B(n_948), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_918), .B(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g1018 ( .A(n_918), .Y(n_1018) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
O2A1O1Ixp33_ASAP7_75t_L g977 ( .A1(n_922), .A2(n_974), .B(n_978), .C(n_979), .Y(n_977) );
A2O1A1Ixp33_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_928), .B(n_930), .C(n_932), .Y(n_925) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_931), .B(n_969), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
INVx1_ASAP7_75t_L g972 ( .A(n_934), .Y(n_972) );
AOI21xp33_ASAP7_75t_SL g936 ( .A1(n_937), .A2(n_940), .B(n_941), .Y(n_936) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
OR2x2_ASAP7_75t_L g990 ( .A(n_939), .B(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g985 ( .A(n_945), .Y(n_985) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
INVx2_ASAP7_75t_L g960 ( .A(n_946), .Y(n_960) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
AOI21xp33_ASAP7_75t_L g1001 ( .A1(n_949), .A2(n_1002), .B(n_1004), .Y(n_1001) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_955), .B(n_956), .Y(n_951) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_953), .Y(n_952) );
NOR3xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_958), .C(n_960), .Y(n_956) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_969), .B(n_984), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g989 ( .A(n_969), .B(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1011 ( .A(n_971), .Y(n_1011) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g983 ( .A(n_974), .Y(n_983) );
OAI221xp5_ASAP7_75t_SL g1006 ( .A1(n_974), .A2(n_1007), .B1(n_1015), .B2(n_1022), .C(n_1023), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_980) );
INVxp67_ASAP7_75t_L g1027 ( .A(n_981), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
CKINVDCx14_ASAP7_75t_R g1013 ( .A(n_982), .Y(n_1013) );
INVx1_ASAP7_75t_L g1016 ( .A(n_986), .Y(n_1016) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_995), .Y(n_993) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
CKINVDCx14_ASAP7_75t_R g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVxp67_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
NOR2x1_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1042), .Y(n_1033) );
NAND4xp25_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .C(n_1037), .D(n_1040), .Y(n_1034) );
NAND4xp25_ASAP7_75t_SL g1042 ( .A(n_1043), .B(n_1045), .C(n_1046), .D(n_1047), .Y(n_1042) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
NOR4xp75_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1063), .C(n_1067), .D(n_1071), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1062), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1066), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1070), .Y(n_1067) );
NAND2xp5_ASAP7_75t_SL g1071 ( .A(n_1072), .B(n_1074), .Y(n_1071) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g1079 ( .A(n_1080), .Y(n_1079) );
endmodule