module fake_jpeg_2864_n_204 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_52),
.B1(n_71),
.B2(n_63),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_69),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_62),
.C(n_48),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_88),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_62),
.C(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_52),
.B1(n_71),
.B2(n_66),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_51),
.B1(n_60),
.B2(n_69),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_95),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_93),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_68),
.B(n_64),
.C(n_67),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_52),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_61),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_60),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_123),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_56),
.B(n_61),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_126),
.B(n_12),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_0),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_23),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_70),
.B(n_22),
.C(n_25),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_70),
.B1(n_2),
.B2(n_4),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_101),
.B(n_8),
.C(n_9),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_7),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_155),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_98),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

AO21x2_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_30),
.B(n_47),
.Y(n_146)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_128),
.B1(n_36),
.B2(n_27),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_29),
.C(n_46),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_154),
.C(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_7),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

OA21x2_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_10),
.B(n_11),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_10),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_120),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_156),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_14),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_133),
.B1(n_126),
.B2(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_169),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_174),
.B1(n_141),
.B2(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_146),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_35),
.C(n_45),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_147),
.C(n_155),
.Y(n_184)
);

XOR2x1_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_17),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_177),
.B(n_179),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_135),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_184),
.Y(n_186)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_185),
.B(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_162),
.Y(n_183)
);

OA21x2_ASAP7_75t_SL g188 ( 
.A1(n_183),
.A2(n_161),
.B(n_163),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_176),
.A3(n_166),
.B1(n_168),
.B2(n_165),
.C1(n_174),
.C2(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_189),
.A2(n_178),
.B1(n_164),
.B2(n_184),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_167),
.C(n_171),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_39),
.B(n_31),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_141),
.C(n_164),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_192),
.A2(n_141),
.B(n_190),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_196),
.B(n_32),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_186),
.C(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_187),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_34),
.Y(n_203)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_203),
.Y(n_204)
);


endmodule