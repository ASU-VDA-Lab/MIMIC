module fake_jpeg_2661_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_42),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_8),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_0),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_66),
.B1(n_51),
.B2(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_62),
.Y(n_86)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_58),
.B1(n_56),
.B2(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_79),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_62),
.B1(n_57),
.B2(n_59),
.Y(n_81)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_67),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_106),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_96),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_71),
.B(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_99),
.C(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_50),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_73),
.C(n_68),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_73),
.C(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_49),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_25),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_51),
.B1(n_49),
.B2(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_115),
.B1(n_105),
.B2(n_65),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_64),
.B1(n_65),
.B2(n_5),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_4),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_7),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_119),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_8),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_26),
.Y(n_123)
);

XOR2x2_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_9),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_94),
.C(n_91),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_138),
.C(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_140),
.Y(n_151)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_27),
.C(n_43),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_65),
.B(n_11),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_143),
.B(n_14),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_22),
.C(n_35),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_10),
.B(n_11),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_12),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_145),
.B(n_13),
.Y(n_149)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_16),
.Y(n_152)
);

AO221x1_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_152),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_18),
.B1(n_20),
.B2(n_28),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_127),
.B1(n_141),
.B2(n_134),
.Y(n_171)
);

XOR2x1_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_29),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_30),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_32),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_142),
.C(n_143),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_33),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_171),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_151),
.B(n_126),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_165),
.B1(n_166),
.B2(n_153),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_162),
.B(n_150),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_170),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_174),
.A2(n_163),
.B(n_156),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_158),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_177),
.B(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_182),
.B1(n_175),
.B2(n_170),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_180),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_189),
.A2(n_190),
.B(n_188),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_186),
.C(n_159),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_159),
.Y(n_193)
);


endmodule