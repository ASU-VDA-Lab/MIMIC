module real_jpeg_29914_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g103 ( 
.A(n_0),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_0),
.Y(n_108)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_0),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_27),
.B1(n_31),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_1),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_118),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_118),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_59),
.B1(n_61),
.B2(n_118),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_2),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_26),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_2),
.B(n_31),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_2),
.A2(n_31),
.B(n_165),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_123),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_56),
.B(n_59),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_2),
.B(n_78),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_100),
.B1(n_103),
.B2(n_216),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_4),
.A2(n_22),
.B1(n_25),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_4),
.A2(n_48),
.B1(n_59),
.B2(n_61),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_4),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_4),
.A2(n_27),
.B1(n_31),
.B2(n_48),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_7),
.A2(n_22),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_7),
.A2(n_27),
.B1(n_31),
.B2(n_37),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_7),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_37),
.B1(n_59),
.B2(n_61),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_8),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_120),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_8),
.A2(n_59),
.B1(n_61),
.B2(n_120),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_8),
.A2(n_22),
.B1(n_25),
.B2(n_120),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_9),
.A2(n_24),
.B1(n_53),
.B2(n_54),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_24),
.B1(n_27),
.B2(n_31),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_9),
.A2(n_24),
.B1(n_59),
.B2(n_61),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_10),
.A2(n_22),
.B1(n_25),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_10),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_10),
.A2(n_46),
.B1(n_59),
.B2(n_61),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_10),
.A2(n_27),
.B1(n_31),
.B2(n_46),
.Y(n_273)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_12),
.A2(n_22),
.B1(n_25),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_12),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_12),
.A2(n_27),
.B1(n_31),
.B2(n_125),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_125),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_12),
.A2(n_59),
.B1(n_61),
.B2(n_125),
.Y(n_216)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_15),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_85),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_83),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_20),
.A2(n_44),
.B(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_21),
.A2(n_33),
.B(n_82),
.Y(n_300)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_26),
.B(n_29),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_29),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g122 ( 
.A(n_22),
.B(n_123),
.CON(n_122),
.SN(n_122)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_26),
.A2(n_33),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_31),
.B1(n_68),
.B2(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_27),
.A2(n_34),
.B1(n_122),
.B2(n_137),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_53),
.A3(n_67),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_29),
.B(n_31),
.Y(n_137)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_32),
.A2(n_45),
.B(n_49),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_33),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_75),
.C(n_80),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_40),
.A2(n_41),
.B1(n_337),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.C(n_64),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_42),
.A2(n_43),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_44),
.A2(n_49),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_44),
.A2(n_49),
.B1(n_131),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_50),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_50),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_50),
.A2(n_64),
.B1(n_309),
.B2(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_58),
.B(n_62),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_51),
.A2(n_62),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_51),
.A2(n_58),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_51),
.A2(n_173),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_51),
.A2(n_58),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_51),
.A2(n_58),
.B1(n_172),
.B2(n_191),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_51),
.A2(n_58),
.B1(n_95),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_51),
.A2(n_113),
.B(n_249),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_54),
.B(n_68),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_54),
.A2(n_57),
.B(n_123),
.C(n_193),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_58),
.B(n_123),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_59),
.Y(n_61)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_61),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_63),
.B(n_114),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_64),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_65),
.A2(n_77),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_66),
.A2(n_73),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_66),
.A2(n_73),
.B1(n_117),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_66),
.A2(n_73),
.B1(n_148),
.B2(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_66),
.B(n_72),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_66),
.A2(n_73),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_71),
.A2(n_78),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_77),
.A2(n_79),
.B(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_77),
.A2(n_259),
.B(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_80),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_334),
.B(n_340),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_304),
.A3(n_326),
.B1(n_332),
.B2(n_333),
.C(n_342),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_285),
.B(n_303),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_263),
.B(n_284),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_155),
.B(n_240),
.C(n_262),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_140),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_91),
.B(n_140),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_126),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_110),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_93),
.B(n_110),
.C(n_126),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_94),
.B(n_99),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_96),
.B(n_183),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B(n_105),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_100),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_100),
.A2(n_208),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_100),
.A2(n_152),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_101),
.A2(n_106),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_101),
.A2(n_203),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_121),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_123),
.B(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_128),
.B(n_133),
.C(n_135),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_138),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_141),
.A2(n_142),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_151),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_153),
.B(n_202),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_239),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_232),
.B(n_238),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_184),
.B(n_231),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_174),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_159),
.B(n_174),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.C(n_170),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_160),
.A2(n_161),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_163),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_181),
.C(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_225),
.B(n_230),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_204),
.B(n_224),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_194),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_194),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_199),
.C(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_201),
.Y(n_209)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_212),
.B(n_223),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_210),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_218),
.B(n_222),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_214),
.B(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_260),
.B2(n_261),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_251),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_251),
.C(n_261),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_254),
.C(n_258),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_283),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_276),
.B2(n_277),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_277),
.C(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_272),
.C(n_274),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_278),
.A2(n_279),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_281),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_297),
.B(n_300),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_287),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_301),
.B2(n_302),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_296),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_296),
.C(n_302),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B(n_295),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_294),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_306),
.C(n_316),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_295),
.A2(n_306),
.B1(n_307),
.B2(n_331),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_295),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_318),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_318),
.Y(n_333)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_311),
.C(n_313),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_313),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_315),
.B1(n_320),
.B2(n_324),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_324),
.C(n_325),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_316),
.A2(n_317),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_325),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.Y(n_340)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);


endmodule