module fake_jpeg_19070_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_19),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_3),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_0),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_45),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_76),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_52),
.B1(n_64),
.B2(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_83),
.B1(n_85),
.B2(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_4),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_65),
.C(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_50),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_56),
.B1(n_62),
.B2(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_46),
.Y(n_87)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_1),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_6),
.C(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_92),
.Y(n_101)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_60),
.B1(n_51),
.B2(n_4),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_5),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_102),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_107),
.B1(n_9),
.B2(n_13),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_16),
.B(n_17),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_58),
.B1(n_10),
.B2(n_11),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.C(n_113),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_26),
.B(n_29),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_99),
.C(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_116),
.B(n_104),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_36),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_38),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_40),
.C(n_42),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_106),
.Y(n_127)
);


endmodule