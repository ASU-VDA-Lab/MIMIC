module fake_jpeg_9117_n_57 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_57);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_57;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_23),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_32),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_9),
.B1(n_20),
.B2(n_19),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_35),
.B1(n_4),
.B2(n_5),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_34),
.B(n_36),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_1),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_44),
.B1(n_45),
.B2(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_41),
.B1(n_4),
.B2(n_5),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_29),
.C(n_28),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_11),
.B1(n_18),
.B2(n_14),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_8),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_6),
.B1(n_7),
.B2(n_22),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_50),
.Y(n_54)
);

A2O1A1O1Ixp25_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_53),
.B(n_43),
.C(n_51),
.D(n_42),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_42),
.C(n_48),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_40),
.CI(n_45),
.CON(n_57),
.SN(n_57)
);


endmodule