module fake_jpeg_11201_n_196 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_196);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_27),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx3_ASAP7_75t_SL g75 ( 
.A(n_2),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_89),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_1),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_1),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_95),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_107),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_104),
.B1(n_108),
.B2(n_83),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_82),
.B1(n_75),
.B2(n_57),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_75),
.B1(n_82),
.B2(n_78),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_115),
.B1(n_124),
.B2(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_83),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_122),
.C(n_4),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_121),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_84),
.B1(n_61),
.B2(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_64),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_85),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_69),
.C(n_67),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_73),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_70),
.B1(n_79),
.B2(n_81),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_60),
.B(n_76),
.C(n_62),
.Y(n_127)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_57),
.B1(n_60),
.B2(n_65),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_76),
.B1(n_62),
.B2(n_65),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_144),
.B1(n_150),
.B2(n_14),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_3),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_138),
.B(n_143),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_10),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_4),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_5),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_8),
.B(n_9),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_149),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_12),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_40),
.C(n_15),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_164),
.C(n_166),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_16),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_134),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_17),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_54),
.C(n_22),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_38),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_140),
.B(n_162),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_174),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_157),
.B(n_156),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_152),
.C(n_41),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_169),
.C(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_184),
.B(n_176),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_156),
.C(n_170),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_189),
.A2(n_180),
.B1(n_183),
.B2(n_178),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_190),
.A2(n_180),
.B1(n_165),
.B2(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_39),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_42),
.C(n_43),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_47),
.C(n_49),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_50),
.B(n_51),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_53),
.Y(n_196)
);


endmodule