module fake_jpeg_24792_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_30),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_1),
.Y(n_30)
);

CKINVDCx9p33_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_13),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_18),
.B1(n_14),
.B2(n_15),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_17),
.B1(n_20),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_18),
.B1(n_14),
.B2(n_15),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_35),
.B1(n_43),
.B2(n_28),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_13),
.B1(n_20),
.B2(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_9),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_26),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_53),
.C(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_57),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_56),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_24),
.B1(n_19),
.B2(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_25),
.C(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_22),
.B1(n_31),
.B2(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_69),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_57),
.B1(n_45),
.B2(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_58),
.B1(n_50),
.B2(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_79),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_50),
.B1(n_47),
.B2(n_40),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_39),
.Y(n_79)
);

XOR2x2_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_39),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_64),
.C(n_65),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_36),
.B1(n_3),
.B2(n_2),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.C(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_65),
.C(n_60),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_90),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_78),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_93),
.Y(n_97)
);

AO221x1_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_77),
.B1(n_3),
.B2(n_74),
.C(n_8),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_86),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_91),
.C(n_94),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_87),
.B(n_95),
.C(n_67),
.D(n_66),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_66),
.C(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_102),
.Y(n_105)
);


endmodule