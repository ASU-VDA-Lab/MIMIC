module fake_jpeg_5932_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_6),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_4),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_23),
.C(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_0),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_28),
.B(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_10),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_1),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_18),
.C(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_15),
.B(n_2),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_13),
.C(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_29),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_24),
.C(n_21),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_17),
.B1(n_19),
.B2(n_18),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_40),
.B1(n_24),
.B2(n_26),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_12),
.C(n_17),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_38),
.C(n_23),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_39),
.B(n_24),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_16),
.B1(n_20),
.B2(n_4),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_21),
.C(n_28),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_20),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_33),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_29),
.B(n_3),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVxp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_32),
.B(n_29),
.C(n_4),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_41),
.C(n_32),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

BUFx24_ASAP7_75t_SL g58 ( 
.A(n_53),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_62),
.B(n_8),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_2),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_50),
.B(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_65),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_51),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_2),
.B(n_3),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_SL g68 ( 
.A1(n_67),
.A2(n_3),
.B(n_5),
.C(n_64),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_5),
.B1(n_63),
.B2(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_70),
.B1(n_64),
.B2(n_66),
.Y(n_72)
);


endmodule