module fake_netlist_6_4537_n_157 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_29, n_25, n_157);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_157;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_145;
wire n_92;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_130;
wire n_78;
wire n_99;
wire n_84;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_30),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

OR2x6_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_0),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_R g61 ( 
.A(n_40),
.B(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_30),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_32),
.B(n_6),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_32),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_8),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_45),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_48),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_47),
.C(n_41),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_48),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_46),
.B(n_53),
.C(n_43),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_10),
.C(n_11),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

AOI221xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_71),
.B1(n_63),
.B2(n_67),
.C(n_74),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_72),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_66),
.Y(n_95)
);

CKINVDCx11_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_70),
.C(n_57),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_72),
.B(n_70),
.Y(n_98)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_66),
.B(n_65),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

OAI21x1_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_78),
.B(n_88),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_87),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_78),
.B(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_81),
.Y(n_107)
);

OR2x6_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_85),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_85),
.B(n_90),
.Y(n_110)
);

NOR2x1_ASAP7_75t_R g111 ( 
.A(n_107),
.B(n_96),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_68),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_93),
.B1(n_80),
.B2(n_75),
.C(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_101),
.B(n_110),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_102),
.B(n_101),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_115),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_113),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_113),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_113),
.Y(n_128)
);

OR2x6_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_114),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_116),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_108),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_108),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_93),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_61),
.B1(n_130),
.B2(n_129),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_129),
.B(n_57),
.C(n_127),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_129),
.B(n_101),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_111),
.B1(n_62),
.B2(n_60),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_62),
.B(n_55),
.C(n_123),
.Y(n_140)
);

AOI222xp33_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_100),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_99),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_23),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_140),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_141),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_92),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_92),
.B1(n_102),
.B2(n_84),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_84),
.Y(n_151)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_152),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_152),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_150),
.B1(n_153),
.B2(n_155),
.Y(n_157)
);


endmodule