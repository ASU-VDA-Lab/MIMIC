module fake_aes_7581_n_1355 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1355);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1355;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g294 ( .A(n_172), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_55), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_47), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_224), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_197), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_246), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_202), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_250), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_289), .Y(n_302) );
NOR2xp67_ASAP7_75t_L g303 ( .A(n_184), .B(n_140), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_118), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_151), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_30), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_56), .Y(n_307) );
BUFx5_ASAP7_75t_L g308 ( .A(n_86), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_109), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_174), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_188), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_193), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_226), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_72), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_169), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_288), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_154), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_210), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_36), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_83), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_80), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_279), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_278), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_139), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_103), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_30), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_235), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_266), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_247), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_106), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_131), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_41), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_102), .B(n_213), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_11), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_113), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_138), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_9), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_97), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_248), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_68), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_82), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_168), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_293), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_6), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_272), .Y(n_346) );
CKINVDCx16_ASAP7_75t_R g347 ( .A(n_205), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_40), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_71), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_208), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_276), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_17), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_243), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_123), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_155), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_115), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_229), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_206), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_263), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_136), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_236), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_50), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_286), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_252), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_201), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_273), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_170), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_231), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_177), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_15), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_86), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_41), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_70), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_0), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_187), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_142), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_260), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_83), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_285), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_251), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_28), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_104), .B(n_7), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_0), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_261), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_274), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_36), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_215), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_173), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_183), .Y(n_389) );
BUFx8_ASAP7_75t_SL g390 ( .A(n_284), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_62), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_232), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_62), .Y(n_393) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_18), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_124), .Y(n_395) );
BUFx5_ASAP7_75t_L g396 ( .A(n_73), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_204), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_75), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_161), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_269), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_84), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_163), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_217), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_262), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_287), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_190), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_121), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_264), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_171), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_141), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_52), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_56), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_58), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_98), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_92), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_176), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_58), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_162), .Y(n_418) );
INVxp33_ASAP7_75t_L g419 ( .A(n_110), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_186), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_245), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_132), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_19), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_258), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_240), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_53), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_66), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_189), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_158), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_153), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_192), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_181), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_209), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_165), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_79), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_195), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_167), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_283), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_111), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_244), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_3), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_280), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_42), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_191), .Y(n_444) );
INVxp67_ASAP7_75t_L g445 ( .A(n_35), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_255), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_6), .Y(n_447) );
CKINVDCx14_ASAP7_75t_R g448 ( .A(n_218), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_39), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_296), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_308), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_413), .A2(n_4), .B1(n_1), .B2(n_2), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_332), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_308), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_332), .B(n_4), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_427), .B(n_5), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_332), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_308), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_419), .B(n_5), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_332), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_308), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_444), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_296), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_463) );
NAND2xp33_ASAP7_75t_L g464 ( .A(n_308), .B(n_93), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_321), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_465) );
NOR2xp33_ASAP7_75t_R g466 ( .A(n_448), .B(n_94), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_427), .B(n_10), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_390), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_333), .B(n_12), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_321), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_444), .Y(n_471) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_325), .A2(n_96), .B(n_95), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_308), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_308), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_333), .B(n_12), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_396), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_327), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_477) );
AND2x6_ASAP7_75t_L g478 ( .A(n_329), .B(n_99), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_444), .Y(n_479) );
CKINVDCx6p67_ASAP7_75t_R g480 ( .A(n_347), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_396), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_396), .Y(n_484) );
CKINVDCx6p67_ASAP7_75t_R g485 ( .A(n_329), .Y(n_485) );
AND2x6_ASAP7_75t_L g486 ( .A(n_416), .B(n_100), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_457), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_459), .B(n_419), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_456), .B(n_325), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_459), .B(n_448), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_478), .Y(n_492) );
AND2x6_ASAP7_75t_L g493 ( .A(n_456), .B(n_416), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_470), .B(n_480), .Y(n_494) );
INVx4_ASAP7_75t_L g495 ( .A(n_478), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_480), .B(n_396), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_451), .B(n_353), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_473), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_485), .B(n_357), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_456), .B(n_396), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_454), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_456), .B(n_396), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_458), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_478), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_458), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_461), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_478), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_461), .B(n_353), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_457), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_467), .B(n_348), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_476), .B(n_481), .Y(n_512) );
XOR2xp5_ASAP7_75t_L g513 ( .A(n_468), .B(n_413), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_485), .B(n_387), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_457), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_467), .A2(n_326), .B1(n_331), .B2(n_313), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_476), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_478), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_457), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_467), .B(n_348), .Y(n_520) );
BUFx3_ASAP7_75t_L g521 ( .A(n_478), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_467), .B(n_360), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_457), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_457), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_484), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_478), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_481), .B(n_360), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_460), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_482), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_486), .Y(n_530) );
INVx4_ASAP7_75t_SL g531 ( .A(n_486), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_482), .B(n_366), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_473), .B(n_366), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_484), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_460), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_468), .B(n_449), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_525), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_495), .B(n_466), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_493), .A2(n_475), .B1(n_469), .B2(n_486), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_492), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_489), .B(n_469), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_496), .B(n_469), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_500), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_489), .B(n_469), .Y(n_544) );
NAND2xp33_ASAP7_75t_SL g545 ( .A(n_495), .B(n_313), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_495), .B(n_475), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_491), .B(n_475), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_493), .Y(n_548) );
OR2x6_ASAP7_75t_L g549 ( .A(n_491), .B(n_452), .Y(n_549) );
BUFx3_ASAP7_75t_L g550 ( .A(n_492), .Y(n_550) );
AND2x6_ASAP7_75t_SL g551 ( .A(n_513), .B(n_452), .Y(n_551) );
OR2x6_ASAP7_75t_L g552 ( .A(n_491), .B(n_465), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_495), .B(n_300), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_500), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_496), .B(n_300), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_525), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_496), .B(n_327), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_492), .Y(n_558) );
NOR2x2_ASAP7_75t_L g559 ( .A(n_513), .B(n_390), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_525), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_500), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_511), .B(n_301), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_536), .B(n_335), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_525), .Y(n_564) );
NOR2x1p5_ASAP7_75t_L g565 ( .A(n_494), .B(n_335), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_536), .B(n_386), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_525), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_511), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_492), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_534), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_503), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_520), .B(n_312), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_494), .Y(n_573) );
AO22x1_ASAP7_75t_L g574 ( .A1(n_493), .A2(n_486), .B1(n_477), .B2(n_377), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_495), .B(n_312), .Y(n_575) );
NOR2x1p5_ASAP7_75t_L g576 ( .A(n_494), .B(n_386), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_503), .B(n_450), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_503), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_487), .A2(n_472), .B(n_486), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_520), .B(n_317), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_513), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_493), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_516), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_520), .B(n_317), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_536), .A2(n_326), .B1(n_415), .B2(n_331), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_495), .B(n_330), .Y(n_586) );
NOR2x2_ASAP7_75t_L g587 ( .A(n_516), .B(n_415), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_490), .A2(n_431), .B1(n_424), .B2(n_450), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_493), .A2(n_431), .B1(n_424), .B2(n_393), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_493), .A2(n_486), .B1(n_474), .B2(n_484), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_518), .B(n_330), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_493), .B(n_343), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_518), .B(n_343), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_534), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_505), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_493), .A2(n_295), .B1(n_314), .B2(n_306), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_493), .A2(n_322), .B1(n_338), .B2(n_320), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_534), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_499), .B(n_392), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_499), .B(n_356), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_497), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_497), .Y(n_602) );
INVxp67_ASAP7_75t_SL g603 ( .A(n_505), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_514), .B(n_356), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_490), .A2(n_342), .B1(n_345), .B2(n_341), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_522), .A2(n_352), .B1(n_362), .B2(n_349), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_522), .A2(n_463), .B1(n_514), .B2(n_518), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_533), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_518), .A2(n_393), .B1(n_417), .B2(n_394), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_505), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_509), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_498), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_518), .B(n_404), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_509), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_533), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_498), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_512), .Y(n_617) );
AND2x4_ASAP7_75t_SL g618 ( .A(n_518), .B(n_463), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_530), .A2(n_371), .B1(n_373), .B2(n_370), .Y(n_619) );
INVx3_ASAP7_75t_L g620 ( .A(n_530), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_512), .B(n_407), .Y(n_621) );
INVx3_ASAP7_75t_L g622 ( .A(n_530), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_530), .A2(n_374), .B1(n_381), .B2(n_378), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_487), .B(n_407), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_501), .Y(n_625) );
INVxp33_ASAP7_75t_L g626 ( .A(n_527), .Y(n_626) );
AO22x1_ASAP7_75t_L g627 ( .A1(n_530), .A2(n_311), .B1(n_425), .B2(n_417), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_501), .Y(n_628) );
INVx4_ASAP7_75t_L g629 ( .A(n_530), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_501), .B(n_425), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_502), .B(n_337), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_531), .B(n_391), .Y(n_632) );
BUFx3_ASAP7_75t_L g633 ( .A(n_505), .Y(n_633) );
INVx5_ASAP7_75t_L g634 ( .A(n_508), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_531), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_508), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_540), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_614), .B(n_508), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_617), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_617), .B(n_502), .Y(n_640) );
OAI22x1_ASAP7_75t_L g641 ( .A1(n_585), .A2(n_307), .B1(n_445), .B2(n_372), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_601), .B(n_502), .Y(n_642) );
BUFx3_ASAP7_75t_L g643 ( .A(n_563), .Y(n_643) );
AO21x1_ASAP7_75t_L g644 ( .A1(n_579), .A2(n_464), .B(n_527), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_602), .B(n_504), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_577), .A2(n_398), .B1(n_401), .B2(n_411), .C1(n_412), .C2(n_423), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_588), .B(n_455), .C(n_435), .Y(n_647) );
NOR2xp33_ASAP7_75t_R g648 ( .A(n_545), .B(n_521), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_563), .B(n_426), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_611), .A2(n_532), .B(n_526), .C(n_521), .Y(n_650) );
OR2x6_ASAP7_75t_L g651 ( .A(n_549), .B(n_521), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_568), .B(n_531), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_543), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_608), .B(n_504), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_615), .A2(n_526), .B1(n_506), .B2(n_507), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_554), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_581), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_607), .A2(n_532), .B(n_506), .C(n_507), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_566), .B(n_441), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_577), .A2(n_504), .B1(n_517), .B2(n_507), .Y(n_660) );
BUFx12f_ASAP7_75t_L g661 ( .A(n_551), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_573), .B(n_517), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_549), .A2(n_552), .B1(n_583), .B2(n_615), .Y(n_663) );
NAND3xp33_ASAP7_75t_SL g664 ( .A(n_589), .B(n_421), .C(n_350), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_554), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_542), .B(n_529), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_542), .B(n_529), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_545), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_570), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_625), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_557), .B(n_566), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_542), .B(n_561), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_610), .A2(n_539), .B1(n_577), .B2(n_618), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_548), .B(n_531), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_549), .A2(n_447), .B1(n_443), .B2(n_383), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_549), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_628), .A2(n_382), .B(n_443), .C(n_383), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_628), .A2(n_472), .B(n_531), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_540), .Y(n_679) );
BUFx8_ASAP7_75t_L g680 ( .A(n_557), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_561), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_541), .A2(n_449), .B(n_418), .C(n_406), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_571), .B(n_531), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_546), .A2(n_472), .B(n_531), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_547), .A2(n_297), .B(n_294), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_544), .A2(n_299), .B(n_298), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_627), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_570), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_627), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_583), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_540), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_571), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_594), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_578), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_613), .A2(n_382), .B(n_304), .C(n_305), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_540), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_619), .B(n_447), .C(n_309), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_631), .A2(n_310), .B(n_302), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_552), .B(n_315), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_565), .B(n_447), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_562), .B(n_447), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_576), .Y(n_702) );
AOI21x1_ASAP7_75t_L g703 ( .A1(n_574), .A2(n_510), .B(n_488), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_598), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_L g705 ( .A1(n_572), .A2(n_316), .B(n_319), .C(n_318), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_552), .B(n_323), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_552), .B(n_13), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_538), .A2(n_328), .B(n_324), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_553), .A2(n_339), .B(n_336), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_610), .A2(n_340), .B1(n_346), .B2(n_344), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_612), .Y(n_711) );
NOR2xp33_ASAP7_75t_R g712 ( .A(n_582), .B(n_14), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_580), .B(n_351), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_623), .B(n_355), .C(n_354), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_575), .A2(n_359), .B(n_358), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_548), .B(n_361), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_618), .A2(n_363), .B1(n_365), .B2(n_364), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_586), .A2(n_368), .B(n_367), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_574), .A2(n_369), .B1(n_376), .B2(n_375), .Y(n_719) );
BUFx2_ASAP7_75t_L g720 ( .A(n_559), .Y(n_720) );
NOR2x1_ASAP7_75t_R g721 ( .A(n_559), .B(n_379), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_621), .A2(n_380), .B1(n_385), .B2(n_384), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_584), .B(n_388), .Y(n_723) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_587), .A2(n_397), .B1(n_399), .B2(n_395), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_591), .A2(n_402), .B(n_400), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_616), .A2(n_405), .B(n_408), .C(n_403), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_593), .A2(n_410), .B(n_409), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_609), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_596), .A2(n_428), .B1(n_429), .B2(n_422), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_555), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_590), .A2(n_433), .B(n_432), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_624), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_600), .Y(n_733) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_630), .A2(n_436), .B(n_437), .C(n_434), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_632), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_605), .B(n_438), .Y(n_736) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_550), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_606), .B(n_439), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_558), .A2(n_446), .B(n_442), .Y(n_739) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_540), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_604), .B(n_389), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_599), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g743 ( .A1(n_537), .A2(n_414), .B(n_389), .Y(n_743) );
OAI21xp33_ASAP7_75t_L g744 ( .A1(n_597), .A2(n_420), .B(n_414), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_634), .B(n_420), .Y(n_745) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_587), .A2(n_430), .B1(n_440), .B2(n_334), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_634), .B(n_430), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_592), .B(n_440), .Y(n_748) );
BUFx3_ASAP7_75t_L g749 ( .A(n_537), .Y(n_749) );
INVx5_ASAP7_75t_L g750 ( .A(n_582), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_626), .B(n_16), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_556), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_582), .B(n_16), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_556), .Y(n_754) );
INVx2_ASAP7_75t_SL g755 ( .A(n_560), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_603), .A2(n_303), .B1(n_334), .B2(n_453), .Y(n_756) );
O2A1O1Ixp33_ASAP7_75t_L g757 ( .A1(n_564), .A2(n_453), .B(n_462), .C(n_483), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_564), .B(n_18), .Y(n_758) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_550), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_567), .B(n_19), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_567), .Y(n_761) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_633), .Y(n_762) );
AO31x2_ASAP7_75t_L g763 ( .A1(n_629), .A2(n_453), .A3(n_462), .B(n_483), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_635), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_629), .B(n_20), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_569), .A2(n_510), .B(n_488), .Y(n_766) );
INVx5_ASAP7_75t_L g767 ( .A(n_634), .Y(n_767) );
BUFx12f_ASAP7_75t_L g768 ( .A(n_634), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g769 ( .A(n_634), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_569), .A2(n_510), .B(n_488), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_620), .A2(n_460), .B1(n_471), .B2(n_479), .Y(n_771) );
AOI22x1_ASAP7_75t_SL g772 ( .A1(n_622), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_622), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_622), .B(n_22), .Y(n_774) );
INVx3_ASAP7_75t_L g775 ( .A(n_633), .Y(n_775) );
OAI21x1_ASAP7_75t_L g776 ( .A1(n_636), .A2(n_519), .B(n_515), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_660), .B(n_636), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_680), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_660), .B(n_636), .Y(n_779) );
O2A1O1Ixp5_ASAP7_75t_L g780 ( .A1(n_644), .A2(n_523), .B(n_535), .C(n_528), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_643), .B(n_23), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_L g782 ( .A1(n_695), .A2(n_595), .B(n_535), .C(n_528), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_640), .A2(n_460), .B1(n_471), .B2(n_479), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_639), .B(n_24), .Y(n_784) );
BUFx2_ASAP7_75t_L g785 ( .A(n_680), .Y(n_785) );
INVx2_ASAP7_75t_SL g786 ( .A(n_707), .Y(n_786) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_678), .A2(n_519), .B(n_515), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_663), .A2(n_460), .B1(n_471), .B2(n_479), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_684), .A2(n_519), .B(n_515), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_654), .A2(n_524), .B(n_523), .Y(n_790) );
INVxp67_ASAP7_75t_L g791 ( .A(n_671), .Y(n_791) );
NOR2xp67_ASAP7_75t_SL g792 ( .A(n_687), .B(n_24), .Y(n_792) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_642), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_653), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_657), .B(n_25), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_742), .B(n_25), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_768), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_703), .A2(n_524), .B(n_523), .Y(n_798) );
BUFx3_ASAP7_75t_L g799 ( .A(n_720), .Y(n_799) );
OAI211xp5_ASAP7_75t_L g800 ( .A1(n_675), .A2(n_479), .B(n_471), .C(n_28), .Y(n_800) );
OAI22x1_ASAP7_75t_L g801 ( .A1(n_676), .A2(n_26), .B1(n_27), .B2(n_29), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_645), .A2(n_479), .B1(n_471), .B2(n_29), .Y(n_802) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_637), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_730), .B(n_26), .Y(n_804) );
O2A1O1Ixp33_ASAP7_75t_SL g805 ( .A1(n_753), .A2(n_150), .B(n_292), .C(n_291), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_732), .A2(n_471), .B(n_479), .C(n_32), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_673), .A2(n_27), .B1(n_31), .B2(n_32), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_656), .Y(n_808) );
INVx1_ASAP7_75t_SL g809 ( .A(n_690), .Y(n_809) );
BUFx3_ASAP7_75t_L g810 ( .A(n_702), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_719), .A2(n_31), .B1(n_33), .B2(n_34), .Y(n_811) );
O2A1O1Ixp33_ASAP7_75t_L g812 ( .A1(n_726), .A2(n_33), .B(n_34), .C(n_35), .Y(n_812) );
A2O1A1Ixp33_ASAP7_75t_L g813 ( .A1(n_658), .A2(n_37), .B(n_38), .C(n_39), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_665), .Y(n_814) );
A2O1A1Ixp33_ASAP7_75t_L g815 ( .A1(n_705), .A2(n_37), .B(n_38), .C(n_40), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_766), .A2(n_105), .B(n_101), .Y(n_816) );
AO32x2_ASAP7_75t_L g817 ( .A1(n_756), .A2(n_42), .A3(n_43), .B1(n_44), .B2(n_45), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_770), .A2(n_108), .B(n_107), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_685), .A2(n_114), .B(n_112), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_646), .B(n_43), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_L g821 ( .A1(n_734), .A2(n_44), .B(n_45), .C(n_46), .Y(n_821) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_637), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_699), .B(n_46), .Y(n_823) );
AOI221xp5_ASAP7_75t_L g824 ( .A1(n_746), .A2(n_47), .B1(n_48), .B2(n_49), .C(n_50), .Y(n_824) );
O2A1O1Ixp33_ASAP7_75t_L g825 ( .A1(n_682), .A2(n_48), .B(n_49), .C(n_51), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_669), .Y(n_826) );
BUFx3_ASAP7_75t_L g827 ( .A(n_767), .Y(n_827) );
OAI22xp5_ASAP7_75t_SL g828 ( .A1(n_724), .A2(n_51), .B1(n_52), .B2(n_53), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_706), .B(n_54), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_651), .B(n_54), .Y(n_830) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_647), .B(n_55), .C(n_57), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_743), .A2(n_166), .B(n_282), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g833 ( .A1(n_728), .A2(n_57), .B1(n_59), .B2(n_60), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_681), .Y(n_834) );
INVx3_ASAP7_75t_L g835 ( .A(n_767), .Y(n_835) );
AO21x2_ASAP7_75t_L g836 ( .A1(n_731), .A2(n_164), .B(n_277), .Y(n_836) );
O2A1O1Ixp33_ASAP7_75t_L g837 ( .A1(n_717), .A2(n_59), .B(n_60), .C(n_61), .Y(n_837) );
A2O1A1Ixp33_ASAP7_75t_L g838 ( .A1(n_698), .A2(n_61), .B(n_63), .C(n_64), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_649), .B(n_63), .Y(n_839) );
AO31x2_ASAP7_75t_L g840 ( .A1(n_670), .A2(n_64), .A3(n_65), .B(n_66), .Y(n_840) );
O2A1O1Ixp33_ASAP7_75t_L g841 ( .A1(n_722), .A2(n_65), .B(n_67), .C(n_68), .Y(n_841) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_637), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_655), .A2(n_178), .B(n_275), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_672), .B(n_67), .Y(n_844) );
O2A1O1Ixp33_ASAP7_75t_L g845 ( .A1(n_713), .A2(n_69), .B(n_70), .C(n_71), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_669), .Y(n_846) );
NOR2xp67_ASAP7_75t_SL g847 ( .A(n_689), .B(n_69), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_746), .A2(n_72), .B1(n_73), .B2(n_74), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_692), .Y(n_849) );
A2O1A1Ixp33_ASAP7_75t_L g850 ( .A1(n_686), .A2(n_74), .B(n_75), .C(n_76), .Y(n_850) );
AOI21xp33_ASAP7_75t_L g851 ( .A1(n_662), .A2(n_76), .B(n_77), .Y(n_851) );
NOR2xp33_ASAP7_75t_SL g852 ( .A(n_721), .B(n_77), .Y(n_852) );
CKINVDCx8_ASAP7_75t_R g853 ( .A(n_651), .Y(n_853) );
NOR2xp67_ASAP7_75t_SL g854 ( .A(n_767), .B(n_78), .Y(n_854) );
O2A1O1Ixp33_ASAP7_75t_SL g855 ( .A1(n_774), .A2(n_185), .B(n_271), .C(n_270), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_760), .A2(n_180), .B(n_268), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_739), .A2(n_179), .B(n_267), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_724), .B(n_78), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_733), .B(n_79), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_748), .A2(n_182), .B(n_265), .Y(n_860) );
NAND2xp5_ASAP7_75t_SL g861 ( .A(n_712), .B(n_80), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_719), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_862) );
A2O1A1Ixp33_ASAP7_75t_L g863 ( .A1(n_708), .A2(n_81), .B(n_82), .C(n_84), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_694), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_741), .A2(n_194), .B(n_259), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_659), .Y(n_866) );
O2A1O1Ixp33_ASAP7_75t_SL g867 ( .A1(n_701), .A2(n_175), .B(n_257), .C(n_256), .Y(n_867) );
INVx4_ASAP7_75t_L g868 ( .A(n_651), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_700), .Y(n_869) );
AOI31xp67_ASAP7_75t_L g870 ( .A1(n_711), .A2(n_160), .A3(n_254), .B(n_253), .Y(n_870) );
OAI21x1_ASAP7_75t_L g871 ( .A1(n_745), .A2(n_159), .B(n_249), .Y(n_871) );
O2A1O1Ixp33_ASAP7_75t_SL g872 ( .A1(n_747), .A2(n_157), .B(n_242), .C(n_241), .Y(n_872) );
BUFx6f_ASAP7_75t_L g873 ( .A(n_679), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_735), .Y(n_874) );
CKINVDCx11_ASAP7_75t_R g875 ( .A(n_661), .Y(n_875) );
BUFx6f_ASAP7_75t_L g876 ( .A(n_679), .Y(n_876) );
O2A1O1Ixp33_ASAP7_75t_SL g877 ( .A1(n_688), .A2(n_152), .B(n_239), .C(n_238), .Y(n_877) );
A2O1A1Ixp33_ASAP7_75t_L g878 ( .A1(n_714), .A2(n_81), .B(n_85), .C(n_87), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g879 ( .A(n_772), .Y(n_879) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_714), .A2(n_85), .B(n_87), .C(n_88), .Y(n_880) );
NAND3x1_ASAP7_75t_L g881 ( .A(n_751), .B(n_88), .C(n_89), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_641), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_638), .A2(n_156), .B(n_237), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_704), .Y(n_884) );
A2O1A1Ixp33_ASAP7_75t_L g885 ( .A1(n_723), .A2(n_89), .B(n_90), .C(n_91), .Y(n_885) );
A2O1A1Ixp33_ASAP7_75t_L g886 ( .A1(n_709), .A2(n_90), .B(n_91), .C(n_116), .Y(n_886) );
OAI21x1_ASAP7_75t_L g887 ( .A1(n_771), .A2(n_117), .B(n_119), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_693), .A2(n_120), .B(n_122), .Y(n_888) );
O2A1O1Ixp33_ASAP7_75t_L g889 ( .A1(n_710), .A2(n_125), .B(n_126), .C(n_127), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_715), .A2(n_128), .B(n_129), .Y(n_890) );
BUFx2_ASAP7_75t_L g891 ( .A(n_765), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_763), .Y(n_892) );
O2A1O1Ixp33_ASAP7_75t_SL g893 ( .A1(n_674), .A2(n_130), .B(n_133), .C(n_134), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_763), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_664), .B(n_135), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_729), .A2(n_137), .B1(n_143), .B2(n_144), .Y(n_896) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_697), .B(n_145), .C(n_146), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_718), .A2(n_147), .B(n_148), .Y(n_898) );
O2A1O1Ixp33_ASAP7_75t_L g899 ( .A1(n_736), .A2(n_149), .B(n_196), .C(n_198), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_763), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_725), .A2(n_199), .B(n_200), .Y(n_901) );
OAI21xp5_ASAP7_75t_L g902 ( .A1(n_773), .A2(n_203), .B(n_207), .Y(n_902) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_727), .A2(n_211), .B(n_212), .Y(n_903) );
BUFx3_ASAP7_75t_L g904 ( .A(n_754), .Y(n_904) );
AO31x2_ASAP7_75t_L g905 ( .A1(n_752), .A2(n_214), .A3(n_216), .B(n_219), .Y(n_905) );
AO31x2_ASAP7_75t_L g906 ( .A1(n_761), .A2(n_220), .A3(n_221), .B(n_222), .Y(n_906) );
AO31x2_ASAP7_75t_L g907 ( .A1(n_738), .A2(n_223), .A3(n_225), .B(n_227), .Y(n_907) );
O2A1O1Ixp33_ASAP7_75t_L g908 ( .A1(n_744), .A2(n_228), .B(n_230), .C(n_233), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_729), .B(n_234), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_758), .B(n_290), .Y(n_910) );
A2O1A1Ixp33_ASAP7_75t_L g911 ( .A1(n_744), .A2(n_757), .B(n_749), .C(n_755), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_716), .B(n_764), .Y(n_912) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_679), .Y(n_913) );
OAI21xp5_ASAP7_75t_L g914 ( .A1(n_683), .A2(n_737), .B(n_652), .Y(n_914) );
AO32x2_ASAP7_75t_L g915 ( .A1(n_648), .A2(n_691), .A3(n_696), .B1(n_740), .B2(n_762), .Y(n_915) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_750), .B(n_762), .C(n_759), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g917 ( .A1(n_750), .A2(n_775), .B1(n_769), .B2(n_762), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_759), .Y(n_918) );
AND2x2_ASAP7_75t_SL g919 ( .A(n_683), .B(n_652), .Y(n_919) );
OAI21x1_ASAP7_75t_L g920 ( .A1(n_775), .A2(n_678), .B(n_776), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_759), .A2(n_640), .B(n_684), .Y(n_921) );
O2A1O1Ixp33_ASAP7_75t_L g922 ( .A1(n_695), .A2(n_677), .B(n_663), .C(n_726), .Y(n_922) );
AND2x4_ASAP7_75t_L g923 ( .A(n_651), .B(n_639), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_639), .Y(n_924) );
NOR2xp33_ASAP7_75t_SL g925 ( .A(n_721), .B(n_680), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g926 ( .A1(n_640), .A2(n_684), .B(n_654), .Y(n_926) );
AO31x2_ASAP7_75t_L g927 ( .A1(n_644), .A2(n_678), .A3(n_677), .B(n_650), .Y(n_927) );
NAND2xp5_ASAP7_75t_SL g928 ( .A(n_660), .B(n_589), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_866), .Y(n_929) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_793), .A2(n_926), .B(n_921), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_928), .A2(n_830), .B1(n_791), .B2(n_820), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_862), .A2(n_828), .B1(n_830), .B2(n_807), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_786), .B(n_924), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g934 ( .A1(n_828), .A2(n_824), .B1(n_804), .B2(n_882), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_788), .A2(n_891), .B1(n_853), .B2(n_779), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_796), .A2(n_923), .B1(n_858), .B2(n_839), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_904), .B(n_859), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_794), .Y(n_938) );
A2O1A1Ixp33_ASAP7_75t_L g939 ( .A1(n_922), .A2(n_825), .B(n_821), .C(n_788), .Y(n_939) );
AOI222xp33_ASAP7_75t_L g940 ( .A1(n_879), .A2(n_925), .B1(n_852), .B2(n_785), .C1(n_809), .C2(n_848), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_811), .A2(n_909), .B1(n_833), .B2(n_829), .Y(n_941) );
OAI22xp33_ASAP7_75t_L g942 ( .A1(n_795), .A2(n_781), .B1(n_868), .B2(n_778), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_808), .B(n_814), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_834), .Y(n_944) );
BUFx2_ASAP7_75t_L g945 ( .A(n_827), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_849), .B(n_864), .Y(n_946) );
AO31x2_ASAP7_75t_L g947 ( .A1(n_892), .A2(n_894), .A3(n_900), .B(n_806), .Y(n_947) );
BUFx2_ASAP7_75t_L g948 ( .A(n_797), .Y(n_948) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_875), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_874), .B(n_923), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_784), .Y(n_951) );
A2O1A1Ixp33_ASAP7_75t_L g952 ( .A1(n_841), .A2(n_812), .B(n_895), .C(n_845), .Y(n_952) );
OR2x2_ASAP7_75t_L g953 ( .A(n_797), .B(n_799), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_868), .A2(n_919), .B1(n_831), .B2(n_823), .Y(n_954) );
OAI21xp5_ASAP7_75t_L g955 ( .A1(n_780), .A2(n_777), .B(n_782), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_789), .A2(n_787), .B(n_920), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_840), .Y(n_957) );
AO21x1_ASAP7_75t_L g958 ( .A1(n_896), .A2(n_889), .B(n_902), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_844), .B(n_869), .Y(n_959) );
A2O1A1Ixp33_ASAP7_75t_L g960 ( .A1(n_837), .A2(n_813), .B(n_815), .C(n_850), .Y(n_960) );
OAI211xp5_ASAP7_75t_SL g961 ( .A1(n_851), .A2(n_885), .B(n_838), .C(n_863), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_861), .A2(n_801), .B1(n_914), .B2(n_792), .Y(n_962) );
OR2x2_ASAP7_75t_L g963 ( .A(n_810), .B(n_835), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_896), .A2(n_881), .B1(n_910), .B2(n_880), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_840), .Y(n_965) );
BUFx2_ASAP7_75t_L g966 ( .A(n_915), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_817), .B(n_840), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_817), .B(n_878), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_912), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_847), .Y(n_970) );
BUFx8_ASAP7_75t_L g971 ( .A(n_915), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_826), .B(n_846), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g973 ( .A1(n_819), .A2(n_800), .B1(n_836), .B2(n_802), .Y(n_973) );
OA21x2_ASAP7_75t_L g974 ( .A1(n_798), .A2(n_832), .B(n_856), .Y(n_974) );
A2O1A1Ixp33_ASAP7_75t_L g975 ( .A1(n_843), .A2(n_886), .B(n_899), .C(n_908), .Y(n_975) );
INVx2_ASAP7_75t_SL g976 ( .A(n_918), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_884), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_927), .B(n_854), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_790), .A2(n_911), .B(n_805), .Y(n_979) );
AOI21xp33_ASAP7_75t_L g980 ( .A1(n_917), .A2(n_836), .B(n_916), .Y(n_980) );
A2O1A1Ixp33_ASAP7_75t_L g981 ( .A1(n_865), .A2(n_857), .B(n_860), .C(n_890), .Y(n_981) );
OAI21xp5_ASAP7_75t_L g982 ( .A1(n_887), .A2(n_883), .B(n_818), .Y(n_982) );
AND2x4_ASAP7_75t_L g983 ( .A(n_803), .B(n_876), .Y(n_983) );
AO31x2_ASAP7_75t_L g984 ( .A1(n_783), .A2(n_816), .A3(n_888), .B(n_901), .Y(n_984) );
OAI221xp5_ASAP7_75t_SL g985 ( .A1(n_898), .A2(n_903), .B1(n_897), .B2(n_906), .C(n_905), .Y(n_985) );
OR2x6_ASAP7_75t_L g986 ( .A(n_803), .B(n_822), .Y(n_986) );
NAND3x1_ASAP7_75t_L g987 ( .A(n_915), .B(n_906), .C(n_907), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_822), .B(n_842), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_906), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_855), .A2(n_867), .B(n_877), .Y(n_990) );
OAI22xp33_ASAP7_75t_L g991 ( .A1(n_822), .A2(n_842), .B1(n_876), .B2(n_873), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_842), .A2(n_873), .B1(n_913), .B2(n_871), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_913), .A2(n_870), .B1(n_893), .B2(n_907), .Y(n_993) );
AOI21xp5_ASAP7_75t_L g994 ( .A1(n_872), .A2(n_913), .B(n_907), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_928), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_866), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_791), .B(n_577), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_866), .Y(n_998) );
AOI21xp5_ASAP7_75t_L g999 ( .A1(n_793), .A2(n_926), .B(n_921), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_866), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_791), .B(n_577), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_928), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_866), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_904), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_866), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_791), .B(n_577), .Y(n_1006) );
NOR2x1_ASAP7_75t_R g1007 ( .A(n_778), .B(n_785), .Y(n_1007) );
A2O1A1Ixp33_ASAP7_75t_L g1008 ( .A1(n_922), .A2(n_793), .B(n_825), .C(n_821), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_820), .B(n_563), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_866), .Y(n_1010) );
AO31x2_ASAP7_75t_L g1011 ( .A1(n_892), .A2(n_644), .A3(n_900), .B(n_894), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_866), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_793), .A2(n_660), .B1(n_862), .B2(n_663), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_866), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_809), .B(n_581), .Y(n_1015) );
OA21x2_ASAP7_75t_L g1016 ( .A1(n_787), .A2(n_780), .B(n_920), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_866), .Y(n_1017) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_904), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_928), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_866), .Y(n_1020) );
INVx2_ASAP7_75t_L g1021 ( .A(n_924), .Y(n_1021) );
INVx2_ASAP7_75t_L g1022 ( .A(n_924), .Y(n_1022) );
INVx4_ASAP7_75t_L g1023 ( .A(n_778), .Y(n_1023) );
AO21x2_ASAP7_75t_L g1024 ( .A1(n_788), .A2(n_787), .B(n_921), .Y(n_1024) );
OA21x2_ASAP7_75t_L g1025 ( .A1(n_787), .A2(n_780), .B(n_920), .Y(n_1025) );
AOI21xp5_ASAP7_75t_L g1026 ( .A1(n_793), .A2(n_926), .B(n_921), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_866), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_809), .B(n_581), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_866), .Y(n_1029) );
AOI21xp5_ASAP7_75t_L g1030 ( .A1(n_793), .A2(n_926), .B(n_921), .Y(n_1030) );
OA21x2_ASAP7_75t_L g1031 ( .A1(n_787), .A2(n_780), .B(n_920), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_866), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_866), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_928), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_809), .B(n_581), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g1036 ( .A(n_778), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_828), .A2(n_724), .B1(n_746), .B2(n_925), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_928), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_866), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_928), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_791), .B(n_577), .Y(n_1041) );
INVx3_ASAP7_75t_L g1042 ( .A(n_835), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_791), .B(n_577), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_928), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_1044) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_828), .A2(n_724), .B1(n_746), .B2(n_925), .Y(n_1045) );
A2O1A1Ixp33_ASAP7_75t_L g1046 ( .A1(n_922), .A2(n_793), .B(n_825), .C(n_821), .Y(n_1046) );
AOI21xp5_ASAP7_75t_L g1047 ( .A1(n_793), .A2(n_926), .B(n_921), .Y(n_1047) );
OAI21xp33_ASAP7_75t_L g1048 ( .A1(n_793), .A2(n_788), .B(n_719), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_866), .Y(n_1049) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_793), .A2(n_724), .B1(n_746), .B2(n_663), .Y(n_1050) );
AND2x4_ASAP7_75t_L g1051 ( .A(n_793), .B(n_923), .Y(n_1051) );
OAI211xp5_ASAP7_75t_L g1052 ( .A1(n_848), .A2(n_824), .B(n_513), .C(n_675), .Y(n_1052) );
OAI21x1_ASAP7_75t_L g1053 ( .A1(n_920), .A2(n_798), .B(n_787), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_820), .B(n_563), .Y(n_1054) );
OAI21x1_ASAP7_75t_L g1055 ( .A1(n_920), .A2(n_798), .B(n_787), .Y(n_1055) );
OAI221xp5_ASAP7_75t_L g1056 ( .A1(n_791), .A2(n_746), .B1(n_671), .B2(n_724), .C(n_549), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_938), .Y(n_1057) );
OAI21xp5_ASAP7_75t_L g1058 ( .A1(n_1008), .A2(n_1046), .B(n_952), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_944), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1004), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1011), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_933), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_1037), .A2(n_1045), .B1(n_995), .B2(n_1002), .Y(n_1063) );
INVx2_ASAP7_75t_SL g1064 ( .A(n_1051), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1009), .B(n_1054), .Y(n_1065) );
OR2x6_ASAP7_75t_L g1066 ( .A(n_1013), .B(n_935), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_931), .B(n_1013), .Y(n_1067) );
AOI211xp5_ASAP7_75t_SL g1068 ( .A1(n_935), .A2(n_1056), .B(n_1050), .C(n_1052), .Y(n_1068) );
INVx2_ASAP7_75t_SL g1069 ( .A(n_1018), .Y(n_1069) );
AO21x2_ASAP7_75t_L g1070 ( .A1(n_989), .A2(n_979), .B(n_978), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1071 ( .A(n_945), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_997), .B(n_1001), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1021), .B(n_1022), .Y(n_1073) );
AO21x2_ASAP7_75t_L g1074 ( .A1(n_930), .A2(n_1047), .B(n_1030), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_929), .Y(n_1075) );
OR2x6_ASAP7_75t_L g1076 ( .A(n_1048), .B(n_986), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_996), .Y(n_1077) );
BUFx3_ASAP7_75t_L g1078 ( .A(n_948), .Y(n_1078) );
INVx4_ASAP7_75t_L g1079 ( .A(n_986), .Y(n_1079) );
OR2x2_ASAP7_75t_L g1080 ( .A(n_1015), .B(n_1028), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_998), .Y(n_1081) );
INVxp67_ASAP7_75t_L g1082 ( .A(n_1007), .Y(n_1082) );
OA21x2_ASAP7_75t_L g1083 ( .A1(n_956), .A2(n_1055), .B(n_1053), .Y(n_1083) );
OA332x1_ASAP7_75t_L g1084 ( .A1(n_1019), .A2(n_1034), .A3(n_1038), .B1(n_1040), .B2(n_1044), .B3(n_964), .C1(n_940), .C2(n_1050), .Y(n_1084) );
AO21x2_ASAP7_75t_L g1085 ( .A1(n_999), .A2(n_1026), .B(n_965), .Y(n_1085) );
NOR2x1_ASAP7_75t_L g1086 ( .A(n_970), .B(n_942), .Y(n_1086) );
AO21x2_ASAP7_75t_L g1087 ( .A1(n_957), .A2(n_994), .B(n_955), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_932), .A2(n_941), .B1(n_934), .B2(n_936), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_947), .Y(n_1089) );
OR2x6_ASAP7_75t_L g1090 ( .A(n_1048), .B(n_986), .Y(n_1090) );
AO21x2_ASAP7_75t_L g1091 ( .A1(n_955), .A2(n_980), .B(n_990), .Y(n_1091) );
AND2x4_ASAP7_75t_SL g1092 ( .A(n_1023), .B(n_1036), .Y(n_1092) );
OR2x6_ASAP7_75t_L g1093 ( .A(n_966), .B(n_964), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1000), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1003), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1005), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_953), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_969), .B(n_932), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_950), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_1006), .A2(n_1041), .B1(n_1043), .B2(n_1049), .C(n_1039), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1016), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1010), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1012), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1014), .B(n_1029), .Y(n_1104) );
OAI21xp5_ASAP7_75t_L g1105 ( .A1(n_939), .A2(n_960), .B(n_941), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1017), .Y(n_1106) );
OAI21xp5_ASAP7_75t_L g1107 ( .A1(n_934), .A2(n_961), .B(n_951), .Y(n_1107) );
AOI221xp5_ASAP7_75t_L g1108 ( .A1(n_1020), .A2(n_1032), .B1(n_1027), .B2(n_1033), .C(n_959), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_943), .Y(n_1109) );
OAI21xp5_ASAP7_75t_L g1110 ( .A1(n_975), .A2(n_954), .B(n_962), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_946), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_977), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_937), .B(n_940), .Y(n_1113) );
OA21x2_ASAP7_75t_L g1114 ( .A1(n_993), .A2(n_967), .B(n_982), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_963), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_972), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1042), .Y(n_1117) );
AO21x2_ASAP7_75t_L g1118 ( .A1(n_1024), .A2(n_982), .B(n_968), .Y(n_1118) );
OAI33xp33_ASAP7_75t_L g1119 ( .A1(n_1035), .A2(n_991), .A3(n_988), .B1(n_987), .B2(n_985), .B3(n_973), .Y(n_1119) );
INVx3_ASAP7_75t_L g1120 ( .A(n_971), .Y(n_1120) );
OA21x2_ASAP7_75t_L g1121 ( .A1(n_992), .A2(n_981), .B(n_958), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_976), .B(n_1031), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_971), .Y(n_1123) );
NAND4xp25_ASAP7_75t_L g1124 ( .A(n_1023), .B(n_949), .C(n_984), .D(n_1025), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1031), .B(n_974), .Y(n_1125) );
INVx8_ASAP7_75t_L g1126 ( .A(n_984), .Y(n_1126) );
INVx3_ASAP7_75t_SL g1127 ( .A(n_1036), .Y(n_1127) );
OAI21xp5_ASAP7_75t_L g1128 ( .A1(n_1008), .A2(n_1046), .B(n_952), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_1051), .B(n_983), .Y(n_1129) );
OAI21xp5_ASAP7_75t_L g1130 ( .A1(n_1008), .A2(n_1046), .B(n_952), .Y(n_1130) );
BUFx2_ASAP7_75t_L g1131 ( .A(n_1018), .Y(n_1131) );
INVxp67_ASAP7_75t_SL g1132 ( .A(n_1051), .Y(n_1132) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1004), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1009), .B(n_1054), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1018), .B(n_1004), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_1004), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1066), .B(n_1067), .Y(n_1137) );
INVxp67_ASAP7_75t_SL g1138 ( .A(n_1132), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1101), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1061), .Y(n_1140) );
INVx1_ASAP7_75t_SL g1141 ( .A(n_1071), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_1060), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1066), .B(n_1067), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_1063), .A2(n_1088), .B1(n_1107), .B2(n_1105), .C(n_1068), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1061), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1066), .B(n_1098), .Y(n_1146) );
BUFx2_ASAP7_75t_L g1147 ( .A(n_1076), .Y(n_1147) );
HB1xp67_ASAP7_75t_L g1148 ( .A(n_1133), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1098), .B(n_1073), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1058), .B(n_1128), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1123), .B(n_1080), .Y(n_1151) );
INVxp67_ASAP7_75t_SL g1152 ( .A(n_1099), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1130), .B(n_1100), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1113), .B(n_1124), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1073), .B(n_1116), .Y(n_1155) );
A2O1A1Ixp33_ASAP7_75t_L g1156 ( .A1(n_1063), .A2(n_1110), .B(n_1086), .C(n_1078), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1109), .B(n_1111), .Y(n_1157) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_1120), .B(n_1122), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1057), .B(n_1059), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1065), .B(n_1134), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1118), .B(n_1075), .Y(n_1161) );
INVx1_ASAP7_75t_SL g1162 ( .A(n_1071), .Y(n_1162) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_1136), .Y(n_1163) );
BUFx2_ASAP7_75t_L g1164 ( .A(n_1076), .Y(n_1164) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_1076), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1118), .B(n_1103), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1118), .B(n_1102), .Y(n_1167) );
BUFx2_ASAP7_75t_L g1168 ( .A(n_1076), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1169 ( .A(n_1078), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1077), .B(n_1096), .Y(n_1170) );
OR2x6_ASAP7_75t_L g1171 ( .A(n_1090), .B(n_1093), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1115), .Y(n_1172) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_1097), .Y(n_1173) );
INVx4_ASAP7_75t_L g1174 ( .A(n_1079), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1081), .B(n_1106), .Y(n_1175) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1108), .B(n_1095), .Y(n_1176) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_1120), .B(n_1090), .Y(n_1177) );
AND2x4_ASAP7_75t_L g1178 ( .A(n_1090), .B(n_1089), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1097), .B(n_1093), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_1064), .A2(n_1093), .B1(n_1090), .B2(n_1062), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1094), .B(n_1112), .Y(n_1181) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_1072), .A2(n_1084), .B1(n_1064), .B2(n_1082), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1104), .B(n_1093), .Y(n_1183) );
AOI21xp5_ASAP7_75t_L g1184 ( .A1(n_1126), .A2(n_1074), .B(n_1083), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1161), .B(n_1114), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1166), .B(n_1114), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1166), .Y(n_1187) );
INVx2_ASAP7_75t_L g1188 ( .A(n_1139), .Y(n_1188) );
INVx1_ASAP7_75t_SL g1189 ( .A(n_1141), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1167), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1183), .B(n_1114), .Y(n_1191) );
BUFx2_ASAP7_75t_L g1192 ( .A(n_1169), .Y(n_1192) );
INVx3_ASAP7_75t_L g1193 ( .A(n_1178), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1167), .B(n_1085), .Y(n_1194) );
INVx1_ASAP7_75t_SL g1195 ( .A(n_1141), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_1144), .A2(n_1119), .B1(n_1084), .B2(n_1131), .Y(n_1196) );
NOR2x1_ASAP7_75t_L g1197 ( .A(n_1174), .B(n_1079), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1183), .B(n_1069), .Y(n_1198) );
AND2x4_ASAP7_75t_SL g1199 ( .A(n_1174), .B(n_1079), .Y(n_1199) );
NAND2xp5_ASAP7_75t_SL g1200 ( .A(n_1162), .B(n_1069), .Y(n_1200) );
AND2x4_ASAP7_75t_L g1201 ( .A(n_1177), .B(n_1087), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1146), .B(n_1085), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1149), .B(n_1146), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1149), .B(n_1070), .Y(n_1204) );
AND2x4_ASAP7_75t_SL g1205 ( .A(n_1174), .B(n_1129), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1153), .B(n_1126), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1140), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1153), .B(n_1126), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1137), .B(n_1135), .Y(n_1209) );
INVx1_ASAP7_75t_SL g1210 ( .A(n_1162), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1176), .B(n_1070), .Y(n_1211) );
BUFx2_ASAP7_75t_L g1212 ( .A(n_1177), .Y(n_1212) );
HB1xp67_ASAP7_75t_L g1213 ( .A(n_1173), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1214 ( .A(n_1142), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1140), .Y(n_1215) );
HB1xp67_ASAP7_75t_L g1216 ( .A(n_1148), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1143), .B(n_1125), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1145), .Y(n_1218) );
HB1xp67_ASAP7_75t_L g1219 ( .A(n_1163), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1176), .B(n_1121), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1150), .B(n_1121), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1158), .B(n_1091), .Y(n_1222) );
INVx1_ASAP7_75t_SL g1223 ( .A(n_1172), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1158), .B(n_1121), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1204), .B(n_1171), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1207), .Y(n_1226) );
INVx2_ASAP7_75t_SL g1227 ( .A(n_1192), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1215), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1204), .B(n_1171), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1214), .B(n_1152), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1214), .B(n_1170), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1204), .B(n_1171), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1202), .B(n_1171), .Y(n_1233) );
AOI22xp5_ASAP7_75t_L g1234 ( .A1(n_1196), .A2(n_1144), .B1(n_1182), .B2(n_1150), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1235 ( .A(n_1192), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1202), .B(n_1171), .Y(n_1236) );
NAND2xp33_ASAP7_75t_SL g1237 ( .A(n_1216), .B(n_1127), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1202), .B(n_1177), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1187), .B(n_1154), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1185), .B(n_1178), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1216), .B(n_1170), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1215), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1218), .Y(n_1243) );
NAND3xp33_ASAP7_75t_L g1244 ( .A(n_1219), .B(n_1156), .C(n_1182), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1187), .B(n_1154), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1190), .B(n_1179), .Y(n_1246) );
AND2x2_ASAP7_75t_SL g1247 ( .A(n_1205), .B(n_1147), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1190), .B(n_1151), .Y(n_1248) );
NOR2x1_ASAP7_75t_L g1249 ( .A(n_1197), .B(n_1174), .Y(n_1249) );
AND2x4_ASAP7_75t_L g1250 ( .A(n_1201), .B(n_1178), .Y(n_1250) );
INVx1_ASAP7_75t_SL g1251 ( .A(n_1223), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1217), .B(n_1151), .Y(n_1252) );
AOI21xp5_ASAP7_75t_L g1253 ( .A1(n_1197), .A2(n_1184), .B(n_1180), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1185), .B(n_1178), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_1213), .Y(n_1255) );
INVx3_ASAP7_75t_L g1256 ( .A(n_1201), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1219), .B(n_1175), .Y(n_1257) );
NOR2xp33_ASAP7_75t_L g1258 ( .A(n_1223), .B(n_1127), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_1213), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1185), .B(n_1164), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1203), .B(n_1175), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1217), .B(n_1180), .Y(n_1262) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1188), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1186), .B(n_1147), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1240), .B(n_1222), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1226), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1239), .B(n_1203), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1226), .Y(n_1268) );
INVx1_ASAP7_75t_SL g1269 ( .A(n_1251), .Y(n_1269) );
NOR3xp33_ASAP7_75t_L g1270 ( .A(n_1244), .B(n_1200), .C(n_1220), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1245), .B(n_1191), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1240), .B(n_1222), .Y(n_1272) );
INVxp67_ASAP7_75t_L g1273 ( .A(n_1258), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1245), .B(n_1194), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1255), .B(n_1194), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1259), .B(n_1220), .Y(n_1276) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_1244), .A2(n_1160), .B1(n_1206), .B2(n_1208), .C(n_1211), .Y(n_1277) );
INVx2_ASAP7_75t_L g1278 ( .A(n_1263), .Y(n_1278) );
INVx1_ASAP7_75t_SL g1279 ( .A(n_1237), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1231), .B(n_1206), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1254), .B(n_1222), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1254), .B(n_1224), .Y(n_1282) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1263), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1228), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1252), .B(n_1191), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1228), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1260), .B(n_1224), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1242), .Y(n_1288) );
INVxp67_ASAP7_75t_L g1289 ( .A(n_1235), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1242), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1243), .Y(n_1291) );
INVx1_ASAP7_75t_SL g1292 ( .A(n_1252), .Y(n_1292) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_1273), .B(n_1230), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1265), .B(n_1256), .Y(n_1294) );
INVx3_ASAP7_75t_L g1295 ( .A(n_1278), .Y(n_1295) );
NAND3xp33_ASAP7_75t_L g1296 ( .A(n_1277), .B(n_1234), .C(n_1227), .Y(n_1296) );
INVx1_ASAP7_75t_SL g1297 ( .A(n_1269), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1270), .B(n_1227), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1266), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1265), .B(n_1256), .Y(n_1300) );
INVxp67_ASAP7_75t_L g1301 ( .A(n_1279), .Y(n_1301) );
OAI21xp5_ASAP7_75t_L g1302 ( .A1(n_1289), .A2(n_1249), .B(n_1234), .Y(n_1302) );
NAND2xp5_ASAP7_75t_SL g1303 ( .A(n_1292), .B(n_1247), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1266), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1285), .B(n_1241), .Y(n_1305) );
OAI211xp5_ASAP7_75t_L g1306 ( .A1(n_1276), .A2(n_1249), .B(n_1253), .C(n_1257), .Y(n_1306) );
AOI21xp5_ASAP7_75t_L g1307 ( .A1(n_1275), .A2(n_1247), .B(n_1205), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1268), .Y(n_1308) );
OAI322xp33_ASAP7_75t_L g1309 ( .A1(n_1285), .A2(n_1248), .A3(n_1262), .B1(n_1261), .B2(n_1246), .C1(n_1209), .C2(n_1208), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1272), .B(n_1256), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1274), .B(n_1264), .Y(n_1311) );
INVxp67_ASAP7_75t_SL g1312 ( .A(n_1278), .Y(n_1312) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1283), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1299), .Y(n_1314) );
O2A1O1Ixp5_ASAP7_75t_L g1315 ( .A1(n_1302), .A2(n_1280), .B(n_1256), .C(n_1267), .Y(n_1315) );
AO21x1_ASAP7_75t_L g1316 ( .A1(n_1298), .A2(n_1199), .B(n_1092), .Y(n_1316) );
OAI221xp5_ASAP7_75t_SL g1317 ( .A1(n_1301), .A2(n_1262), .B1(n_1271), .B2(n_1209), .C(n_1233), .Y(n_1317) );
INVxp67_ASAP7_75t_L g1318 ( .A(n_1297), .Y(n_1318) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1295), .Y(n_1319) );
OAI32xp33_ASAP7_75t_L g1320 ( .A1(n_1297), .A2(n_1296), .A3(n_1303), .B1(n_1293), .B2(n_1305), .Y(n_1320) );
AOI322xp5_ASAP7_75t_L g1321 ( .A1(n_1294), .A2(n_1287), .A3(n_1282), .B1(n_1281), .B2(n_1264), .C1(n_1232), .C2(n_1229), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1305), .Y(n_1322) );
INVxp67_ASAP7_75t_L g1323 ( .A(n_1312), .Y(n_1323) );
OAI221xp5_ASAP7_75t_SL g1324 ( .A1(n_1306), .A2(n_1233), .B1(n_1236), .B2(n_1225), .C(n_1229), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1299), .Y(n_1325) );
INVx1_ASAP7_75t_SL g1326 ( .A(n_1307), .Y(n_1326) );
OAI211xp5_ASAP7_75t_L g1327 ( .A1(n_1320), .A2(n_1195), .B(n_1189), .C(n_1210), .Y(n_1327) );
AOI221xp5_ASAP7_75t_L g1328 ( .A1(n_1320), .A2(n_1309), .B1(n_1308), .B2(n_1304), .C(n_1295), .Y(n_1328) );
AOI21xp5_ASAP7_75t_L g1329 ( .A1(n_1316), .A2(n_1247), .B(n_1092), .Y(n_1329) );
AOI222xp33_ASAP7_75t_L g1330 ( .A1(n_1326), .A2(n_1310), .B1(n_1300), .B2(n_1294), .C1(n_1295), .C2(n_1311), .Y(n_1330) );
OAI221xp5_ASAP7_75t_L g1331 ( .A1(n_1315), .A2(n_1310), .B1(n_1300), .B2(n_1313), .C(n_1195), .Y(n_1331) );
AOI221x1_ASAP7_75t_L g1332 ( .A1(n_1322), .A2(n_1313), .B1(n_1291), .B2(n_1284), .C(n_1290), .Y(n_1332) );
AOI221xp5_ASAP7_75t_L g1333 ( .A1(n_1317), .A2(n_1288), .B1(n_1286), .B2(n_1284), .C(n_1268), .Y(n_1333) );
AOI22xp5_ASAP7_75t_L g1334 ( .A1(n_1316), .A2(n_1236), .B1(n_1232), .B2(n_1225), .Y(n_1334) );
NOR2x1_ASAP7_75t_L g1335 ( .A(n_1327), .B(n_1319), .Y(n_1335) );
NOR5xp2_ASAP7_75t_L g1336 ( .A(n_1331), .B(n_1318), .C(n_1324), .D(n_1323), .E(n_1314), .Y(n_1336) );
OAI221xp5_ASAP7_75t_L g1337 ( .A1(n_1328), .A2(n_1321), .B1(n_1319), .B2(n_1314), .C(n_1325), .Y(n_1337) );
NAND2xp5_ASAP7_75t_SL g1338 ( .A(n_1329), .B(n_1189), .Y(n_1338) );
NOR3xp33_ASAP7_75t_L g1339 ( .A(n_1333), .B(n_1157), .C(n_1211), .Y(n_1339) );
NOR3x1_ASAP7_75t_L g1340 ( .A(n_1337), .B(n_1330), .C(n_1212), .Y(n_1340) );
NAND5xp2_ASAP7_75t_L g1341 ( .A(n_1336), .B(n_1334), .C(n_1165), .D(n_1168), .E(n_1164), .Y(n_1341) );
NOR3xp33_ASAP7_75t_L g1342 ( .A(n_1338), .B(n_1157), .C(n_1221), .Y(n_1342) );
NOR3xp33_ASAP7_75t_L g1343 ( .A(n_1335), .B(n_1221), .C(n_1159), .Y(n_1343) );
NOR2x1_ASAP7_75t_L g1344 ( .A(n_1341), .B(n_1332), .Y(n_1344) );
NAND4xp75_ASAP7_75t_L g1345 ( .A(n_1340), .B(n_1339), .C(n_1238), .D(n_1181), .Y(n_1345) );
OAI22xp5_ASAP7_75t_SL g1346 ( .A1(n_1343), .A2(n_1138), .B1(n_1168), .B2(n_1165), .Y(n_1346) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1345), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_1344), .A2(n_1342), .B1(n_1198), .B2(n_1199), .Y(n_1348) );
HB1xp67_ASAP7_75t_L g1349 ( .A(n_1347), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1348), .Y(n_1350) );
AOI222xp33_ASAP7_75t_SL g1351 ( .A1(n_1349), .A2(n_1350), .B1(n_1346), .B2(n_1212), .C1(n_1193), .C2(n_1117), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1350), .Y(n_1352) );
XNOR2xp5_ASAP7_75t_L g1353 ( .A(n_1352), .B(n_1205), .Y(n_1353) );
XNOR2x1_ASAP7_75t_L g1354 ( .A(n_1353), .B(n_1351), .Y(n_1354) );
AOI22xp5_ASAP7_75t_L g1355 ( .A1(n_1354), .A2(n_1250), .B1(n_1155), .B2(n_1201), .Y(n_1355) );
endmodule