module fake_ariane_407_n_4585 (n_295, n_356, n_556, n_170, n_190, n_698, n_1072, n_695, n_913, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_1008, n_581, n_294, n_1020, n_646, n_197, n_640, n_463, n_1024, n_830, n_176, n_691, n_34, n_404, n_172, n_943, n_678, n_1058, n_651, n_987, n_936, n_347, n_423, n_1042, n_961, n_183, n_469, n_1046, n_479, n_726, n_603, n_878, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_850, n_908, n_771, n_1036, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_1029, n_985, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_906, n_416, n_969, n_283, n_919, n_50, n_187, n_525, n_806, n_367, n_970, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_924, n_927, n_781, n_220, n_261, n_1095, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_864, n_952, n_1096, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_940, n_346, n_1016, n_214, n_764, n_979, n_348, n_552, n_1077, n_2, n_462, n_607, n_670, n_897, n_32, n_949, n_956, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_891, n_737, n_137, n_885, n_122, n_198, n_232, n_52, n_441, n_568, n_1032, n_385, n_637, n_917, n_73, n_327, n_77, n_1088, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_960, n_520, n_980, n_870, n_87, n_714, n_279, n_905, n_702, n_945, n_958, n_207, n_790, n_857, n_898, n_363, n_720, n_968, n_1067, n_354, n_41, n_813, n_926, n_140, n_725, n_419, n_151, n_28, n_146, n_1009, n_230, n_270, n_194, n_1064, n_633, n_900, n_154, n_883, n_338, n_142, n_995, n_285, n_1093, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_871, n_315, n_903, n_1073, n_594, n_311, n_239, n_402, n_35, n_1052, n_1068, n_272, n_54, n_829, n_1062, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_879, n_167, n_90, n_38, n_422, n_1106, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_1018, n_855, n_158, n_1047, n_69, n_259, n_835, n_95, n_808, n_953, n_446, n_553, n_1076, n_143, n_753, n_1050, n_566, n_814, n_578, n_701, n_1003, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_1107, n_173, n_858, n_242, n_645, n_989, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_1035, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_1053, n_1084, n_398, n_62, n_210, n_1090, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_928, n_1099, n_3, n_271, n_465, n_486, n_507, n_901, n_759, n_247, n_569, n_567, n_825, n_732, n_1103, n_91, n_971, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_894, n_31, n_1105, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_1061, n_1045, n_831, n_256, n_868, n_326, n_681, n_778, n_227, n_48, n_874, n_188, n_323, n_550, n_1023, n_988, n_635, n_707, n_997, n_330, n_914, n_400, n_689, n_694, n_884, n_11, n_129, n_126, n_983, n_282, n_328, n_368, n_1034, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_1085, n_432, n_545, n_1015, n_536, n_644, n_293, n_823, n_921, n_620, n_228, n_325, n_276, n_93, n_688, n_1074, n_859, n_636, n_427, n_108, n_587, n_497, n_1098, n_693, n_863, n_303, n_671, n_442, n_777, n_929, n_168, n_81, n_1, n_206, n_352, n_538, n_899, n_920, n_576, n_843, n_1080, n_511, n_1086, n_611, n_1092, n_238, n_365, n_429, n_455, n_654, n_588, n_1013, n_986, n_1104, n_638, n_136, n_334, n_192, n_729, n_887, n_661, n_488, n_1048, n_775, n_667, n_1049, n_300, n_533, n_904, n_505, n_14, n_163, n_88, n_869, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_1059, n_314, n_684, n_16, n_440, n_627, n_1039, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_957, n_977, n_512, n_715, n_889, n_1066, n_935, n_579, n_844, n_1012, n_459, n_685, n_221, n_321, n_911, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_861, n_175, n_950, n_1017, n_711, n_877, n_1021, n_1065, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_1055, n_260, n_362, n_543, n_942, n_310, n_709, n_236, n_601, n_683, n_565, n_1089, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_907, n_235, n_1006, n_881, n_660, n_464, n_735, n_575, n_546, n_1019, n_297, n_962, n_662, n_641, n_1005, n_503, n_941, n_700, n_910, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_939, n_371, n_845, n_888, n_199, n_918, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_1038, n_70, n_572, n_343, n_865, n_10, n_1041, n_414, n_571, n_680, n_287, n_302, n_993, n_380, n_6, n_948, n_582, n_94, n_284, n_922, n_1004, n_4, n_448, n_593, n_755, n_1097, n_710, n_860, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_851, n_1043, n_255, n_560, n_450, n_890, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_1022, n_135, n_1033, n_896, n_409, n_171, n_947, n_930, n_519, n_902, n_384, n_1031, n_468, n_1056, n_853, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_1040, n_674, n_1081, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_872, n_933, n_13, n_27, n_916, n_254, n_596, n_954, n_912, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_982, n_915, n_215, n_252, n_629, n_664, n_161, n_1075, n_454, n_966, n_992, n_298, n_955, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_1091, n_514, n_418, n_984, n_537, n_1063, n_223, n_403, n_25, n_750, n_834, n_991, n_83, n_389, n_1007, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_951, n_1026, n_213, n_938, n_862, n_110, n_304, n_895, n_659, n_67, n_509, n_583, n_1014, n_724, n_306, n_666, n_1000, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_946, n_757, n_375, n_113, n_114, n_33, n_324, n_1030, n_1100, n_585, n_875, n_669, n_785, n_827, n_931, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_967, n_998, n_999, n_1083, n_472, n_937, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_880, n_793, n_852, n_1079, n_174, n_275, n_100, n_704, n_1060, n_132, n_1044, n_147, n_204, n_751, n_615, n_1027, n_1070, n_996, n_521, n_963, n_873, n_51, n_1082, n_496, n_739, n_1028, n_76, n_342, n_866, n_26, n_246, n_517, n_925, n_530, n_1094, n_0, n_792, n_1001, n_824, n_428, n_159, n_1002, n_358, n_105, n_580, n_892, n_608, n_959, n_30, n_494, n_1051, n_719, n_131, n_263, n_434, n_360, n_1101, n_975, n_1102, n_563, n_229, n_394, n_923, n_250, n_932, n_773, n_165, n_1037, n_144, n_981, n_1010, n_882, n_990, n_317, n_867, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_944, n_749, n_994, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_973, n_523, n_1078, n_268, n_972, n_266, n_470, n_457, n_1087, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_856, n_425, n_431, n_811, n_1054, n_508, n_624, n_118, n_121, n_791, n_876, n_618, n_1071, n_411, n_484, n_712, n_849, n_909, n_976, n_353, n_22, n_736, n_767, n_1025, n_241, n_29, n_357, n_412, n_687, n_447, n_964, n_1057, n_191, n_382, n_797, n_489, n_80, n_480, n_978, n_211, n_642, n_1011, n_97, n_408, n_828, n_595, n_322, n_251, n_974, n_506, n_893, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_854, n_471, n_351, n_886, n_965, n_39, n_393, n_1069, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_934, n_783, n_675, n_4585);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_1072;
input n_695;
input n_913;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_1008;
input n_581;
input n_294;
input n_1020;
input n_646;
input n_197;
input n_640;
input n_463;
input n_1024;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_943;
input n_678;
input n_1058;
input n_651;
input n_987;
input n_936;
input n_347;
input n_423;
input n_1042;
input n_961;
input n_183;
input n_469;
input n_1046;
input n_479;
input n_726;
input n_603;
input n_878;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_850;
input n_908;
input n_771;
input n_1036;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_1029;
input n_985;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_906;
input n_416;
input n_969;
input n_283;
input n_919;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_970;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_924;
input n_927;
input n_781;
input n_220;
input n_261;
input n_1095;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_864;
input n_952;
input n_1096;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_940;
input n_346;
input n_1016;
input n_214;
input n_764;
input n_979;
input n_348;
input n_552;
input n_1077;
input n_2;
input n_462;
input n_607;
input n_670;
input n_897;
input n_32;
input n_949;
input n_956;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_891;
input n_737;
input n_137;
input n_885;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_1032;
input n_385;
input n_637;
input n_917;
input n_73;
input n_327;
input n_77;
input n_1088;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_960;
input n_520;
input n_980;
input n_870;
input n_87;
input n_714;
input n_279;
input n_905;
input n_702;
input n_945;
input n_958;
input n_207;
input n_790;
input n_857;
input n_898;
input n_363;
input n_720;
input n_968;
input n_1067;
input n_354;
input n_41;
input n_813;
input n_926;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_1009;
input n_230;
input n_270;
input n_194;
input n_1064;
input n_633;
input n_900;
input n_154;
input n_883;
input n_338;
input n_142;
input n_995;
input n_285;
input n_1093;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_871;
input n_315;
input n_903;
input n_1073;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_1052;
input n_1068;
input n_272;
input n_54;
input n_829;
input n_1062;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_879;
input n_167;
input n_90;
input n_38;
input n_422;
input n_1106;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_1018;
input n_855;
input n_158;
input n_1047;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_953;
input n_446;
input n_553;
input n_1076;
input n_143;
input n_753;
input n_1050;
input n_566;
input n_814;
input n_578;
input n_701;
input n_1003;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_1107;
input n_173;
input n_858;
input n_242;
input n_645;
input n_989;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_1035;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_1053;
input n_1084;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_928;
input n_1099;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_901;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_1103;
input n_91;
input n_971;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_894;
input n_31;
input n_1105;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_1061;
input n_1045;
input n_831;
input n_256;
input n_868;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_874;
input n_188;
input n_323;
input n_550;
input n_1023;
input n_988;
input n_635;
input n_707;
input n_997;
input n_330;
input n_914;
input n_400;
input n_689;
input n_694;
input n_884;
input n_11;
input n_129;
input n_126;
input n_983;
input n_282;
input n_328;
input n_368;
input n_1034;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_1085;
input n_432;
input n_545;
input n_1015;
input n_536;
input n_644;
input n_293;
input n_823;
input n_921;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_1074;
input n_859;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_1098;
input n_693;
input n_863;
input n_303;
input n_671;
input n_442;
input n_777;
input n_929;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_899;
input n_920;
input n_576;
input n_843;
input n_1080;
input n_511;
input n_1086;
input n_611;
input n_1092;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_1013;
input n_986;
input n_1104;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_887;
input n_661;
input n_488;
input n_1048;
input n_775;
input n_667;
input n_1049;
input n_300;
input n_533;
input n_904;
input n_505;
input n_14;
input n_163;
input n_88;
input n_869;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_1059;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_1039;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_957;
input n_977;
input n_512;
input n_715;
input n_889;
input n_1066;
input n_935;
input n_579;
input n_844;
input n_1012;
input n_459;
input n_685;
input n_221;
input n_321;
input n_911;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_861;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_877;
input n_1021;
input n_1065;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_1055;
input n_260;
input n_362;
input n_543;
input n_942;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_1089;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_907;
input n_235;
input n_1006;
input n_881;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_1019;
input n_297;
input n_962;
input n_662;
input n_641;
input n_1005;
input n_503;
input n_941;
input n_700;
input n_910;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_939;
input n_371;
input n_845;
input n_888;
input n_199;
input n_918;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_1038;
input n_70;
input n_572;
input n_343;
input n_865;
input n_10;
input n_1041;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_993;
input n_380;
input n_6;
input n_948;
input n_582;
input n_94;
input n_284;
input n_922;
input n_1004;
input n_4;
input n_448;
input n_593;
input n_755;
input n_1097;
input n_710;
input n_860;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_851;
input n_1043;
input n_255;
input n_560;
input n_450;
input n_890;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_1022;
input n_135;
input n_1033;
input n_896;
input n_409;
input n_171;
input n_947;
input n_930;
input n_519;
input n_902;
input n_384;
input n_1031;
input n_468;
input n_1056;
input n_853;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_1040;
input n_674;
input n_1081;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_872;
input n_933;
input n_13;
input n_27;
input n_916;
input n_254;
input n_596;
input n_954;
input n_912;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_982;
input n_915;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_1075;
input n_454;
input n_966;
input n_992;
input n_298;
input n_955;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_1091;
input n_514;
input n_418;
input n_984;
input n_537;
input n_1063;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_991;
input n_83;
input n_389;
input n_1007;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_951;
input n_1026;
input n_213;
input n_938;
input n_862;
input n_110;
input n_304;
input n_895;
input n_659;
input n_67;
input n_509;
input n_583;
input n_1014;
input n_724;
input n_306;
input n_666;
input n_1000;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_1030;
input n_1100;
input n_585;
input n_875;
input n_669;
input n_785;
input n_827;
input n_931;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_967;
input n_998;
input n_999;
input n_1083;
input n_472;
input n_937;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_880;
input n_793;
input n_852;
input n_1079;
input n_174;
input n_275;
input n_100;
input n_704;
input n_1060;
input n_132;
input n_1044;
input n_147;
input n_204;
input n_751;
input n_615;
input n_1027;
input n_1070;
input n_996;
input n_521;
input n_963;
input n_873;
input n_51;
input n_1082;
input n_496;
input n_739;
input n_1028;
input n_76;
input n_342;
input n_866;
input n_26;
input n_246;
input n_517;
input n_925;
input n_530;
input n_1094;
input n_0;
input n_792;
input n_1001;
input n_824;
input n_428;
input n_159;
input n_1002;
input n_358;
input n_105;
input n_580;
input n_892;
input n_608;
input n_959;
input n_30;
input n_494;
input n_1051;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_1101;
input n_975;
input n_1102;
input n_563;
input n_229;
input n_394;
input n_923;
input n_250;
input n_932;
input n_773;
input n_165;
input n_1037;
input n_144;
input n_981;
input n_1010;
input n_882;
input n_990;
input n_317;
input n_867;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_944;
input n_749;
input n_994;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_973;
input n_523;
input n_1078;
input n_268;
input n_972;
input n_266;
input n_470;
input n_457;
input n_1087;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_856;
input n_425;
input n_431;
input n_811;
input n_1054;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_876;
input n_618;
input n_1071;
input n_411;
input n_484;
input n_712;
input n_849;
input n_909;
input n_976;
input n_353;
input n_22;
input n_736;
input n_767;
input n_1025;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_964;
input n_1057;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_978;
input n_211;
input n_642;
input n_1011;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_974;
input n_506;
input n_893;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_854;
input n_471;
input n_351;
input n_886;
input n_965;
input n_39;
input n_393;
input n_1069;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_934;
input n_783;
input n_675;

output n_4585;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_4030;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_4342;
wire n_4557;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_4382;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2680;
wire n_2334;
wire n_4259;
wire n_3264;
wire n_4475;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_3181;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_4403;
wire n_1713;
wire n_2818;
wire n_1436;
wire n_2407;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_1430;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_1837;
wire n_4178;
wire n_2013;
wire n_2786;
wire n_4547;
wire n_1566;
wire n_2837;
wire n_3765;
wire n_4058;
wire n_2006;
wire n_4090;
wire n_2446;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_2461;
wire n_2207;
wire n_2702;
wire n_1706;
wire n_3719;
wire n_4363;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3888;
wire n_3954;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_2529;
wire n_2238;
wire n_2374;
wire n_4103;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_2873;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_2278;
wire n_4028;
wire n_3330;
wire n_3514;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_4416;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4439;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_4575;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_4106;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_4581;
wire n_2960;
wire n_4260;
wire n_3270;
wire n_2323;
wire n_4549;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_4148;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_1736;
wire n_4512;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_4038;
wire n_4132;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_4500;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_2832;
wire n_1688;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_4515;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_2878;
wire n_1284;
wire n_1428;
wire n_1241;
wire n_3890;
wire n_3830;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_2782;
wire n_4136;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_4353;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_4567;
wire n_4176;
wire n_1207;
wire n_4124;
wire n_3606;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_3474;
wire n_2232;
wire n_4488;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_1512;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_3412;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_2988;
wire n_1636;
wire n_4560;
wire n_3482;
wire n_1900;
wire n_3948;
wire n_3230;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_4546;
wire n_1889;
wire n_1977;
wire n_2650;
wire n_1254;
wire n_3960;
wire n_4454;
wire n_4147;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_2332;
wire n_1703;
wire n_2391;
wire n_3828;
wire n_3975;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_3883;
wire n_4032;
wire n_4018;
wire n_4576;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_4117;
wire n_3049;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_2341;
wire n_2899;
wire n_1654;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_4572;
wire n_4505;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3739;
wire n_1840;
wire n_1230;
wire n_2739;
wire n_3728;
wire n_3962;
wire n_1597;
wire n_4082;
wire n_4476;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_4541;
wire n_4360;
wire n_1544;
wire n_3271;
wire n_4540;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_1267;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1790;
wire n_2956;
wire n_2382;
wire n_1354;
wire n_1213;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_4443;
wire n_1443;
wire n_4000;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_3458;
wire n_2727;
wire n_4562;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_2909;
wire n_1121;
wire n_1416;
wire n_1378;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1830;
wire n_3850;
wire n_4529;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_4498;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_2969;
wire n_1669;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_4432;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_4495;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_4357;
wire n_1594;
wire n_2806;
wire n_1935;
wire n_4109;
wire n_3191;
wire n_1716;
wire n_4108;
wire n_3777;
wire n_4502;
wire n_4530;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_3900;
wire n_4115;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_4394;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_2134;
wire n_3862;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_4513;
wire n_1179;
wire n_3284;
wire n_3909;
wire n_4311;
wire n_4220;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2810;
wire n_1386;
wire n_3391;
wire n_3506;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_2791;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_4378;
wire n_2683;
wire n_3212;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_4354;
wire n_4405;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_4459;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_3306;
wire n_2748;
wire n_2185;
wire n_4345;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_2398;
wire n_4233;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_1972;
wire n_1178;
wire n_2015;
wire n_2925;
wire n_1292;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_4029;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_2628;
wire n_1491;
wire n_3219;
wire n_3362;
wire n_3937;
wire n_4130;
wire n_2161;
wire n_1418;
wire n_4175;
wire n_1357;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_4456;
wire n_1312;
wire n_4508;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_1812;
wire n_3651;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_1880;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1567;
wire n_1343;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3629;
wire n_3666;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_2224;
wire n_1226;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_3046;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_4055;
wire n_3980;
wire n_4410;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_3741;
wire n_2388;
wire n_4352;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_2695;
wire n_2557;
wire n_2898;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_3567;
wire n_4003;
wire n_1832;
wire n_2795;
wire n_1392;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2762;
wire n_2302;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_4438;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_3884;
wire n_4433;
wire n_1147;
wire n_2829;
wire n_4367;
wire n_4492;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_4445;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_4254;
wire n_4462;
wire n_2507;
wire n_4219;
wire n_4484;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_2328;
wire n_4043;
wire n_4336;
wire n_4451;
wire n_2434;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_2649;
wire n_3981;
wire n_1247;
wire n_4234;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_2681;
wire n_1363;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3031;
wire n_3179;
wire n_2262;
wire n_2565;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_2980;
wire n_3078;
wire n_2335;
wire n_1728;
wire n_3699;
wire n_3971;
wire n_4315;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_4442;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_4494;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_4207;
wire n_4201;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_2312;
wire n_2677;
wire n_4296;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_3994;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1217;
wire n_2558;
wire n_2996;
wire n_1496;
wire n_2812;
wire n_1592;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_4386;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_4049;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_4522;
wire n_2718;
wire n_4263;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_4426;
wire n_3876;
wire n_3615;
wire n_4362;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_3946;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4089;
wire n_1501;
wire n_4186;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1198;
wire n_4096;
wire n_4506;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_1879;
wire n_1886;
wire n_4346;
wire n_4138;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_2476;
wire n_1365;
wire n_3968;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_2122;
wire n_1611;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_4337;
wire n_2399;
wire n_4543;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_4555;
wire n_1901;
wire n_2055;
wire n_4486;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_4359;
wire n_3118;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4441;
wire n_1906;
wire n_4323;
wire n_1899;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_4447;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_1467;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_4458;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_4523;
wire n_3007;
wire n_2267;
wire n_3599;
wire n_3618;
wire n_3705;
wire n_3983;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3286;
wire n_4480;
wire n_3734;
wire n_3370;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_4583;
wire n_3788;
wire n_3939;
wire n_2075;
wire n_3542;
wire n_3263;
wire n_1726;
wire n_3569;
wire n_3837;
wire n_2523;
wire n_1945;
wire n_3835;
wire n_2418;
wire n_2496;
wire n_1614;
wire n_1162;
wire n_1377;
wire n_2031;
wire n_3260;
wire n_3819;
wire n_3349;
wire n_3761;
wire n_3996;
wire n_4292;
wire n_2118;
wire n_3222;
wire n_1740;
wire n_1602;
wire n_4348;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_3764;
wire n_1553;
wire n_1760;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_1963;
wire n_2802;
wire n_4374;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_3403;
wire n_4261;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4344;
wire n_4084;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_1402;
wire n_1242;
wire n_3957;
wire n_2774;
wire n_2707;
wire n_2754;
wire n_4580;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_4393;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_1431;
wire n_4389;
wire n_3995;
wire n_1119;
wire n_4460;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_1500;
wire n_2214;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4461;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3501;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_3931;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_2949;
wire n_2894;
wire n_2300;
wire n_1667;
wire n_3896;
wire n_4067;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_4551;
wire n_3214;
wire n_3551;
wire n_4521;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_4525;
wire n_2283;
wire n_3364;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1219;
wire n_1711;
wire n_4387;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_4369;
wire n_2124;
wire n_1894;
wire n_2594;
wire n_1239;
wire n_1460;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_4324;
wire n_3626;
wire n_1898;
wire n_4428;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_4464;
wire n_4463;
wire n_1793;
wire n_4446;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1975;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_2119;
wire n_1719;
wire n_2742;
wire n_1540;
wire n_3671;
wire n_4396;
wire n_4440;
wire n_2366;
wire n_1797;
wire n_2493;
wire n_4425;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_4565;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_1800;
wire n_3791;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_4114;
wire n_2460;
wire n_4552;
wire n_2840;
wire n_1580;
wire n_3135;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_4482;
wire n_2480;
wire n_3024;
wire n_4528;
wire n_2772;
wire n_3564;
wire n_1700;
wire n_2637;
wire n_3795;
wire n_1332;
wire n_2306;
wire n_4328;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_3990;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_4400;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_3208;
wire n_3161;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4568;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_2958;
wire n_3365;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_4351;
wire n_4424;
wire n_3340;
wire n_4429;
wire n_4192;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_2581;
wire n_1527;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_4524;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_4221;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_4436;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_4035;
wire n_4160;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_3836;
wire n_4190;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_4545;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_2489;
wire n_1161;
wire n_3685;
wire n_4145;
wire n_3097;
wire n_4395;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_2492;
wire n_3864;
wire n_4385;
wire n_2939;
wire n_3425;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_2627;
wire n_1786;
wire n_4050;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_2106;
wire n_1804;
wire n_1406;
wire n_4306;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_4558;
wire n_1318;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2691;
wire n_2264;
wire n_3789;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_4511;
wire n_4358;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_4289;
wire n_1873;
wire n_1137;
wire n_1733;
wire n_2723;
wire n_1258;
wire n_1856;
wire n_1524;
wire n_1476;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_3925;
wire n_2928;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_3167;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3746;
wire n_4537;
wire n_1807;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3753;
wire n_3893;
wire n_2307;
wire n_1488;
wire n_1330;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_4076;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_2720;
wire n_1561;
wire n_2412;
wire n_1556;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_2907;
wire n_2386;
wire n_1971;
wire n_2945;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1324;
wire n_3543;
wire n_2528;
wire n_1778;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_1154;
wire n_3609;
wire n_1759;
wire n_1557;
wire n_2325;
wire n_1829;
wire n_4330;
wire n_1130;
wire n_1450;
wire n_4152;
wire n_3718;
wire n_2022;
wire n_3390;
wire n_3879;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_4343;
wire n_3017;
wire n_2320;
wire n_2986;
wire n_2570;
wire n_2329;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2890;
wire n_2546;
wire n_2454;
wire n_1493;
wire n_2813;
wire n_2911;
wire n_3381;
wire n_3455;
wire n_3736;
wire n_4466;
wire n_3313;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_3233;
wire n_1864;
wire n_2760;
wire n_3907;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_4419;
wire n_1151;
wire n_4420;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_3605;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4404;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_4372;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_4377;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_4563;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4301;
wire n_3573;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_4561;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_4188;
wire n_3654;
wire n_2001;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_4399;
wire n_2413;
wire n_4008;
wire n_2610;
wire n_1593;
wire n_3715;
wire n_4140;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_3982;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3973;
wire n_3134;
wire n_2771;
wire n_2403;
wire n_3842;
wire n_2947;
wire n_1367;
wire n_3755;
wire n_4202;
wire n_4536;
wire n_2044;
wire n_4534;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_3769;
wire n_4078;
wire n_2619;
wire n_1565;
wire n_4437;
wire n_1192;
wire n_3738;
wire n_3098;
wire n_1380;
wire n_4503;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_4070;
wire n_2020;
wire n_3987;
wire n_2310;
wire n_4249;
wire n_4418;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_3386;
wire n_4139;
wire n_4582;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_2177;
wire n_1511;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_4450;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3967;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_1517;
wire n_2036;
wire n_4412;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_4370;
wire n_3444;
wire n_4368;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_4091;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_4184;
wire n_4430;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_1752;
wire n_1955;
wire n_1504;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_4538;
wire n_4544;
wire n_1370;
wire n_1603;
wire n_4191;
wire n_4409;
wire n_4478;
wire n_2401;
wire n_2935;
wire n_4246;
wire n_3822;
wire n_4355;
wire n_3255;
wire n_3818;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_4061;
wire n_2658;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_4518;
wire n_4155;
wire n_3376;
wire n_4278;
wire n_4531;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_3770;
wire n_4375;
wire n_4542;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_2121;
wire n_1559;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_4532;
wire n_2692;
wire n_3927;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_2645;
wire n_2553;
wire n_1420;
wire n_3790;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_3490;
wire n_2459;
wire n_4413;
wire n_3396;
wire n_1210;
wire n_4241;
wire n_2751;
wire n_1135;
wire n_2566;
wire n_1622;
wire n_3113;
wire n_4183;
wire n_3101;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_4341;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3904;
wire n_3887;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_4126;
wire n_4164;
wire n_1336;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_1749;
wire n_1653;
wire n_3409;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4381;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_4469;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_4455;
wire n_3241;
wire n_3802;
wire n_3899;
wire n_4366;
wire n_1157;
wire n_1584;
wire n_4384;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_1814;
wire n_4577;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_4208;
wire n_3972;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_3926;
wire n_4209;
wire n_1687;
wire n_4457;
wire n_2073;
wire n_2150;
wire n_4481;
wire n_4004;
wire n_1552;
wire n_2938;
wire n_3630;
wire n_2498;
wire n_1612;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_4350;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_2455;
wire n_3092;
wire n_2600;
wire n_1617;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_2828;
wire n_4212;
wire n_4270;
wire n_1626;
wire n_3436;
wire n_4509;
wire n_4584;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_1175;
wire n_2299;
wire n_3751;
wire n_4388;
wire n_3402;
wire n_2406;
wire n_3247;
wire n_4477;
wire n_1621;
wire n_4110;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_1221;
wire n_4217;
wire n_1785;
wire n_1262;
wire n_4271;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_4317;
wire n_4406;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_2974;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_2503;
wire n_1758;
wire n_3873;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_2465;
wire n_1407;
wire n_3610;
wire n_2865;
wire n_1204;
wire n_1554;
wire n_3279;
wire n_2428;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_3178;
wire n_2858;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_3100;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3676;
wire n_1564;
wire n_2010;
wire n_3677;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_2356;
wire n_1361;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_2941;
wire n_1509;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_3536;
wire n_2564;
wire n_1721;
wire n_3576;
wire n_3558;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_3034;
wire n_1317;
wire n_1445;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_4435;
wire n_4053;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_3091;
wire n_4496;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_4210;
wire n_2604;
wire n_1775;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_4554;
wire n_2630;
wire n_4105;
wire n_4526;
wire n_2794;
wire n_3663;
wire n_2028;
wire n_3114;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_4578;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_2409;
wire n_1720;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_3360;
wire n_4470;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_1809;
wire n_2787;
wire n_4092;
wire n_3585;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_4057;
wire n_2770;
wire n_4550;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_4347;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3633;
wire n_3042;
wire n_4144;
wire n_4335;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_4379;
wire n_3111;
wire n_2212;
wire n_3838;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_4434;
wire n_2835;
wire n_1452;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_4499;
wire n_2569;
wire n_4504;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_2009;
wire n_4339;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_4497;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_4510;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4472;
wire n_4253;
wire n_1865;
wire n_1710;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_2580;
wire n_1792;
wire n_4064;
wire n_3351;
wire n_2062;
wire n_4489;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_2973;
wire n_2153;
wire n_1459;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_4519;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_4197;
wire n_4564;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_3776;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_4566;
wire n_3970;
wire n_4371;
wire n_2351;
wire n_1619;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_1902;
wire n_2206;
wire n_2784;
wire n_3898;
wire n_4414;
wire n_2541;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_4448;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_2538;
wire n_1845;
wire n_4295;
wire n_3932;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_4579;
wire n_4507;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_2552;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1470;
wire n_3445;
wire n_4087;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_4473;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_4398;
wire n_3253;
wire n_4471;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_4392;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_4238;
wire n_4365;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_4349;
wire n_3148;
wire n_3775;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3966;
wire n_4397;
wire n_4449;
wire n_3285;
wire n_3824;
wire n_3825;
wire n_4198;
wire n_2246;
wire n_3616;
wire n_1150;
wire n_4266;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_2971;
wire n_2532;
wire n_2191;
wire n_1831;
wire n_3874;
wire n_4373;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_4407;
wire n_2472;
wire n_2705;
wire n_2664;
wire n_4165;
wire n_4154;
wire n_4479;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_4390;
wire n_3845;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_4380;
wire n_4361;
wire n_3941;
wire n_1915;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_2240;
wire n_4168;
wire n_1369;
wire n_4258;
wire n_2846;
wire n_4298;
wire n_3371;
wire n_1781;
wire n_4571;
wire n_3137;
wire n_2917;
wire n_4250;
wire n_2544;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_4415;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_2188;
wire n_1777;
wire n_1477;
wire n_2097;
wire n_1982;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_2297;
wire n_1410;
wire n_4276;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_4408;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_4569;
wire n_1862;
wire n_2017;
wire n_3752;
wire n_4483;
wire n_3672;
wire n_3061;
wire n_1810;
wire n_2587;
wire n_3504;
wire n_2839;
wire n_1347;
wire n_3237;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_4128;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_4036;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_4487;
wire n_4548;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_4539;
wire n_4574;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_3071;
wire n_1638;
wire n_3918;
wire n_4010;
wire n_4329;
wire n_1571;
wire n_4501;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_2148;
wire n_1946;
wire n_3244;
wire n_4383;
wire n_3499;
wire n_4391;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_4095;
wire n_4444;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3910;
wire n_3947;
wire n_4485;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_2585;
wire n_1591;
wire n_3293;
wire n_3361;
wire n_2995;
wire n_4287;
wire n_4533;
wire n_1683;
wire n_1229;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_4356;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_2381;
wire n_1732;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_3707;
wire n_2052;
wire n_2485;
wire n_3779;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_4338;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_4573;
wire n_1891;
wire n_4520;
wire n_1328;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_4042;
wire n_1581;
wire n_3849;
wire n_4244;
wire n_1928;
wire n_3058;
wire n_2047;
wire n_4072;
wire n_2792;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_3398;
wire n_3709;
wire n_4465;
wire n_4553;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_1699;
wire n_1598;
wire n_3592;
wire n_3557;
wire n_3725;
wire n_3986;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_3399;
wire n_1702;
wire n_3894;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_3772;
wire n_1264;
wire n_2891;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_4120;
wire n_4149;
wire n_2361;
wire n_1313;
wire n_2819;
wire n_2880;
wire n_1115;
wire n_2229;
wire n_1722;
wire n_3030;
wire n_3075;
wire n_3505;
wire n_3722;
wire n_4277;
wire n_1339;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_2551;
wire n_2255;
wire n_4516;
wire n_1129;
wire n_2239;
wire n_1252;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_2830;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4222;
wire n_1871;
wire n_2514;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_3201;
wire n_1569;
wire n_3334;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1870;
wire n_1299;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_4046;
wire n_4467;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_4570;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_3041;
wire n_1251;
wire n_1989;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_1421;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_4493;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_4376;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_2479;
wire n_3204;
wire n_1981;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_2345;
wire n_4417;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g1108 ( 
.A(n_999),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_837),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1071),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1096),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1038),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_775),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_975),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_928),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_711),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_319),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_599),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_584),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_884),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_940),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_922),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_924),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_636),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_336),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1082),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_781),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_121),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_515),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_608),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_888),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_210),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_120),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_811),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_830),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1078),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1080),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1057),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_741),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_96),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_477),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1027),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_721),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_584),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_963),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_849),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_624),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_411),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_88),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1088),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_270),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_691),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_65),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1000),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_583),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_729),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_915),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1064),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_270),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1026),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_943),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_838),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_602),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_835),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_977),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_626),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_907),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1098),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1049),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_100),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_956),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_874),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_425),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_356),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_957),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_968),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1003),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1011),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_205),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1007),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_163),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_878),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_851),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_138),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_185),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_354),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1021),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1091),
.Y(n_1188)
);

BUFx10_ASAP7_75t_L g1189 ( 
.A(n_836),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1024),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_740),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_451),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_742),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_112),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_314),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1054),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1103),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_107),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_13),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_457),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_856),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_390),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_367),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_997),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_764),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_868),
.Y(n_1206)
);

CKINVDCx16_ASAP7_75t_R g1207 ( 
.A(n_274),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_396),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_921),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_4),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_746),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_735),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_978),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_616),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_538),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_783),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_942),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_846),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_326),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_933),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1001),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_40),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_245),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_630),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1101),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_923),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_209),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_479),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_189),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1029),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_400),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_868),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_391),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_468),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_945),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_446),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_115),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_670),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1061),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_505),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_771),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_351),
.Y(n_1242)
);

CKINVDCx16_ASAP7_75t_R g1243 ( 
.A(n_850),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_449),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_678),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_259),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1073),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_841),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_656),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1053),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_117),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_59),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_180),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_899),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_958),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_971),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_316),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_824),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_118),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_315),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_136),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_906),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_844),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_89),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_613),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_652),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_919),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1068),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_520),
.Y(n_1269)
);

BUFx5_ASAP7_75t_L g1270 ( 
.A(n_54),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_821),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_329),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_973),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_102),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_817),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_564),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1048),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_598),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_896),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_214),
.Y(n_1280)
);

INVxp67_ASAP7_75t_SL g1281 ( 
.A(n_1017),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_886),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_820),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1041),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_144),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_173),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_782),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_961),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_151),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_674),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_829),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_932),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_825),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_76),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_538),
.Y(n_1295)
);

CKINVDCx16_ASAP7_75t_R g1296 ( 
.A(n_1065),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_393),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_716),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_842),
.Y(n_1299)
);

BUFx5_ASAP7_75t_L g1300 ( 
.A(n_245),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_898),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_697),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_627),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1047),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_818),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_438),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1032),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1090),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_901),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1086),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_900),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_591),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_981),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1075),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_982),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_585),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_362),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1023),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1070),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_534),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_551),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_617),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_602),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_232),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_920),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_768),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_870),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_199),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_326),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_267),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1094),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1079),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_224),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_722),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1035),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_827),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_976),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_863),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_46),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1107),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1102),
.Y(n_1341)
);

CKINVDCx16_ASAP7_75t_R g1342 ( 
.A(n_804),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_481),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_986),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_828),
.Y(n_1345)
);

CKINVDCx16_ASAP7_75t_R g1346 ( 
.A(n_696),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_314),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_64),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_464),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1063),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_833),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_950),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_89),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_510),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1010),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_704),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_364),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_930),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_893),
.Y(n_1359)
);

CKINVDCx14_ASAP7_75t_R g1360 ( 
.A(n_1067),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_826),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_578),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_335),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1036),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_711),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_914),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_767),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_259),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_412),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_853),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_37),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_298),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_655),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_681),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_939),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_876),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_916),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_480),
.Y(n_1378)
);

CKINVDCx16_ASAP7_75t_R g1379 ( 
.A(n_1037),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_966),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_65),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_970),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_483),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_390),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_741),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_411),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_242),
.Y(n_1387)
);

BUFx10_ASAP7_75t_L g1388 ( 
.A(n_587),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_858),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_379),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1093),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_365),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_780),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_214),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_475),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_974),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_363),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_892),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_869),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_56),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_605),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1046),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_708),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_987),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_988),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_285),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_805),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_475),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_671),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_460),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_894),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_84),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_577),
.Y(n_1413)
);

BUFx5_ASAP7_75t_L g1414 ( 
.A(n_575),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_935),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_189),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_849),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_766),
.Y(n_1418)
);

CKINVDCx16_ASAP7_75t_R g1419 ( 
.A(n_745),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_492),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_684),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_790),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_905),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_953),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_854),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1059),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_573),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_40),
.Y(n_1428)
);

BUFx10_ASAP7_75t_L g1429 ( 
.A(n_885),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1052),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_359),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_33),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_464),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_263),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_347),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1008),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_807),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1015),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_993),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_173),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_840),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_879),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_823),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_949),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_995),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_269),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_182),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_882),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_598),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_881),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_56),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_642),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_430),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_817),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_128),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_445),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_632),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1055),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_877),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_927),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_772),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_394),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1072),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_349),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1033),
.Y(n_1465)
);

CKINVDCx14_ASAP7_75t_R g1466 ( 
.A(n_238),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_685),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_677),
.Y(n_1468)
);

BUFx10_ASAP7_75t_L g1469 ( 
.A(n_150),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_52),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1022),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_955),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_682),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1084),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_461),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_815),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_808),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1077),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_872),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_685),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1014),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_331),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_78),
.Y(n_1483)
);

CKINVDCx14_ASAP7_75t_R g1484 ( 
.A(n_443),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_679),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_960),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_887),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_647),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_839),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_827),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1092),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_607),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_288),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_447),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_403),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1004),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_121),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1016),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_374),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_190),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_865),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_242),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_965),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_829),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_36),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_343),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_133),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_810),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_848),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_771),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_426),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_235),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_600),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_309),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1006),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_349),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_228),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_951),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_57),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_655),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1018),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_859),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_193),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_917),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_135),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_897),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_783),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_738),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_392),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_864),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_809),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_830),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_86),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_421),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_225),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_92),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_248),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_238),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_80),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_952),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_185),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_271),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_702),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_269),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_298),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_524),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1062),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1039),
.Y(n_1548)
);

CKINVDCx16_ASAP7_75t_R g1549 ( 
.A(n_266),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_855),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_880),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_904),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1085),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1042),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_867),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_782),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_918),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_833),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_566),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_883),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_759),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_132),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_293),
.Y(n_1563)
);

BUFx10_ASAP7_75t_L g1564 ( 
.A(n_126),
.Y(n_1564)
);

CKINVDCx16_ASAP7_75t_R g1565 ( 
.A(n_211),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_292),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_183),
.Y(n_1567)
);

BUFx10_ASAP7_75t_L g1568 ( 
.A(n_1019),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1106),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_980),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_926),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_825),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_171),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1097),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_341),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_990),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_544),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_447),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_723),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1076),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_536),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_330),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_802),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1066),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_959),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_677),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_819),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_402),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_875),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_346),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_55),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_929),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_701),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_372),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_550),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_217),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_832),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_133),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_936),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_937),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_195),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_931),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_284),
.Y(n_1604)
);

BUFx10_ASAP7_75t_L g1605 ( 
.A(n_910),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_397),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1087),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_178),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_902),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_903),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_38),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_792),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_992),
.Y(n_1613)
);

INVxp33_ASAP7_75t_SL g1614 ( 
.A(n_53),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_82),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_10),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_599),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_363),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_311),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_97),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_9),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_623),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_969),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_271),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_4),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1028),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_913),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_444),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_813),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_962),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_534),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_805),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_733),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_600),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1009),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_142),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_486),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_454),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_765),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_847),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_967),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_588),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1020),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_372),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_590),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1013),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_67),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_806),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_636),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_842),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_786),
.Y(n_1651)
);

BUFx10_ASAP7_75t_L g1652 ( 
.A(n_1069),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_181),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_228),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_834),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_444),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1105),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_671),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_925),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_139),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_811),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_160),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_188),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1095),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_604),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1051),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_666),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_809),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1044),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_834),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_895),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_781),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_578),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1012),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_934),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_540),
.Y(n_1676)
);

BUFx5_ASAP7_75t_L g1677 ( 
.A(n_255),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_627),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_330),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1089),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_401),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1056),
.Y(n_1682)
);

CKINVDCx14_ASAP7_75t_R g1683 ( 
.A(n_588),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_707),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_192),
.Y(n_1685)
);

CKINVDCx16_ASAP7_75t_R g1686 ( 
.A(n_543),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1002),
.Y(n_1687)
);

CKINVDCx16_ASAP7_75t_R g1688 ( 
.A(n_404),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1050),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_0),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_726),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1104),
.Y(n_1692)
);

BUFx5_ASAP7_75t_L g1693 ( 
.A(n_743),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_177),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_279),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_954),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_670),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_801),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_857),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_891),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1034),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_909),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_137),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_712),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_796),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_994),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_241),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_323),
.Y(n_1708)
);

CKINVDCx16_ASAP7_75t_R g1709 ( 
.A(n_732),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_28),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_335),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1045),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_964),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_646),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_52),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_617),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_533),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_350),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_153),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_151),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_701),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_606),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_713),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_972),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_692),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1058),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_790),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_908),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_142),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_761),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_983),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_946),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_410),
.Y(n_1733)
);

CKINVDCx5p33_ASAP7_75t_R g1734 ( 
.A(n_768),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1099),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_488),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_742),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_388),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_637),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_948),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1074),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_633),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_748),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_348),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_773),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_865),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_989),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_149),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_667),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_55),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_71),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_938),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_816),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_663),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_991),
.Y(n_1756)
);

BUFx10_ASAP7_75t_L g1757 ( 
.A(n_784),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_859),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_862),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_375),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_268),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_780),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_712),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_226),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_614),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_92),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_686),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_493),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_223),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_365),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_375),
.Y(n_1771)
);

BUFx5_ASAP7_75t_L g1772 ( 
.A(n_401),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_574),
.Y(n_1773)
);

CKINVDCx20_ASAP7_75t_R g1774 ( 
.A(n_719),
.Y(n_1774)
);

BUFx10_ASAP7_75t_L g1775 ( 
.A(n_647),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_682),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_814),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_246),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_871),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_488),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1060),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_746),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_521),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_764),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_860),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1043),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_696),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_996),
.Y(n_1788)
);

INVxp33_ASAP7_75t_SL g1789 ( 
.A(n_873),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_50),
.Y(n_1790)
);

CKINVDCx20_ASAP7_75t_R g1791 ( 
.A(n_985),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_835),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_649),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_852),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1025),
.Y(n_1795)
);

BUFx10_ASAP7_75t_L g1796 ( 
.A(n_911),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_947),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_166),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_814),
.Y(n_1799)
);

BUFx2_ASAP7_75t_R g1800 ( 
.A(n_760),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_831),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_775),
.Y(n_1802)
);

BUFx10_ASAP7_75t_L g1803 ( 
.A(n_555),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_889),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_979),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_554),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_33),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_843),
.Y(n_1808)
);

INVx1_ASAP7_75t_SL g1809 ( 
.A(n_159),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_941),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_944),
.Y(n_1811)
);

BUFx8_ASAP7_75t_SL g1812 ( 
.A(n_209),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_747),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_861),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_619),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_984),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1083),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_550),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_215),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_998),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_767),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1081),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_735),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_845),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_607),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_890),
.Y(n_1826)
);

BUFx10_ASAP7_75t_L g1827 ( 
.A(n_721),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_380),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1030),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1031),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_162),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_738),
.Y(n_1832)
);

INVx4_ASAP7_75t_R g1833 ( 
.A(n_912),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_413),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_730),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_531),
.Y(n_1836)
);

INVxp33_ASAP7_75t_L g1837 ( 
.A(n_287),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_528),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_474),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_473),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_533),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_7),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_17),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_72),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_449),
.Y(n_1845)
);

BUFx10_ASAP7_75t_L g1846 ( 
.A(n_866),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_279),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_812),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_348),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_822),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_608),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_540),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_437),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1005),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_616),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_747),
.Y(n_1856)
);

CKINVDCx14_ASAP7_75t_R g1857 ( 
.A(n_1100),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1040),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_255),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_799),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_489),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_433),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1270),
.Y(n_1863)
);

CKINVDCx14_ASAP7_75t_R g1864 ( 
.A(n_1466),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1484),
.Y(n_1865)
);

INVxp33_ASAP7_75t_SL g1866 ( 
.A(n_1395),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1270),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1812),
.Y(n_1868)
);

BUFx3_ASAP7_75t_L g1869 ( 
.A(n_1255),
.Y(n_1869)
);

CKINVDCx20_ASAP7_75t_R g1870 ( 
.A(n_1683),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1270),
.Y(n_1871)
);

CKINVDCx16_ASAP7_75t_R g1872 ( 
.A(n_1207),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1426),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1270),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1243),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1270),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1800),
.Y(n_1877)
);

CKINVDCx14_ASAP7_75t_R g1878 ( 
.A(n_1360),
.Y(n_1878)
);

CKINVDCx16_ASAP7_75t_R g1879 ( 
.A(n_1342),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1429),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1546),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1300),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1346),
.Y(n_1883)
);

CKINVDCx20_ASAP7_75t_R g1884 ( 
.A(n_1282),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1300),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1300),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1300),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1300),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1414),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1414),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1419),
.Y(n_1891)
);

NOR2xp67_ASAP7_75t_L g1892 ( 
.A(n_1550),
.B(n_0),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1284),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1549),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1414),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1565),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1614),
.B(n_3),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1414),
.Y(n_1898)
);

INVxp67_ASAP7_75t_SL g1899 ( 
.A(n_1166),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1686),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1414),
.Y(n_1901)
);

CKINVDCx14_ASAP7_75t_R g1902 ( 
.A(n_1857),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1268),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1677),
.Y(n_1904)
);

CKINVDCx14_ASAP7_75t_R g1905 ( 
.A(n_1429),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1677),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1677),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1566),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1677),
.Y(n_1909)
);

CKINVDCx20_ASAP7_75t_R g1910 ( 
.A(n_1288),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1677),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1688),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1693),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1693),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1709),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1314),
.Y(n_1916)
);

INVxp67_ASAP7_75t_SL g1917 ( 
.A(n_1166),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1693),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1693),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1693),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1772),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1772),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1772),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1772),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1772),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1113),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1119),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1133),
.Y(n_1928)
);

INVxp33_ASAP7_75t_SL g1929 ( 
.A(n_1144),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1427),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1152),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1490),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1325),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1174),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1424),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1179),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1186),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1194),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1200),
.Y(n_1939)
);

INVxp33_ASAP7_75t_SL g1940 ( 
.A(n_1530),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1203),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1232),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1536),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1471),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1205),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1229),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1231),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1234),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1246),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1257),
.Y(n_1950)
);

INVxp33_ASAP7_75t_L g1951 ( 
.A(n_1624),
.Y(n_1951)
);

CKINVDCx16_ASAP7_75t_R g1952 ( 
.A(n_1296),
.Y(n_1952)
);

INVxp33_ASAP7_75t_L g1953 ( 
.A(n_1690),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1264),
.Y(n_1954)
);

INVxp67_ASAP7_75t_SL g1955 ( 
.A(n_1166),
.Y(n_1955)
);

INVxp33_ASAP7_75t_SL g1956 ( 
.A(n_1737),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1268),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1265),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1268),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1521),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1266),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1222),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1289),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1290),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1293),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1553),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1294),
.Y(n_1967)
);

HB1xp67_ASAP7_75t_L g1968 ( 
.A(n_1237),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1295),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1560),
.Y(n_1970)
);

CKINVDCx16_ASAP7_75t_R g1971 ( 
.A(n_1379),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1222),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1297),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1263),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1576),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1370),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1371),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1384),
.Y(n_1978)
);

BUFx10_ASAP7_75t_L g1979 ( 
.A(n_1222),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1979),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1903),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1899),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1917),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1955),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1876),
.A2(n_1114),
.B(n_1108),
.Y(n_1985)
);

INVx5_ASAP7_75t_L g1986 ( 
.A(n_1872),
.Y(n_1986)
);

BUFx3_ASAP7_75t_L g1987 ( 
.A(n_1979),
.Y(n_1987)
);

OAI22x1_ASAP7_75t_R g1988 ( 
.A1(n_1868),
.A2(n_1208),
.B1(n_1245),
.B2(n_1173),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1863),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1903),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1880),
.B(n_1441),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1968),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1903),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1867),
.Y(n_1994)
);

BUFx3_ASAP7_75t_L g1995 ( 
.A(n_1942),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1916),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1957),
.Y(n_1997)
);

OAI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1904),
.A2(n_1136),
.B(n_1126),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1875),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1883),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1957),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1871),
.Y(n_2002)
);

AND2x2_ASAP7_75t_SL g2003 ( 
.A(n_1952),
.B(n_1157),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1942),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1933),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1874),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1957),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1891),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1869),
.B(n_1533),
.Y(n_2009)
);

AOI22x1_ASAP7_75t_SL g2010 ( 
.A1(n_1884),
.A2(n_1271),
.B1(n_1278),
.B2(n_1269),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1894),
.Y(n_2011)
);

BUFx12f_ASAP7_75t_L g2012 ( 
.A(n_1935),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1896),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1878),
.B(n_1311),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1882),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1930),
.A2(n_1837),
.B1(n_1316),
.B2(n_1323),
.Y(n_2016)
);

INVx6_ASAP7_75t_L g2017 ( 
.A(n_1879),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1959),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1905),
.B(n_1568),
.Y(n_2019)
);

XOR2xp5_ASAP7_75t_L g2020 ( 
.A(n_1893),
.B(n_1779),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1959),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1959),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1910),
.Y(n_2023)
);

INVx5_ASAP7_75t_L g2024 ( 
.A(n_1971),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1864),
.B(n_1568),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1925),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1944),
.Y(n_2027)
);

OAI21x1_ASAP7_75t_L g2028 ( 
.A1(n_1885),
.A2(n_1168),
.B(n_1160),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1929),
.A2(n_1336),
.B1(n_1372),
.B2(n_1322),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1940),
.A2(n_1408),
.B1(n_1489),
.B2(n_1473),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1902),
.B(n_1605),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1960),
.Y(n_2032)
);

BUFx12f_ASAP7_75t_L g2033 ( 
.A(n_1970),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1951),
.B(n_1605),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1900),
.Y(n_2035)
);

INVx5_ASAP7_75t_L g2036 ( 
.A(n_1873),
.Y(n_2036)
);

INVx5_ASAP7_75t_L g2037 ( 
.A(n_1962),
.Y(n_2037)
);

INVx5_ASAP7_75t_L g2038 ( 
.A(n_1972),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1953),
.B(n_1652),
.Y(n_2039)
);

OAI22x1_ASAP7_75t_SL g2040 ( 
.A1(n_1956),
.A2(n_1597),
.B1(n_1599),
.B2(n_1539),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1926),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1974),
.B(n_1545),
.Y(n_2042)
);

AND2x6_ASAP7_75t_L g2043 ( 
.A(n_1927),
.B(n_1562),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1866),
.A2(n_1649),
.B1(n_1658),
.B2(n_1633),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1886),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1928),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1931),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1966),
.Y(n_2048)
);

BUFx8_ASAP7_75t_L g2049 ( 
.A(n_1934),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1936),
.Y(n_2050)
);

BUFx12f_ASAP7_75t_L g2051 ( 
.A(n_1912),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1932),
.B(n_1575),
.Y(n_2052)
);

INVx4_ASAP7_75t_L g2053 ( 
.A(n_1915),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1943),
.B(n_1652),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1887),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_1881),
.B(n_1604),
.Y(n_2056)
);

CKINVDCx20_ASAP7_75t_R g2057 ( 
.A(n_1975),
.Y(n_2057)
);

OA21x2_ASAP7_75t_L g2058 ( 
.A1(n_1888),
.A2(n_1176),
.B(n_1169),
.Y(n_2058)
);

BUFx3_ASAP7_75t_L g2059 ( 
.A(n_1889),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1890),
.Y(n_2060)
);

BUFx12f_ASAP7_75t_L g2061 ( 
.A(n_1865),
.Y(n_2061)
);

BUFx6f_ASAP7_75t_L g2062 ( 
.A(n_1937),
.Y(n_2062)
);

OA21x2_ASAP7_75t_L g2063 ( 
.A1(n_1895),
.A2(n_1190),
.B(n_1182),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1898),
.Y(n_2064)
);

AOI22x1_ASAP7_75t_SL g2065 ( 
.A1(n_1877),
.A2(n_1665),
.B1(n_1678),
.B2(n_1660),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1901),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1906),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1907),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1909),
.Y(n_2069)
);

HB1xp67_ASAP7_75t_L g2070 ( 
.A(n_1908),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1911),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1938),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1939),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1913),
.Y(n_2074)
);

BUFx8_ASAP7_75t_L g2075 ( 
.A(n_1941),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1945),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1914),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1918),
.B(n_1789),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1919),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1946),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1920),
.Y(n_2081)
);

BUFx12f_ASAP7_75t_L g2082 ( 
.A(n_1870),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1921),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_1947),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1922),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1948),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1949),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1923),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1897),
.A2(n_1774),
.B1(n_1840),
.B2(n_1710),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1924),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1950),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1954),
.B(n_1784),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1958),
.Y(n_2093)
);

INVxp67_ASAP7_75t_L g2094 ( 
.A(n_1961),
.Y(n_2094)
);

BUFx12f_ASAP7_75t_L g2095 ( 
.A(n_1892),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1963),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1964),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1965),
.B(n_1217),
.Y(n_2098)
);

INVx2_ASAP7_75t_SL g2099 ( 
.A(n_1967),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_1969),
.B(n_1806),
.Y(n_2100)
);

BUFx12f_ASAP7_75t_L g2101 ( 
.A(n_1973),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1976),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1977),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1978),
.Y(n_2104)
);

OAI21x1_ASAP7_75t_L g2105 ( 
.A1(n_1876),
.A2(n_1225),
.B(n_1221),
.Y(n_2105)
);

OAI22x1_ASAP7_75t_L g2106 ( 
.A1(n_1877),
.A2(n_1212),
.B1(n_1367),
.B2(n_1287),
.Y(n_2106)
);

INVx2_ASAP7_75t_SL g2107 ( 
.A(n_1880),
.Y(n_2107)
);

INVx5_ASAP7_75t_L g2108 ( 
.A(n_1872),
.Y(n_2108)
);

INVx3_ASAP7_75t_L g2109 ( 
.A(n_1979),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1899),
.Y(n_2110)
);

BUFx12f_ASAP7_75t_L g2111 ( 
.A(n_1868),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1903),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1899),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1875),
.Y(n_2114)
);

AND2x6_ASAP7_75t_L g2115 ( 
.A(n_1880),
.B(n_1814),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1899),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1979),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1899),
.Y(n_2118)
);

INVx5_ASAP7_75t_L g2119 ( 
.A(n_1979),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1929),
.A2(n_1791),
.B1(n_1519),
.B2(n_1584),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1979),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1903),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_1979),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_1875),
.Y(n_2124)
);

INVx2_ASAP7_75t_SL g2125 ( 
.A(n_1880),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1979),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1905),
.B(n_1796),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1878),
.B(n_1230),
.Y(n_2128)
);

BUFx12f_ASAP7_75t_L g2129 ( 
.A(n_1868),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1905),
.B(n_1796),
.Y(n_2130)
);

AOI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_1929),
.A2(n_1715),
.B1(n_1760),
.B2(n_1457),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_1880),
.B(n_1236),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_1875),
.Y(n_2133)
);

OAI22x1_ASAP7_75t_L g2134 ( 
.A1(n_1877),
.A2(n_1790),
.B1(n_1809),
.B2(n_1793),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_1880),
.B(n_1356),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1916),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1903),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1903),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1979),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1880),
.B(n_1180),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1979),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1905),
.B(n_1189),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1880),
.B(n_1383),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1899),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_1875),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1979),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_1979),
.Y(n_2147)
);

CKINVDCx16_ASAP7_75t_R g2148 ( 
.A(n_1952),
.Y(n_2148)
);

BUFx12f_ASAP7_75t_L g2149 ( 
.A(n_1868),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1979),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1899),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_1875),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1899),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1903),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1878),
.B(n_1235),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_1979),
.Y(n_2156)
);

INVxp67_ASAP7_75t_SL g2157 ( 
.A(n_1974),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1899),
.Y(n_2158)
);

INVx6_ASAP7_75t_L g2159 ( 
.A(n_1979),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1880),
.B(n_1443),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1899),
.Y(n_2161)
);

CKINVDCx20_ASAP7_75t_R g2162 ( 
.A(n_1884),
.Y(n_2162)
);

INVxp67_ASAP7_75t_L g2163 ( 
.A(n_1968),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_L g2164 ( 
.A1(n_1876),
.A2(n_1273),
.B(n_1250),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1899),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_1979),
.Y(n_2166)
);

OAI21x1_ASAP7_75t_L g2167 ( 
.A1(n_1876),
.A2(n_1308),
.B(n_1304),
.Y(n_2167)
);

BUFx3_ASAP7_75t_L g2168 ( 
.A(n_1979),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1899),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1899),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1905),
.B(n_1189),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1899),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1903),
.Y(n_2173)
);

INVx2_ASAP7_75t_SL g2174 ( 
.A(n_1880),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1905),
.B(n_1388),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_1875),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1905),
.B(n_1388),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_1916),
.Y(n_2178)
);

INVx2_ASAP7_75t_SL g2179 ( 
.A(n_1880),
.Y(n_2179)
);

BUFx12f_ASAP7_75t_L g2180 ( 
.A(n_1868),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1899),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1903),
.Y(n_2182)
);

INVx4_ASAP7_75t_L g2183 ( 
.A(n_1880),
.Y(n_2183)
);

AOI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_1929),
.A2(n_1828),
.B1(n_1849),
.B2(n_1821),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_1929),
.A2(n_1116),
.B1(n_1117),
.B2(n_1109),
.Y(n_2185)
);

AOI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_1929),
.A2(n_1127),
.B1(n_1128),
.B2(n_1124),
.Y(n_2186)
);

BUFx3_ASAP7_75t_L g2187 ( 
.A(n_1979),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1899),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_1875),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1903),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1899),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1903),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_1875),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1905),
.B(n_1469),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1916),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1979),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_L g2197 ( 
.A(n_1979),
.Y(n_2197)
);

AOI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_1929),
.A2(n_1129),
.B1(n_1132),
.B2(n_1130),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_1880),
.B(n_1513),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1899),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_1968),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1903),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1905),
.B(n_1469),
.Y(n_2203)
);

BUFx8_ASAP7_75t_L g2204 ( 
.A(n_1880),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1878),
.B(n_1309),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1905),
.B(n_1564),
.Y(n_2206)
);

BUFx6f_ASAP7_75t_L g2207 ( 
.A(n_1979),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_1875),
.Y(n_2208)
);

BUFx6f_ASAP7_75t_L g2209 ( 
.A(n_1979),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1903),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1903),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1899),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1878),
.B(n_1310),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1878),
.B(n_1313),
.Y(n_2214)
);

AND2x2_ASAP7_75t_SL g2215 ( 
.A(n_1952),
.B(n_1118),
.Y(n_2215)
);

INVxp67_ASAP7_75t_SL g2216 ( 
.A(n_1974),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_1979),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1899),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1979),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1899),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_1880),
.B(n_1795),
.Y(n_2221)
);

INVx2_ASAP7_75t_SL g2222 ( 
.A(n_1880),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_1905),
.B(n_1564),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1899),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1903),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1905),
.B(n_1757),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1878),
.B(n_1315),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_1979),
.Y(n_2228)
);

CKINVDCx20_ASAP7_75t_R g2229 ( 
.A(n_1884),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_1880),
.B(n_1591),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1979),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_1875),
.Y(n_2232)
);

HB1xp67_ASAP7_75t_L g2233 ( 
.A(n_1875),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1876),
.A2(n_1341),
.B(n_1337),
.Y(n_2234)
);

INVx5_ASAP7_75t_L g2235 ( 
.A(n_1979),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_1875),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_1880),
.B(n_1733),
.Y(n_2237)
);

OAI22x1_ASAP7_75t_R g2238 ( 
.A1(n_1868),
.A2(n_1134),
.B1(n_1139),
.B2(n_1135),
.Y(n_2238)
);

AOI22x1_ASAP7_75t_SL g2239 ( 
.A1(n_1884),
.A2(n_1141),
.B1(n_1143),
.B2(n_1140),
.Y(n_2239)
);

OAI22x1_ASAP7_75t_R g2240 ( 
.A1(n_1868),
.A2(n_1146),
.B1(n_1148),
.B2(n_1147),
.Y(n_2240)
);

INVx4_ASAP7_75t_L g2241 ( 
.A(n_1880),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1929),
.A2(n_1153),
.B1(n_1155),
.B2(n_1149),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1899),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_1979),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_1875),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1878),
.B(n_1344),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_1979),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1979),
.Y(n_2248)
);

AOI22x1_ASAP7_75t_SL g2249 ( 
.A1(n_1884),
.A2(n_1156),
.B1(n_1163),
.B2(n_1159),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1899),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1989),
.B(n_1570),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1996),
.Y(n_2252)
);

AND2x4_ASAP7_75t_SL g2253 ( 
.A(n_2142),
.B(n_1757),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2091),
.Y(n_2254)
);

OA21x2_ASAP7_75t_L g2255 ( 
.A1(n_2028),
.A2(n_1998),
.B(n_1985),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2093),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1994),
.B(n_1112),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2102),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2022),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_2117),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2103),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2026),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1981),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2041),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2002),
.B(n_1171),
.Y(n_2265)
);

HB1xp67_ASAP7_75t_L g2266 ( 
.A(n_2005),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_1986),
.B(n_2108),
.Y(n_2267)
);

BUFx6f_ASAP7_75t_L g2268 ( 
.A(n_2121),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2046),
.Y(n_2269)
);

OA21x2_ASAP7_75t_L g2270 ( 
.A1(n_2105),
.A2(n_1352),
.B(n_1350),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2006),
.B(n_1279),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1990),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_2139),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2047),
.Y(n_2274)
);

INVx3_ASAP7_75t_L g2275 ( 
.A(n_1995),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1993),
.Y(n_2276)
);

OR2x2_ASAP7_75t_SL g2277 ( 
.A(n_2148),
.B(n_1151),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2015),
.B(n_2060),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2001),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_1980),
.B(n_1125),
.Y(n_2280)
);

OAI21x1_ASAP7_75t_L g2281 ( 
.A1(n_2164),
.A2(n_1382),
.B(n_1364),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2050),
.Y(n_2282)
);

BUFx8_ASAP7_75t_L g2283 ( 
.A(n_2111),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2064),
.B(n_1335),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_2141),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2062),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_2027),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_2032),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2072),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_2146),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_1987),
.B(n_1729),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2076),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2080),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2147),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2018),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_2156),
.B(n_1390),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2021),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2084),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_2196),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2112),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2034),
.B(n_1775),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2086),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2122),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2087),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2166),
.B(n_1394),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_2197),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2096),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_L g2308 ( 
.A(n_2207),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2137),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_SL g2310 ( 
.A(n_2003),
.B(n_1775),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2097),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2067),
.B(n_1458),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2071),
.B(n_1486),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2104),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2079),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2083),
.Y(n_2316)
);

OAI21x1_ASAP7_75t_L g2317 ( 
.A1(n_2167),
.A2(n_1396),
.B(n_1391),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_2209),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2085),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2088),
.Y(n_2320)
);

OR2x6_ASAP7_75t_L g2321 ( 
.A(n_2017),
.B(n_1162),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2136),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2168),
.B(n_1401),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2090),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1982),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1983),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1984),
.Y(n_2327)
);

INVx3_ASAP7_75t_L g2328 ( 
.A(n_2219),
.Y(n_2328)
);

INVx3_ASAP7_75t_L g2329 ( 
.A(n_2228),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2138),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2110),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2154),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2113),
.Y(n_2333)
);

BUFx6f_ASAP7_75t_L g2334 ( 
.A(n_1997),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2116),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2118),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2078),
.B(n_2055),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_2004),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_2007),
.Y(n_2339)
);

INVxp67_ASAP7_75t_L g2340 ( 
.A(n_2039),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2144),
.Y(n_2341)
);

INVx3_ASAP7_75t_L g2342 ( 
.A(n_2159),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2173),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2151),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_1992),
.B(n_1803),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2153),
.Y(n_2346)
);

AND2x6_ASAP7_75t_L g2347 ( 
.A(n_2019),
.B(n_1353),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_2178),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2158),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2161),
.Y(n_2350)
);

BUFx6f_ASAP7_75t_L g2351 ( 
.A(n_2187),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2182),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2165),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2169),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2190),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2192),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2170),
.Y(n_2357)
);

NAND3xp33_ASAP7_75t_L g2358 ( 
.A(n_2094),
.B(n_2186),
.C(n_2185),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2172),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2202),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2059),
.B(n_2069),
.Y(n_2361)
);

BUFx2_ASAP7_75t_L g2362 ( 
.A(n_2195),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2163),
.B(n_1803),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2107),
.B(n_1164),
.Y(n_2364)
);

HB1xp67_ASAP7_75t_L g2365 ( 
.A(n_2070),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_2101),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2201),
.Y(n_2367)
);

INVx3_ASAP7_75t_L g2368 ( 
.A(n_2217),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2181),
.Y(n_2369)
);

OAI21x1_ASAP7_75t_L g2370 ( 
.A1(n_2234),
.A2(n_1404),
.B(n_1402),
.Y(n_2370)
);

HB1xp67_ASAP7_75t_L g2371 ( 
.A(n_2008),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_2231),
.B(n_1433),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2054),
.B(n_1827),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2188),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2191),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2210),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2045),
.B(n_1110),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2066),
.B(n_1111),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2119),
.Y(n_2379)
);

BUFx6f_ASAP7_75t_L g2380 ( 
.A(n_2119),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2013),
.Y(n_2381)
);

INVx3_ASAP7_75t_L g2382 ( 
.A(n_2073),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2024),
.B(n_1437),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2211),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2200),
.Y(n_2385)
);

BUFx6f_ASAP7_75t_L g2386 ( 
.A(n_2235),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2225),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2068),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2074),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2212),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2077),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2127),
.B(n_2130),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2171),
.B(n_1827),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2081),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_2114),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2218),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2175),
.B(n_1846),
.Y(n_2397)
);

OAI21x1_ASAP7_75t_L g2398 ( 
.A1(n_2058),
.A2(n_1423),
.B(n_1405),
.Y(n_2398)
);

AOI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2198),
.A2(n_1181),
.B1(n_1184),
.B2(n_1170),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2220),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2024),
.B(n_1447),
.Y(n_2401)
);

NOR2xp33_ASAP7_75t_L g2402 ( 
.A(n_2128),
.B(n_2155),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_2205),
.B(n_1442),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2224),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2157),
.B(n_1115),
.Y(n_2405)
);

OA21x2_ASAP7_75t_L g2406 ( 
.A1(n_2213),
.A2(n_1463),
.B(n_1459),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2243),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_2235),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2177),
.B(n_1846),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2250),
.Y(n_2410)
);

INVx4_ASAP7_75t_L g2411 ( 
.A(n_2109),
.Y(n_2411)
);

INVx3_ASAP7_75t_L g2412 ( 
.A(n_2123),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2099),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2194),
.B(n_1451),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2063),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2098),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2092),
.Y(n_2417)
);

INVx3_ASAP7_75t_L g2418 ( 
.A(n_2126),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_2129),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2100),
.Y(n_2420)
);

NAND2xp33_ASAP7_75t_SL g2421 ( 
.A(n_2053),
.B(n_1185),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2037),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2037),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2038),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2216),
.Y(n_2425)
);

BUFx2_ASAP7_75t_L g2426 ( 
.A(n_2145),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2140),
.B(n_1120),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2125),
.B(n_1453),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2038),
.Y(n_2429)
);

OAI22xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2030),
.A2(n_2089),
.B1(n_2044),
.B2(n_2029),
.Y(n_2430)
);

INVx3_ASAP7_75t_L g2431 ( 
.A(n_2150),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2042),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_2244),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_L g2434 ( 
.A(n_2051),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2247),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2248),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2221),
.B(n_1121),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2174),
.B(n_1454),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2031),
.B(n_1122),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2214),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2227),
.Y(n_2441)
);

BUFx6f_ASAP7_75t_L g2442 ( 
.A(n_2149),
.Y(n_2442)
);

NAND2x1_ASAP7_75t_L g2443 ( 
.A(n_2115),
.B(n_1833),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1991),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2246),
.Y(n_2445)
);

HB1xp67_ASAP7_75t_L g2446 ( 
.A(n_2152),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_2180),
.Y(n_2447)
);

INVx2_ASAP7_75t_SL g2448 ( 
.A(n_2203),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_2009),
.Y(n_2449)
);

INVx1_ASAP7_75t_SL g2450 ( 
.A(n_2023),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2132),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2135),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2025),
.B(n_1123),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2057),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2043),
.B(n_1131),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2014),
.B(n_1465),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_2012),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2143),
.Y(n_2458)
);

HB1xp67_ASAP7_75t_L g2459 ( 
.A(n_2189),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_2033),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2043),
.B(n_2179),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2095),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2160),
.Y(n_2463)
);

AND2x4_ASAP7_75t_L g2464 ( 
.A(n_2222),
.B(n_1456),
.Y(n_2464)
);

AND2x6_ASAP7_75t_L g2465 ( 
.A(n_2206),
.B(n_1353),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2199),
.B(n_1137),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2230),
.Y(n_2467)
);

INVx1_ASAP7_75t_SL g2468 ( 
.A(n_2162),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2223),
.B(n_1467),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2226),
.B(n_1475),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2237),
.Y(n_2471)
);

CKINVDCx14_ASAP7_75t_R g2472 ( 
.A(n_2229),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2115),
.B(n_1138),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2183),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_2036),
.Y(n_2475)
);

BUFx6f_ASAP7_75t_L g2476 ( 
.A(n_2036),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2061),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2056),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2241),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2052),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_2048),
.Y(n_2481)
);

BUFx6f_ASAP7_75t_L g2482 ( 
.A(n_2082),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_1999),
.B(n_1480),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2215),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2242),
.B(n_1142),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2131),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2184),
.B(n_1145),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2120),
.B(n_1150),
.Y(n_2488)
);

BUFx2_ASAP7_75t_L g2489 ( 
.A(n_2000),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2011),
.B(n_1158),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2342),
.B(n_2035),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2262),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2402),
.B(n_2124),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2260),
.Y(n_2494)
);

AOI22xp33_ASAP7_75t_L g2495 ( 
.A1(n_2430),
.A2(n_2016),
.B1(n_2134),
.B2(n_2106),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2419),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2325),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2388),
.Y(n_2498)
);

NOR3xp33_ASAP7_75t_L g2499 ( 
.A(n_2395),
.B(n_2426),
.C(n_2489),
.Y(n_2499)
);

INVxp67_ASAP7_75t_L g2500 ( 
.A(n_2371),
.Y(n_2500)
);

INVx3_ASAP7_75t_L g2501 ( 
.A(n_2260),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2389),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2326),
.Y(n_2503)
);

OA22x2_ASAP7_75t_L g2504 ( 
.A1(n_2486),
.A2(n_2020),
.B1(n_2176),
.B2(n_2133),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_R g2505 ( 
.A(n_2252),
.B(n_2193),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2391),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2394),
.Y(n_2507)
);

INVx2_ASAP7_75t_SL g2508 ( 
.A(n_2381),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2327),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2331),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2254),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2333),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_2440),
.B(n_2208),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2256),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2335),
.Y(n_2515)
);

BUFx4f_ASAP7_75t_L g2516 ( 
.A(n_2442),
.Y(n_2516)
);

AND2x2_ASAP7_75t_SL g2517 ( 
.A(n_2310),
.B(n_2232),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2441),
.A2(n_2236),
.B1(n_2245),
.B2(n_2233),
.Y(n_2518)
);

INVx8_ASAP7_75t_L g2519 ( 
.A(n_2267),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2416),
.B(n_1353),
.Y(n_2520)
);

INVx2_ASAP7_75t_SL g2521 ( 
.A(n_2446),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2258),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2261),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2336),
.Y(n_2524)
);

INVxp67_ASAP7_75t_SL g2525 ( 
.A(n_2268),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2341),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2263),
.Y(n_2527)
);

INVx2_ASAP7_75t_SL g2528 ( 
.A(n_2459),
.Y(n_2528)
);

AOI22xp33_ASAP7_75t_L g2529 ( 
.A1(n_2445),
.A2(n_1224),
.B1(n_1240),
.B2(n_1183),
.Y(n_2529)
);

CKINVDCx5p33_ASAP7_75t_R g2530 ( 
.A(n_2287),
.Y(n_2530)
);

OAI22xp5_ASAP7_75t_L g2531 ( 
.A1(n_2358),
.A2(n_1191),
.B1(n_1193),
.B2(n_1192),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2272),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2276),
.Y(n_2533)
);

BUFx8_ASAP7_75t_SL g2534 ( 
.A(n_2362),
.Y(n_2534)
);

INVx2_ASAP7_75t_SL g2535 ( 
.A(n_2268),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2279),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2344),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2373),
.B(n_2367),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_2481),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2295),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2346),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2273),
.Y(n_2542)
);

NAND2xp33_ASAP7_75t_L g2543 ( 
.A(n_2337),
.B(n_2427),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2349),
.Y(n_2544)
);

AOI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2456),
.A2(n_1281),
.B1(n_1481),
.B2(n_1472),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2350),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2403),
.B(n_1417),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2353),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2273),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2297),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2354),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_SL g2552 ( 
.A(n_2340),
.B(n_2411),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2300),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2439),
.B(n_2049),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_2472),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_L g2556 ( 
.A(n_2485),
.B(n_2204),
.Y(n_2556)
);

AOI22xp33_ASAP7_75t_SL g2557 ( 
.A1(n_2488),
.A2(n_2010),
.B1(n_2249),
.B2(n_2239),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2301),
.A2(n_1526),
.B1(n_1551),
.B2(n_1503),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2453),
.B(n_2075),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2357),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2303),
.Y(n_2561)
);

AOI22xp33_ASAP7_75t_L g2562 ( 
.A1(n_2315),
.A2(n_1406),
.B1(n_1416),
.B2(n_1285),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2484),
.B(n_1195),
.Y(n_2563)
);

INVx2_ASAP7_75t_SL g2564 ( 
.A(n_2306),
.Y(n_2564)
);

AOI22xp33_ASAP7_75t_L g2565 ( 
.A1(n_2316),
.A2(n_1425),
.B1(n_1483),
.B2(n_1434),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_2306),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2359),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2400),
.B(n_1417),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_L g2569 ( 
.A1(n_2319),
.A2(n_1561),
.B1(n_1787),
.B2(n_1512),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_2283),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2320),
.B(n_1417),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2345),
.B(n_1485),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2363),
.B(n_1493),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2369),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_L g2575 ( 
.A(n_2425),
.B(n_1198),
.Y(n_2575)
);

AOI22xp33_ASAP7_75t_L g2576 ( 
.A1(n_2324),
.A2(n_1819),
.B1(n_1832),
.B2(n_1802),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2374),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2309),
.Y(n_2578)
);

NAND2xp33_ASAP7_75t_L g2579 ( 
.A(n_2437),
.B(n_1199),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2330),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2375),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2385),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2390),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2368),
.B(n_1201),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2332),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2396),
.Y(n_2586)
);

INVx5_ASAP7_75t_L g2587 ( 
.A(n_2442),
.Y(n_2587)
);

BUFx2_ASAP7_75t_L g2588 ( 
.A(n_2365),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2404),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2308),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2343),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2352),
.Y(n_2592)
);

INVxp67_ASAP7_75t_SL g2593 ( 
.A(n_2308),
.Y(n_2593)
);

INVx5_ASAP7_75t_L g2594 ( 
.A(n_2447),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2407),
.B(n_1431),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2487),
.B(n_1202),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2410),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2450),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2311),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_2266),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2314),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2318),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2406),
.A2(n_1859),
.B1(n_1578),
.B2(n_1647),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2449),
.B(n_1206),
.Y(n_2604)
);

NAND2xp33_ASAP7_75t_SL g2605 ( 
.A(n_2288),
.B(n_1210),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2278),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2355),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2356),
.Y(n_2608)
);

NOR3xp33_ASAP7_75t_L g2609 ( 
.A(n_2322),
.B(n_2348),
.C(n_2412),
.Y(n_2609)
);

OR2x6_ASAP7_75t_L g2610 ( 
.A(n_2447),
.B(n_1988),
.Y(n_2610)
);

INVx3_ASAP7_75t_L g2611 ( 
.A(n_2318),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2393),
.B(n_2397),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2360),
.Y(n_2613)
);

NOR2xp33_ASAP7_75t_L g2614 ( 
.A(n_2418),
.B(n_2431),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2251),
.B(n_1431),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2376),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2384),
.Y(n_2617)
);

OAI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2413),
.A2(n_1211),
.B1(n_1215),
.B2(n_1214),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2433),
.B(n_1216),
.Y(n_2619)
);

INVxp67_ASAP7_75t_L g2620 ( 
.A(n_2454),
.Y(n_2620)
);

INVx5_ASAP7_75t_L g2621 ( 
.A(n_2434),
.Y(n_2621)
);

INVxp33_ASAP7_75t_SL g2622 ( 
.A(n_2468),
.Y(n_2622)
);

OAI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2399),
.A2(n_2382),
.B1(n_2452),
.B2(n_2451),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2387),
.Y(n_2624)
);

OR2x2_ASAP7_75t_L g2625 ( 
.A(n_2321),
.B(n_1494),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_L g2626 ( 
.A(n_2448),
.B(n_1218),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2259),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2409),
.B(n_1499),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2415),
.Y(n_2629)
);

BUFx10_ASAP7_75t_L g2630 ( 
.A(n_2434),
.Y(n_2630)
);

INVx4_ASAP7_75t_L g2631 ( 
.A(n_2457),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2366),
.B(n_2462),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2270),
.Y(n_2633)
);

NAND3xp33_ASAP7_75t_L g2634 ( 
.A(n_2490),
.B(n_1223),
.C(n_1219),
.Y(n_2634)
);

INVx2_ASAP7_75t_SL g2635 ( 
.A(n_2392),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2338),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2414),
.B(n_2469),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2422),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2423),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2280),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2424),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2429),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_2351),
.B(n_1227),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2351),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_2361),
.B(n_1228),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_SL g2646 ( 
.A(n_2457),
.Y(n_2646)
);

AOI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2470),
.A2(n_1571),
.B1(n_1574),
.B2(n_1554),
.Y(n_2647)
);

NAND2xp33_ASAP7_75t_L g2648 ( 
.A(n_2435),
.B(n_1233),
.Y(n_2648)
);

INVx5_ASAP7_75t_L g2649 ( 
.A(n_2460),
.Y(n_2649)
);

OR2x2_ASAP7_75t_L g2650 ( 
.A(n_2478),
.B(n_1502),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2405),
.B(n_1238),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2398),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_2460),
.Y(n_2653)
);

INVx2_ASAP7_75t_SL g2654 ( 
.A(n_2428),
.Y(n_2654)
);

INVx6_ASAP7_75t_L g2655 ( 
.A(n_2462),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2629),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2497),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2493),
.B(n_2347),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2516),
.Y(n_2659)
);

INVx3_ASAP7_75t_L g2660 ( 
.A(n_2630),
.Y(n_2660)
);

INVx3_ASAP7_75t_L g2661 ( 
.A(n_2496),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2566),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2503),
.Y(n_2663)
);

INVx2_ASAP7_75t_SL g2664 ( 
.A(n_2519),
.Y(n_2664)
);

BUFx2_ASAP7_75t_L g2665 ( 
.A(n_2588),
.Y(n_2665)
);

OAI221xp5_ASAP7_75t_L g2666 ( 
.A1(n_2495),
.A2(n_2458),
.B1(n_2467),
.B2(n_2471),
.C(n_2463),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2509),
.Y(n_2667)
);

BUFx2_ASAP7_75t_L g2668 ( 
.A(n_2598),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_2530),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2510),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2492),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2566),
.Y(n_2672)
);

BUFx2_ASAP7_75t_L g2673 ( 
.A(n_2508),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2498),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2512),
.Y(n_2675)
);

BUFx2_ASAP7_75t_L g2676 ( 
.A(n_2521),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2515),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2606),
.B(n_2347),
.Y(n_2678)
);

BUFx6f_ASAP7_75t_L g2679 ( 
.A(n_2519),
.Y(n_2679)
);

BUFx4_ASAP7_75t_L g2680 ( 
.A(n_2646),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2524),
.Y(n_2681)
);

HB1xp67_ASAP7_75t_L g2682 ( 
.A(n_2528),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2502),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2506),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2526),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2537),
.Y(n_2686)
);

HB1xp67_ASAP7_75t_L g2687 ( 
.A(n_2500),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2541),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_2505),
.B(n_2438),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2620),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2544),
.Y(n_2691)
);

INVx4_ASAP7_75t_L g2692 ( 
.A(n_2587),
.Y(n_2692)
);

AND2x6_ASAP7_75t_L g2693 ( 
.A(n_2612),
.B(n_2477),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2546),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2548),
.Y(n_2695)
);

AND2x6_ASAP7_75t_L g2696 ( 
.A(n_2653),
.B(n_2477),
.Y(n_2696)
);

INVx5_ASAP7_75t_L g2697 ( 
.A(n_2534),
.Y(n_2697)
);

AOI22xp33_ASAP7_75t_SL g2698 ( 
.A1(n_2517),
.A2(n_2065),
.B1(n_2465),
.B2(n_2253),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2622),
.B(n_2275),
.Y(n_2699)
);

BUFx6f_ASAP7_75t_L g2700 ( 
.A(n_2587),
.Y(n_2700)
);

INVx4_ASAP7_75t_L g2701 ( 
.A(n_2594),
.Y(n_2701)
);

BUFx3_ASAP7_75t_L g2702 ( 
.A(n_2594),
.Y(n_2702)
);

NAND3x1_ASAP7_75t_L g2703 ( 
.A(n_2499),
.B(n_2040),
.C(n_2461),
.Y(n_2703)
);

BUFx3_ASAP7_75t_L g2704 ( 
.A(n_2621),
.Y(n_2704)
);

BUFx6f_ASAP7_75t_L g2705 ( 
.A(n_2621),
.Y(n_2705)
);

INVxp67_ASAP7_75t_SL g2706 ( 
.A(n_2654),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2551),
.Y(n_2707)
);

INVx3_ASAP7_75t_L g2708 ( 
.A(n_2631),
.Y(n_2708)
);

INVx4_ASAP7_75t_L g2709 ( 
.A(n_2649),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2538),
.B(n_2483),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2600),
.B(n_2464),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2628),
.B(n_2291),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2507),
.Y(n_2713)
);

INVxp67_ASAP7_75t_L g2714 ( 
.A(n_2637),
.Y(n_2714)
);

OR2x2_ASAP7_75t_L g2715 ( 
.A(n_2539),
.B(n_2480),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2511),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2560),
.B(n_2465),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2567),
.Y(n_2718)
);

INVx4_ASAP7_75t_L g2719 ( 
.A(n_2649),
.Y(n_2719)
);

INVx4_ASAP7_75t_L g2720 ( 
.A(n_2655),
.Y(n_2720)
);

INVx3_ASAP7_75t_L g2721 ( 
.A(n_2655),
.Y(n_2721)
);

INVx3_ASAP7_75t_L g2722 ( 
.A(n_2632),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2574),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2491),
.B(n_2640),
.Y(n_2724)
);

OR2x2_ASAP7_75t_L g2725 ( 
.A(n_2650),
.B(n_2444),
.Y(n_2725)
);

INVx3_ASAP7_75t_L g2726 ( 
.A(n_2590),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2577),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2581),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2582),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2514),
.Y(n_2730)
);

OAI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_2599),
.A2(n_2601),
.B1(n_2586),
.B2(n_2589),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2583),
.Y(n_2732)
);

BUFx2_ASAP7_75t_L g2733 ( 
.A(n_2555),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2597),
.B(n_2473),
.Y(n_2734)
);

AND2x6_ASAP7_75t_L g2735 ( 
.A(n_2572),
.B(n_2482),
.Y(n_2735)
);

INVx4_ASAP7_75t_L g2736 ( 
.A(n_2570),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2522),
.Y(n_2737)
);

INVx1_ASAP7_75t_SL g2738 ( 
.A(n_2625),
.Y(n_2738)
);

OR2x6_ASAP7_75t_L g2739 ( 
.A(n_2610),
.B(n_2482),
.Y(n_2739)
);

INVx3_ASAP7_75t_L g2740 ( 
.A(n_2494),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2523),
.Y(n_2741)
);

INVxp33_ASAP7_75t_L g2742 ( 
.A(n_2626),
.Y(n_2742)
);

INVx4_ASAP7_75t_L g2743 ( 
.A(n_2501),
.Y(n_2743)
);

AND2x4_ASAP7_75t_L g2744 ( 
.A(n_2535),
.B(n_2285),
.Y(n_2744)
);

NOR2xp33_ASAP7_75t_L g2745 ( 
.A(n_2513),
.B(n_2436),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2596),
.A2(n_2265),
.B1(n_2271),
.B2(n_2257),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_L g2747 ( 
.A(n_2635),
.B(n_2277),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2556),
.B(n_2432),
.Y(n_2748)
);

AND2x4_ASAP7_75t_L g2749 ( 
.A(n_2549),
.B(n_2290),
.Y(n_2749)
);

INVx1_ASAP7_75t_SL g2750 ( 
.A(n_2564),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2527),
.Y(n_2751)
);

AO21x2_ASAP7_75t_L g2752 ( 
.A1(n_2633),
.A2(n_2317),
.B(n_2281),
.Y(n_2752)
);

AO22x2_ASAP7_75t_L g2753 ( 
.A1(n_2531),
.A2(n_2420),
.B1(n_2417),
.B2(n_2401),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_SL g2754 ( 
.A(n_2742),
.B(n_2609),
.Y(n_2754)
);

INVx2_ASAP7_75t_SL g2755 ( 
.A(n_2680),
.Y(n_2755)
);

NAND2xp33_ASAP7_75t_L g2756 ( 
.A(n_2669),
.B(n_2634),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2697),
.Y(n_2757)
);

AOI21xp5_ASAP7_75t_L g2758 ( 
.A1(n_2746),
.A2(n_2543),
.B(n_2651),
.Y(n_2758)
);

NAND3xp33_ASAP7_75t_L g2759 ( 
.A(n_2748),
.B(n_2545),
.C(n_2645),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2716),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2657),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2714),
.B(n_2573),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2730),
.Y(n_2763)
);

INVx2_ASAP7_75t_SL g2764 ( 
.A(n_2679),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2665),
.B(n_2518),
.Y(n_2765)
);

OR2x6_ASAP7_75t_L g2766 ( 
.A(n_2739),
.B(n_2659),
.Y(n_2766)
);

BUFx12f_ASAP7_75t_L g2767 ( 
.A(n_2696),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2687),
.B(n_2619),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2673),
.B(n_2614),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2668),
.B(n_2623),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2663),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2667),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2712),
.B(n_2575),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2670),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2676),
.B(n_2554),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2710),
.B(n_2563),
.Y(n_2776)
);

INVx2_ASAP7_75t_SL g2777 ( 
.A(n_2702),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2675),
.B(n_2558),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2741),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2677),
.B(n_2647),
.Y(n_2780)
);

INVx4_ASAP7_75t_L g2781 ( 
.A(n_2700),
.Y(n_2781)
);

AOI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2689),
.A2(n_2605),
.B1(n_2604),
.B2(n_2559),
.Y(n_2782)
);

INVx4_ASAP7_75t_L g2783 ( 
.A(n_2705),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2725),
.B(n_2296),
.Y(n_2784)
);

BUFx3_ASAP7_75t_L g2785 ( 
.A(n_2704),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2681),
.B(n_2529),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2685),
.B(n_2547),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2686),
.B(n_2644),
.Y(n_2788)
);

NOR2x2_ASAP7_75t_L g2789 ( 
.A(n_2733),
.B(n_2610),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2688),
.B(n_2636),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2691),
.B(n_2455),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_R g2792 ( 
.A(n_2660),
.B(n_2294),
.Y(n_2792)
);

CKINVDCx5p33_ASAP7_75t_R g2793 ( 
.A(n_2696),
.Y(n_2793)
);

INVx2_ASAP7_75t_SL g2794 ( 
.A(n_2692),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2682),
.B(n_2305),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2694),
.B(n_2638),
.Y(n_2796)
);

OR2x2_ASAP7_75t_L g2797 ( 
.A(n_2738),
.B(n_2602),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2695),
.B(n_2639),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_SL g2799 ( 
.A(n_2699),
.B(n_2542),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_L g2800 ( 
.A(n_2658),
.B(n_2552),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2656),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2707),
.B(n_2641),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2718),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2723),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2727),
.B(n_2642),
.Y(n_2805)
);

NOR2xp33_ASAP7_75t_L g2806 ( 
.A(n_2715),
.B(n_2611),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2728),
.B(n_2562),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2729),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2732),
.B(n_2565),
.Y(n_2809)
);

AND2x2_ASAP7_75t_SL g2810 ( 
.A(n_2736),
.B(n_2724),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2731),
.B(n_2569),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2737),
.A2(n_2504),
.B1(n_2557),
.B2(n_2383),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2662),
.B(n_2323),
.Y(n_2813)
);

BUFx6f_ASAP7_75t_L g2814 ( 
.A(n_2672),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2698),
.A2(n_2532),
.B1(n_2536),
.B2(n_2533),
.Y(n_2815)
);

AOI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_2747),
.A2(n_2540),
.B1(n_2553),
.B2(n_2550),
.Y(n_2816)
);

INVx2_ASAP7_75t_SL g2817 ( 
.A(n_2701),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2709),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2690),
.Y(n_2819)
);

O2A1O1Ixp5_ASAP7_75t_L g2820 ( 
.A1(n_2717),
.A2(n_2571),
.B(n_2520),
.C(n_2584),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2734),
.B(n_2576),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2671),
.Y(n_2822)
);

CKINVDCx5p33_ASAP7_75t_R g2823 ( 
.A(n_2693),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2745),
.B(n_2627),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2674),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2720),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2711),
.B(n_2525),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2683),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2684),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2713),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_SL g2831 ( 
.A(n_2664),
.B(n_2372),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2735),
.B(n_2593),
.Y(n_2832)
);

OR2x2_ASAP7_75t_L g2833 ( 
.A(n_2722),
.B(n_2299),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2735),
.B(n_2648),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2753),
.B(n_2618),
.Y(n_2835)
);

BUFx6f_ASAP7_75t_L g2836 ( 
.A(n_2719),
.Y(n_2836)
);

AND2x4_ASAP7_75t_L g2837 ( 
.A(n_2661),
.B(n_2328),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2761),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2762),
.B(n_2750),
.Y(n_2839)
);

BUFx6f_ASAP7_75t_L g2840 ( 
.A(n_2767),
.Y(n_2840)
);

O2A1O1Ixp33_ASAP7_75t_L g2841 ( 
.A1(n_2759),
.A2(n_2579),
.B(n_2643),
.C(n_2364),
.Y(n_2841)
);

HB1xp67_ASAP7_75t_L g2842 ( 
.A(n_2819),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2760),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2763),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2773),
.B(n_2776),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2771),
.Y(n_2846)
);

NOR2xp33_ASAP7_75t_L g2847 ( 
.A(n_2770),
.B(n_2726),
.Y(n_2847)
);

AND2x4_ASAP7_75t_L g2848 ( 
.A(n_2766),
.B(n_2721),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2779),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2772),
.Y(n_2850)
);

INVx1_ASAP7_75t_SL g2851 ( 
.A(n_2797),
.Y(n_2851)
);

OR2x6_ASAP7_75t_L g2852 ( 
.A(n_2766),
.B(n_2708),
.Y(n_2852)
);

AND2x4_ASAP7_75t_L g2853 ( 
.A(n_2785),
.B(n_2744),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2774),
.Y(n_2854)
);

NAND2x1p5_ASAP7_75t_L g2855 ( 
.A(n_2826),
.B(n_2743),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2784),
.B(n_2706),
.Y(n_2856)
);

CKINVDCx20_ASAP7_75t_R g2857 ( 
.A(n_2793),
.Y(n_2857)
);

AND3x2_ASAP7_75t_SL g2858 ( 
.A(n_2789),
.B(n_2751),
.C(n_2578),
.Y(n_2858)
);

NAND2x1p5_ASAP7_75t_L g2859 ( 
.A(n_2826),
.B(n_2749),
.Y(n_2859)
);

CKINVDCx5p33_ASAP7_75t_R g2860 ( 
.A(n_2757),
.Y(n_2860)
);

BUFx2_ASAP7_75t_L g2861 ( 
.A(n_2792),
.Y(n_2861)
);

BUFx6f_ASAP7_75t_L g2862 ( 
.A(n_2814),
.Y(n_2862)
);

OAI22xp5_ASAP7_75t_SL g2863 ( 
.A1(n_2782),
.A2(n_2666),
.B1(n_2678),
.B2(n_2240),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2801),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2822),
.Y(n_2865)
);

OR2x2_ASAP7_75t_SL g2866 ( 
.A(n_2834),
.B(n_2475),
.Y(n_2866)
);

AND2x4_ASAP7_75t_L g2867 ( 
.A(n_2764),
.B(n_2740),
.Y(n_2867)
);

BUFx4f_ASAP7_75t_L g2868 ( 
.A(n_2810),
.Y(n_2868)
);

BUFx12f_ASAP7_75t_L g2869 ( 
.A(n_2823),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2765),
.B(n_2329),
.Y(n_2870)
);

AND2x6_ASAP7_75t_L g2871 ( 
.A(n_2803),
.B(n_2804),
.Y(n_2871)
);

OR2x6_ASAP7_75t_SL g2872 ( 
.A(n_2832),
.B(n_1241),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2768),
.B(n_2693),
.Y(n_2873)
);

AOI22xp33_ASAP7_75t_L g2874 ( 
.A1(n_2812),
.A2(n_2580),
.B1(n_2585),
.B2(n_2561),
.Y(n_2874)
);

NAND2x1p5_ASAP7_75t_L g2875 ( 
.A(n_2814),
.B(n_2443),
.Y(n_2875)
);

AOI22xp5_ASAP7_75t_L g2876 ( 
.A1(n_2775),
.A2(n_2421),
.B1(n_2703),
.B2(n_2466),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_2755),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_L g2878 ( 
.A(n_2754),
.B(n_2474),
.Y(n_2878)
);

BUFx3_ASAP7_75t_L g2879 ( 
.A(n_2836),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2806),
.B(n_2778),
.Y(n_2880)
);

AOI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2795),
.A2(n_2269),
.B1(n_2274),
.B2(n_2264),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2825),
.Y(n_2882)
);

AND2x4_ASAP7_75t_L g2883 ( 
.A(n_2777),
.B(n_2282),
.Y(n_2883)
);

AOI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2827),
.A2(n_2289),
.B1(n_2292),
.B2(n_2286),
.Y(n_2884)
);

A2O1A1Ixp33_ASAP7_75t_L g2885 ( 
.A1(n_2758),
.A2(n_2615),
.B(n_2595),
.C(n_2312),
.Y(n_2885)
);

AOI211xp5_ASAP7_75t_L g2886 ( 
.A1(n_2756),
.A2(n_1507),
.B(n_1511),
.C(n_1505),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2808),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2796),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2829),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2780),
.B(n_2293),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2824),
.B(n_2298),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2798),
.Y(n_2892)
);

CKINVDCx20_ASAP7_75t_R g2893 ( 
.A(n_2781),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2828),
.Y(n_2894)
);

AOI211xp5_ASAP7_75t_L g2895 ( 
.A1(n_2835),
.A2(n_1528),
.B(n_1532),
.C(n_1522),
.Y(n_2895)
);

INVx5_ASAP7_75t_L g2896 ( 
.A(n_2836),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2830),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2783),
.Y(n_2898)
);

INVx4_ASAP7_75t_L g2899 ( 
.A(n_2837),
.Y(n_2899)
);

BUFx4f_ASAP7_75t_SL g2900 ( 
.A(n_2799),
.Y(n_2900)
);

AND2x4_ASAP7_75t_L g2901 ( 
.A(n_2794),
.B(n_2302),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2802),
.Y(n_2902)
);

BUFx6f_ASAP7_75t_SL g2903 ( 
.A(n_2840),
.Y(n_2903)
);

NAND3xp33_ASAP7_75t_L g2904 ( 
.A(n_2886),
.B(n_2800),
.C(n_2769),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2845),
.B(n_2821),
.Y(n_2905)
);

NOR2xp67_ASAP7_75t_L g2906 ( 
.A(n_2896),
.B(n_2817),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_SL g2907 ( 
.A(n_2880),
.B(n_2811),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2873),
.B(n_2818),
.Y(n_2908)
);

O2A1O1Ixp33_ASAP7_75t_L g2909 ( 
.A1(n_2841),
.A2(n_2895),
.B(n_2831),
.C(n_2870),
.Y(n_2909)
);

BUFx6f_ASAP7_75t_L g2910 ( 
.A(n_2862),
.Y(n_2910)
);

A2O1A1Ixp33_ASAP7_75t_L g2911 ( 
.A1(n_2878),
.A2(n_2791),
.B(n_2820),
.C(n_2787),
.Y(n_2911)
);

AOI22x1_ASAP7_75t_L g2912 ( 
.A1(n_2842),
.A2(n_1244),
.B1(n_1248),
.B2(n_1242),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2862),
.Y(n_2913)
);

AND2x4_ASAP7_75t_L g2914 ( 
.A(n_2861),
.B(n_2833),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2838),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2847),
.B(n_2805),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2885),
.A2(n_2752),
.B(n_2652),
.Y(n_2917)
);

INVx3_ASAP7_75t_L g2918 ( 
.A(n_2899),
.Y(n_2918)
);

INVx4_ASAP7_75t_L g2919 ( 
.A(n_2896),
.Y(n_2919)
);

OAI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2863),
.A2(n_2815),
.B1(n_2788),
.B2(n_2786),
.Y(n_2920)
);

BUFx3_ASAP7_75t_L g2921 ( 
.A(n_2893),
.Y(n_2921)
);

AOI21xp5_ASAP7_75t_L g2922 ( 
.A1(n_2888),
.A2(n_2790),
.B(n_2370),
.Y(n_2922)
);

O2A1O1Ixp5_ASAP7_75t_SL g2923 ( 
.A1(n_2846),
.A2(n_1534),
.B(n_1541),
.C(n_1537),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_R g2924 ( 
.A(n_2857),
.B(n_2475),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2850),
.Y(n_2925)
);

O2A1O1Ixp33_ASAP7_75t_L g2926 ( 
.A1(n_2890),
.A2(n_2813),
.B(n_1559),
.C(n_1588),
.Y(n_2926)
);

A2O1A1Ixp33_ASAP7_75t_L g2927 ( 
.A1(n_2876),
.A2(n_2809),
.B(n_2807),
.C(n_2313),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2868),
.B(n_2476),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2900),
.B(n_2379),
.Y(n_2929)
);

AOI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2892),
.A2(n_2255),
.B(n_2284),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2848),
.B(n_2379),
.Y(n_2931)
);

OA21x2_ASAP7_75t_L g2932 ( 
.A1(n_2854),
.A2(n_2568),
.B(n_2603),
.Y(n_2932)
);

INVx3_ASAP7_75t_L g2933 ( 
.A(n_2879),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2884),
.B(n_2839),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2887),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2894),
.Y(n_2936)
);

NOR2x1_ASAP7_75t_L g2937 ( 
.A(n_2891),
.B(n_1580),
.Y(n_2937)
);

A2O1A1Ixp33_ASAP7_75t_L g2938 ( 
.A1(n_2902),
.A2(n_2816),
.B(n_1592),
.C(n_1594),
.Y(n_2938)
);

INVx3_ASAP7_75t_L g2939 ( 
.A(n_2852),
.Y(n_2939)
);

O2A1O1Ixp33_ASAP7_75t_L g2940 ( 
.A1(n_2898),
.A2(n_1598),
.B(n_1608),
.C(n_1543),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2871),
.A2(n_2378),
.B(n_2377),
.Y(n_2941)
);

O2A1O1Ixp33_ASAP7_75t_L g2942 ( 
.A1(n_2855),
.A2(n_1616),
.B(n_1618),
.C(n_1611),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2897),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2843),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2856),
.B(n_1622),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2851),
.B(n_1625),
.Y(n_2946)
);

OAI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2866),
.A2(n_1636),
.B1(n_1642),
.B2(n_1629),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2871),
.B(n_1650),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2844),
.Y(n_2949)
);

BUFx2_ASAP7_75t_L g2950 ( 
.A(n_2871),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2849),
.B(n_1655),
.Y(n_2951)
);

NAND3xp33_ASAP7_75t_SL g2952 ( 
.A(n_2877),
.B(n_1251),
.C(n_1249),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2864),
.B(n_1662),
.Y(n_2953)
);

BUFx8_ASAP7_75t_SL g2954 ( 
.A(n_2860),
.Y(n_2954)
);

AOI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2865),
.A2(n_2608),
.B(n_2607),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2882),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2889),
.Y(n_2957)
);

O2A1O1Ixp33_ASAP7_75t_SL g2958 ( 
.A1(n_2881),
.A2(n_1679),
.B(n_1697),
.C(n_1676),
.Y(n_2958)
);

AOI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2875),
.A2(n_2613),
.B(n_1603),
.Y(n_2959)
);

OR2x2_ASAP7_75t_L g2960 ( 
.A(n_2859),
.B(n_2853),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2874),
.A2(n_1607),
.B(n_1585),
.Y(n_2961)
);

HB1xp67_ASAP7_75t_L g2962 ( 
.A(n_2883),
.Y(n_2962)
);

CKINVDCx11_ASAP7_75t_R g2963 ( 
.A(n_2872),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2943),
.Y(n_2964)
);

BUFx12f_ASAP7_75t_L g2965 ( 
.A(n_2963),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2916),
.B(n_2901),
.Y(n_2966)
);

INVx5_ASAP7_75t_L g2967 ( 
.A(n_2954),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2945),
.B(n_2915),
.Y(n_2968)
);

NAND2xp33_ASAP7_75t_L g2969 ( 
.A(n_2924),
.B(n_2840),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2905),
.B(n_2867),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2907),
.B(n_1699),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2936),
.Y(n_2972)
);

BUFx6f_ASAP7_75t_L g2973 ( 
.A(n_2910),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2925),
.B(n_1704),
.Y(n_2974)
);

OAI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_2904),
.A2(n_2869),
.B1(n_1718),
.B2(n_1720),
.Y(n_2975)
);

INVx4_ASAP7_75t_L g2976 ( 
.A(n_2910),
.Y(n_2976)
);

BUFx3_ASAP7_75t_L g2977 ( 
.A(n_2921),
.Y(n_2977)
);

BUFx2_ASAP7_75t_L g2978 ( 
.A(n_2950),
.Y(n_2978)
);

AOI22xp33_ASAP7_75t_L g2979 ( 
.A1(n_2920),
.A2(n_2592),
.B1(n_2616),
.B2(n_2591),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2935),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2944),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2917),
.A2(n_1722),
.B(n_1716),
.Y(n_2982)
);

INVx3_ASAP7_75t_L g2983 ( 
.A(n_2919),
.Y(n_2983)
);

BUFx6f_ASAP7_75t_L g2984 ( 
.A(n_2914),
.Y(n_2984)
);

O2A1O1Ixp33_ASAP7_75t_L g2985 ( 
.A1(n_2909),
.A2(n_1744),
.B(n_1745),
.C(n_1723),
.Y(n_2985)
);

INVx3_ASAP7_75t_L g2986 ( 
.A(n_2933),
.Y(n_2986)
);

BUFx2_ASAP7_75t_L g2987 ( 
.A(n_2962),
.Y(n_2987)
);

O2A1O1Ixp33_ASAP7_75t_SL g2988 ( 
.A1(n_2928),
.A2(n_1754),
.B(n_1761),
.C(n_1746),
.Y(n_2988)
);

AND2x4_ASAP7_75t_L g2989 ( 
.A(n_2939),
.B(n_2858),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_SL g2990 ( 
.A1(n_2948),
.A2(n_2947),
.B1(n_2912),
.B2(n_2946),
.Y(n_2990)
);

CKINVDCx5p33_ASAP7_75t_R g2991 ( 
.A(n_2903),
.Y(n_2991)
);

AOI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2937),
.A2(n_2624),
.B1(n_2617),
.B2(n_2307),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2934),
.B(n_1763),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_2960),
.B(n_2334),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2908),
.B(n_1770),
.Y(n_2995)
);

AOI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2911),
.A2(n_1799),
.B(n_1777),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2949),
.Y(n_2997)
);

OAI21xp5_ASAP7_75t_L g2998 ( 
.A1(n_2927),
.A2(n_1807),
.B(n_1801),
.Y(n_2998)
);

BUFx2_ASAP7_75t_L g2999 ( 
.A(n_2918),
.Y(n_2999)
);

OR2x2_ASAP7_75t_L g3000 ( 
.A(n_2956),
.B(n_1815),
.Y(n_3000)
);

BUFx2_ASAP7_75t_SL g3001 ( 
.A(n_2906),
.Y(n_3001)
);

BUFx3_ASAP7_75t_L g3002 ( 
.A(n_2913),
.Y(n_3002)
);

INVx4_ASAP7_75t_L g3003 ( 
.A(n_2929),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2938),
.A2(n_1835),
.B1(n_1844),
.B2(n_1834),
.Y(n_3004)
);

BUFx3_ASAP7_75t_L g3005 ( 
.A(n_2931),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2957),
.A2(n_2304),
.B1(n_1165),
.B2(n_1712),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2951),
.Y(n_3007)
);

AND2x4_ASAP7_75t_L g3008 ( 
.A(n_2953),
.B(n_2334),
.Y(n_3008)
);

INVx4_ASAP7_75t_L g3009 ( 
.A(n_2952),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2922),
.B(n_1845),
.Y(n_3010)
);

INVx3_ASAP7_75t_L g3011 ( 
.A(n_2932),
.Y(n_3011)
);

BUFx3_ASAP7_75t_L g3012 ( 
.A(n_2932),
.Y(n_3012)
);

BUFx3_ASAP7_75t_L g3013 ( 
.A(n_2942),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2926),
.B(n_1847),
.Y(n_3014)
);

AOI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2958),
.A2(n_1252),
.B1(n_1258),
.B2(n_1253),
.Y(n_3015)
);

NAND2x1p5_ASAP7_75t_L g3016 ( 
.A(n_2955),
.B(n_2339),
.Y(n_3016)
);

AOI221xp5_ASAP7_75t_L g3017 ( 
.A1(n_2940),
.A2(n_1856),
.B1(n_1260),
.B2(n_1272),
.C(n_1261),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_2959),
.Y(n_3018)
);

AOI21xp5_ASAP7_75t_L g3019 ( 
.A1(n_3010),
.A2(n_2982),
.B(n_2941),
.Y(n_3019)
);

AO31x2_ASAP7_75t_L g3020 ( 
.A1(n_2972),
.A2(n_2930),
.A3(n_2961),
.B(n_2923),
.Y(n_3020)
);

AOI221x1_ASAP7_75t_L g3021 ( 
.A1(n_2993),
.A2(n_1626),
.B1(n_1646),
.B2(n_1643),
.C(n_1641),
.Y(n_3021)
);

AOI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_3013),
.A2(n_1578),
.B1(n_1647),
.B2(n_1431),
.Y(n_3022)
);

AO31x2_ASAP7_75t_L g3023 ( 
.A1(n_2981),
.A2(n_1671),
.A3(n_1675),
.B(n_1657),
.Y(n_3023)
);

AND2x4_ASAP7_75t_L g3024 ( 
.A(n_2978),
.B(n_2339),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2980),
.Y(n_3025)
);

AND2x4_ASAP7_75t_L g3026 ( 
.A(n_2987),
.B(n_3005),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_3018),
.B(n_2476),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_2996),
.A2(n_1692),
.B(n_1682),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2985),
.A2(n_2998),
.B(n_3014),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2968),
.B(n_1578),
.Y(n_3030)
);

AND2x4_ASAP7_75t_L g3031 ( 
.A(n_2999),
.B(n_1702),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_3007),
.A2(n_1647),
.B1(n_1848),
.B2(n_1769),
.Y(n_3032)
);

OAI21xp33_ASAP7_75t_SL g3033 ( 
.A1(n_2976),
.A2(n_1748),
.B(n_1724),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2964),
.Y(n_3034)
);

AOI21xp5_ASAP7_75t_L g3035 ( 
.A1(n_2971),
.A2(n_1797),
.B(n_1786),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2984),
.B(n_1769),
.Y(n_3036)
);

OAI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_2975),
.A2(n_1830),
.B(n_1817),
.Y(n_3037)
);

AOI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2966),
.A2(n_1274),
.B(n_1259),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2995),
.B(n_2970),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2990),
.A2(n_1848),
.B1(n_1769),
.B2(n_1275),
.Y(n_3040)
);

O2A1O1Ixp33_ASAP7_75t_SL g3041 ( 
.A1(n_2983),
.A2(n_5),
.B(n_2),
.C(n_3),
.Y(n_3041)
);

AOI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_3016),
.A2(n_1280),
.B(n_1276),
.Y(n_3042)
);

OAI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_3015),
.A2(n_1301),
.B(n_1154),
.Y(n_3043)
);

CKINVDCx6p67_ASAP7_75t_R g3044 ( 
.A(n_2967),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2989),
.A2(n_1848),
.B1(n_1590),
.B2(n_1674),
.Y(n_3045)
);

A2O1A1Ixp33_ASAP7_75t_L g3046 ( 
.A1(n_3004),
.A2(n_1687),
.B(n_1700),
.C(n_1664),
.Y(n_3046)
);

OR2x2_ASAP7_75t_L g3047 ( 
.A(n_3000),
.B(n_2),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2988),
.A2(n_1286),
.B(n_1283),
.Y(n_3048)
);

OAI22xp5_ASAP7_75t_SL g3049 ( 
.A1(n_2965),
.A2(n_1298),
.B1(n_1299),
.B2(n_1291),
.Y(n_3049)
);

AO21x2_ASAP7_75t_L g3050 ( 
.A1(n_2974),
.A2(n_1826),
.B(n_1804),
.Y(n_3050)
);

A2O1A1Ixp33_ASAP7_75t_L g3051 ( 
.A1(n_3017),
.A2(n_1858),
.B(n_1302),
.C(n_1305),
.Y(n_3051)
);

AO31x2_ASAP7_75t_L g3052 ( 
.A1(n_2997),
.A2(n_3009),
.A3(n_3012),
.B(n_3011),
.Y(n_3052)
);

OAI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_3003),
.A2(n_2984),
.B1(n_3002),
.B2(n_2977),
.Y(n_3053)
);

AO31x2_ASAP7_75t_L g3054 ( 
.A1(n_3001),
.A2(n_2479),
.A3(n_1306),
.B(n_1312),
.Y(n_3054)
);

CKINVDCx5p33_ASAP7_75t_R g3055 ( 
.A(n_2991),
.Y(n_3055)
);

NAND2xp33_ASAP7_75t_L g3056 ( 
.A(n_2967),
.B(n_1303),
.Y(n_3056)
);

O2A1O1Ixp33_ASAP7_75t_SL g3057 ( 
.A1(n_2986),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_3057)
);

A2O1A1Ixp33_ASAP7_75t_L g3058 ( 
.A1(n_2969),
.A2(n_1317),
.B(n_1321),
.C(n_1320),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2979),
.A2(n_1326),
.B(n_1324),
.Y(n_3059)
);

INVx4_ASAP7_75t_L g3060 ( 
.A(n_2973),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_3008),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2973),
.Y(n_3062)
);

NOR2xp33_ASAP7_75t_L g3063 ( 
.A(n_2994),
.B(n_6),
.Y(n_3063)
);

BUFx8_ASAP7_75t_L g3064 ( 
.A(n_2992),
.Y(n_3064)
);

O2A1O1Ixp33_ASAP7_75t_SL g3065 ( 
.A1(n_3006),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_3065)
);

OR2x6_ASAP7_75t_L g3066 ( 
.A(n_3026),
.B(n_3027),
.Y(n_3066)
);

OAI22xp33_ASAP7_75t_L g3067 ( 
.A1(n_3029),
.A2(n_1328),
.B1(n_1330),
.B2(n_1329),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_3025),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_3044),
.B(n_8),
.Y(n_3069)
);

CKINVDCx5p33_ASAP7_75t_R g3070 ( 
.A(n_3055),
.Y(n_3070)
);

CKINVDCx20_ASAP7_75t_R g3071 ( 
.A(n_3062),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_3034),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3052),
.Y(n_3073)
);

INVx2_ASAP7_75t_SL g3074 ( 
.A(n_3024),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_3052),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_3040),
.A2(n_1524),
.B1(n_1635),
.B2(n_1277),
.Y(n_3076)
);

OAI221xp5_ASAP7_75t_L g3077 ( 
.A1(n_3043),
.A2(n_1410),
.B1(n_1422),
.B2(n_1393),
.C(n_1378),
.Y(n_3077)
);

AOI221xp5_ASAP7_75t_L g3078 ( 
.A1(n_3035),
.A2(n_1334),
.B1(n_1339),
.B2(n_1338),
.C(n_1333),
.Y(n_3078)
);

A2O1A1Ixp33_ASAP7_75t_L g3079 ( 
.A1(n_3033),
.A2(n_1361),
.B(n_1374),
.C(n_1348),
.Y(n_3079)
);

AND2x4_ASAP7_75t_L g3080 ( 
.A(n_3061),
.B(n_3060),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_3030),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_3036),
.Y(n_3082)
);

AOI22xp33_ASAP7_75t_L g3083 ( 
.A1(n_3050),
.A2(n_3064),
.B1(n_3037),
.B2(n_3019),
.Y(n_3083)
);

AOI22xp33_ASAP7_75t_L g3084 ( 
.A1(n_3022),
.A2(n_1524),
.B1(n_1635),
.B2(n_1277),
.Y(n_3084)
);

OAI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_3045),
.A2(n_1343),
.B1(n_1347),
.B2(n_1345),
.Y(n_3085)
);

AOI22xp33_ASAP7_75t_L g3086 ( 
.A1(n_3038),
.A2(n_1524),
.B1(n_1635),
.B2(n_1277),
.Y(n_3086)
);

NOR2x1_ASAP7_75t_L g3087 ( 
.A(n_3053),
.B(n_2380),
.Y(n_3087)
);

INVx4_ASAP7_75t_L g3088 ( 
.A(n_3031),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_3039),
.B(n_11),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_L g3090 ( 
.A1(n_3028),
.A2(n_1810),
.B1(n_1351),
.B2(n_1354),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_3063),
.B(n_11),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_3047),
.B(n_12),
.Y(n_3092)
);

OAI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_3051),
.A2(n_1357),
.B1(n_1362),
.B2(n_1349),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3023),
.Y(n_3094)
);

AOI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_3065),
.A2(n_1365),
.B(n_1363),
.Y(n_3095)
);

AOI22xp33_ASAP7_75t_L g3096 ( 
.A1(n_3032),
.A2(n_1810),
.B1(n_1369),
.B2(n_1373),
.Y(n_3096)
);

OAI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_3058),
.A2(n_3049),
.B1(n_3046),
.B2(n_3042),
.Y(n_3097)
);

CKINVDCx11_ASAP7_75t_R g3098 ( 
.A(n_3056),
.Y(n_3098)
);

INVx4_ASAP7_75t_L g3099 ( 
.A(n_3041),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_3023),
.Y(n_3100)
);

AND2x4_ASAP7_75t_L g3101 ( 
.A(n_3054),
.B(n_1810),
.Y(n_3101)
);

BUFx6f_ASAP7_75t_L g3102 ( 
.A(n_3057),
.Y(n_3102)
);

AOI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_3059),
.A2(n_1381),
.B1(n_1385),
.B2(n_1368),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_3054),
.B(n_12),
.Y(n_3104)
);

INVx1_ASAP7_75t_SL g3105 ( 
.A(n_3048),
.Y(n_3105)
);

OAI22xp5_ASAP7_75t_L g3106 ( 
.A1(n_3021),
.A2(n_1387),
.B1(n_1389),
.B2(n_1386),
.Y(n_3106)
);

OR2x6_ASAP7_75t_L g3107 ( 
.A(n_3020),
.B(n_2380),
.Y(n_3107)
);

AND2x4_ASAP7_75t_L g3108 ( 
.A(n_3020),
.B(n_13),
.Y(n_3108)
);

OAI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_3029),
.A2(n_1850),
.B1(n_1851),
.B2(n_1843),
.Y(n_3109)
);

OAI221xp5_ASAP7_75t_L g3110 ( 
.A1(n_3040),
.A2(n_1477),
.B1(n_1495),
.B2(n_1428),
.C(n_1409),
.Y(n_3110)
);

OAI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_3029),
.A2(n_1397),
.B(n_1392),
.Y(n_3111)
);

INVx1_ASAP7_75t_SL g3112 ( 
.A(n_3026),
.Y(n_3112)
);

NOR2xp33_ASAP7_75t_L g3113 ( 
.A(n_3044),
.B(n_14),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3025),
.Y(n_3114)
);

AOI22xp33_ASAP7_75t_L g3115 ( 
.A1(n_3029),
.A2(n_1400),
.B1(n_1403),
.B2(n_1399),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_L g3116 ( 
.A1(n_3029),
.A2(n_1412),
.B1(n_1413),
.B2(n_1407),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_3025),
.Y(n_3117)
);

INVx2_ASAP7_75t_SL g3118 ( 
.A(n_3026),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_3026),
.Y(n_3119)
);

OAI22xp5_ASAP7_75t_L g3120 ( 
.A1(n_3029),
.A2(n_1420),
.B1(n_1421),
.B2(n_1418),
.Y(n_3120)
);

O2A1O1Ixp33_ASAP7_75t_SL g3121 ( 
.A1(n_3053),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_3034),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_3034),
.Y(n_3123)
);

INVxp67_ASAP7_75t_L g3124 ( 
.A(n_3119),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3068),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_3114),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_3122),
.Y(n_3127)
);

BUFx2_ASAP7_75t_L g3128 ( 
.A(n_3066),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_3123),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_3117),
.Y(n_3130)
);

OA21x2_ASAP7_75t_L g3131 ( 
.A1(n_3073),
.A2(n_1435),
.B(n_1432),
.Y(n_3131)
);

OAI22xp5_ASAP7_75t_L g3132 ( 
.A1(n_3099),
.A2(n_1446),
.B1(n_1449),
.B2(n_1440),
.Y(n_3132)
);

OAI21x1_ASAP7_75t_L g3133 ( 
.A1(n_3075),
.A2(n_3087),
.B(n_3100),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_3081),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_3072),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3094),
.Y(n_3136)
);

OAI221xp5_ASAP7_75t_L g3137 ( 
.A1(n_3111),
.A2(n_1461),
.B1(n_1462),
.B2(n_1455),
.C(n_1452),
.Y(n_3137)
);

HB1xp67_ASAP7_75t_SL g3138 ( 
.A(n_3070),
.Y(n_3138)
);

BUFx2_ASAP7_75t_L g3139 ( 
.A(n_3066),
.Y(n_3139)
);

AOI22xp5_ASAP7_75t_L g3140 ( 
.A1(n_3120),
.A2(n_1468),
.B1(n_1470),
.B2(n_1464),
.Y(n_3140)
);

INVx1_ASAP7_75t_SL g3141 ( 
.A(n_3098),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3082),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3108),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3080),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3112),
.Y(n_3145)
);

OR2x2_ASAP7_75t_L g3146 ( 
.A(n_3118),
.B(n_15),
.Y(n_3146)
);

AND2x4_ASAP7_75t_L g3147 ( 
.A(n_3074),
.B(n_16),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_3089),
.B(n_1476),
.Y(n_3148)
);

HB1xp67_ASAP7_75t_L g3149 ( 
.A(n_3107),
.Y(n_3149)
);

AO21x2_ASAP7_75t_L g3150 ( 
.A1(n_3092),
.A2(n_2238),
.B(n_1488),
.Y(n_3150)
);

BUFx6f_ASAP7_75t_L g3151 ( 
.A(n_3088),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3107),
.Y(n_3152)
);

AOI22xp33_ASAP7_75t_L g3153 ( 
.A1(n_3101),
.A2(n_1852),
.B1(n_1492),
.B2(n_1497),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_3104),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_3071),
.B(n_17),
.Y(n_3155)
);

HB1xp67_ASAP7_75t_L g3156 ( 
.A(n_3091),
.Y(n_3156)
);

BUFx2_ASAP7_75t_L g3157 ( 
.A(n_3069),
.Y(n_3157)
);

OAI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_3115),
.A2(n_1500),
.B1(n_1501),
.B2(n_1482),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_3083),
.B(n_2386),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_3113),
.B(n_18),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_3105),
.Y(n_3161)
);

OAI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_3067),
.A2(n_1506),
.B(n_1504),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_3102),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3102),
.Y(n_3164)
);

NOR2x1_ASAP7_75t_L g3165 ( 
.A(n_3109),
.B(n_2386),
.Y(n_3165)
);

HB1xp67_ASAP7_75t_L g3166 ( 
.A(n_3097),
.Y(n_3166)
);

BUFx2_ASAP7_75t_L g3167 ( 
.A(n_3079),
.Y(n_3167)
);

OA21x2_ASAP7_75t_L g3168 ( 
.A1(n_3116),
.A2(n_1509),
.B(n_1508),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3121),
.Y(n_3169)
);

INVxp67_ASAP7_75t_L g3170 ( 
.A(n_3110),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_3086),
.B(n_1510),
.Y(n_3171)
);

INVx1_ASAP7_75t_SL g3172 ( 
.A(n_3103),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3106),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3076),
.B(n_3084),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3095),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_3077),
.Y(n_3176)
);

OA21x2_ASAP7_75t_L g3177 ( 
.A1(n_3096),
.A2(n_1516),
.B(n_1514),
.Y(n_3177)
);

OAI21x1_ASAP7_75t_L g3178 ( 
.A1(n_3085),
.A2(n_18),
.B(n_19),
.Y(n_3178)
);

OAI21x1_ASAP7_75t_L g3179 ( 
.A1(n_3090),
.A2(n_19),
.B(n_20),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_3078),
.B(n_20),
.Y(n_3180)
);

OAI221xp5_ASAP7_75t_L g3181 ( 
.A1(n_3166),
.A2(n_3093),
.B1(n_1523),
.B2(n_1525),
.C(n_1520),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_3133),
.Y(n_3182)
);

INVx3_ASAP7_75t_L g3183 ( 
.A(n_3151),
.Y(n_3183)
);

AOI211xp5_ASAP7_75t_L g3184 ( 
.A1(n_3132),
.A2(n_3169),
.B(n_3167),
.C(n_3173),
.Y(n_3184)
);

AOI21xp33_ASAP7_75t_L g3185 ( 
.A1(n_3152),
.A2(n_1527),
.B(n_1517),
.Y(n_3185)
);

AOI22xp33_ASAP7_75t_L g3186 ( 
.A1(n_3154),
.A2(n_1531),
.B1(n_1535),
.B2(n_1529),
.Y(n_3186)
);

AOI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_3161),
.A2(n_1542),
.B1(n_1544),
.B2(n_1538),
.Y(n_3187)
);

OAI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_3128),
.A2(n_3139),
.B1(n_3157),
.B2(n_3124),
.Y(n_3188)
);

OAI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_3156),
.A2(n_1556),
.B1(n_1558),
.B2(n_1555),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3144),
.B(n_21),
.Y(n_3190)
);

AOI222xp33_ASAP7_75t_L g3191 ( 
.A1(n_3176),
.A2(n_1573),
.B1(n_1567),
.B2(n_1577),
.C1(n_1572),
.C2(n_1563),
.Y(n_3191)
);

OAI221xp5_ASAP7_75t_L g3192 ( 
.A1(n_3170),
.A2(n_1582),
.B1(n_1583),
.B2(n_1581),
.C(n_1579),
.Y(n_3192)
);

INVx3_ASAP7_75t_L g3193 ( 
.A(n_3151),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3136),
.Y(n_3194)
);

HB1xp67_ASAP7_75t_L g3195 ( 
.A(n_3125),
.Y(n_3195)
);

BUFx8_ASAP7_75t_SL g3196 ( 
.A(n_3147),
.Y(n_3196)
);

A2O1A1Ixp33_ASAP7_75t_L g3197 ( 
.A1(n_3165),
.A2(n_1589),
.B(n_1595),
.C(n_1587),
.Y(n_3197)
);

OR2x2_ASAP7_75t_L g3198 ( 
.A(n_3135),
.B(n_21),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_3127),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_3143),
.A2(n_1602),
.B1(n_1606),
.B2(n_1596),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_3141),
.Y(n_3201)
);

OAI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_3146),
.A2(n_1637),
.B1(n_1653),
.B2(n_1621),
.Y(n_3202)
);

AOI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_3175),
.A2(n_1615),
.B1(n_1617),
.B2(n_1612),
.Y(n_3203)
);

AO31x2_ASAP7_75t_L g3204 ( 
.A1(n_3163),
.A2(n_30),
.A3(n_39),
.B(n_22),
.Y(n_3204)
);

AOI22xp33_ASAP7_75t_L g3205 ( 
.A1(n_3131),
.A2(n_1620),
.B1(n_1628),
.B2(n_1619),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_SL g3206 ( 
.A1(n_3160),
.A2(n_3150),
.B1(n_3172),
.B2(n_3168),
.Y(n_3206)
);

OAI221xp5_ASAP7_75t_L g3207 ( 
.A1(n_3153),
.A2(n_1634),
.B1(n_1638),
.B2(n_1632),
.C(n_1631),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3126),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_L g3209 ( 
.A1(n_3159),
.A2(n_1640),
.B1(n_1644),
.B2(n_1639),
.Y(n_3209)
);

AOI22xp33_ASAP7_75t_L g3210 ( 
.A1(n_3177),
.A2(n_1648),
.B1(n_1651),
.B2(n_1645),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3130),
.Y(n_3211)
);

OA21x2_ASAP7_75t_L g3212 ( 
.A1(n_3129),
.A2(n_1656),
.B(n_1654),
.Y(n_3212)
);

OR2x2_ASAP7_75t_L g3213 ( 
.A(n_3145),
.B(n_22),
.Y(n_3213)
);

OAI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_3164),
.A2(n_1698),
.B1(n_1739),
.B2(n_1681),
.Y(n_3214)
);

A2O1A1Ixp33_ASAP7_75t_L g3215 ( 
.A1(n_3155),
.A2(n_1663),
.B(n_1667),
.C(n_1661),
.Y(n_3215)
);

AOI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_3180),
.A2(n_1670),
.B1(n_1672),
.B2(n_1668),
.Y(n_3216)
);

AOI211xp5_ASAP7_75t_L g3217 ( 
.A1(n_3137),
.A2(n_1684),
.B(n_1685),
.C(n_1673),
.Y(n_3217)
);

OAI22xp33_ASAP7_75t_L g3218 ( 
.A1(n_3149),
.A2(n_1719),
.B1(n_1743),
.B2(n_1705),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3142),
.B(n_23),
.Y(n_3219)
);

BUFx3_ASAP7_75t_L g3220 ( 
.A(n_3148),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_3138),
.B(n_23),
.Y(n_3221)
);

OAI22xp33_ASAP7_75t_L g3222 ( 
.A1(n_3140),
.A2(n_1736),
.B1(n_1751),
.B2(n_1707),
.Y(n_3222)
);

A2O1A1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_3178),
.A2(n_1694),
.B(n_1695),
.C(n_1691),
.Y(n_3223)
);

OR2x2_ASAP7_75t_L g3224 ( 
.A(n_3134),
.B(n_24),
.Y(n_3224)
);

AND2x4_ASAP7_75t_L g3225 ( 
.A(n_3179),
.B(n_24),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_3171),
.A2(n_1708),
.B(n_1703),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3174),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_3162),
.Y(n_3228)
);

AOI221xp5_ASAP7_75t_L g3229 ( 
.A1(n_3158),
.A2(n_1717),
.B1(n_1721),
.B2(n_1714),
.C(n_1711),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3166),
.A2(n_1727),
.B1(n_1730),
.B2(n_1725),
.Y(n_3230)
);

AOI22xp33_ASAP7_75t_L g3231 ( 
.A1(n_3166),
.A2(n_1738),
.B1(n_1742),
.B2(n_1734),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_3156),
.B(n_25),
.Y(n_3232)
);

OAI22xp33_ASAP7_75t_L g3233 ( 
.A1(n_3166),
.A2(n_1767),
.B1(n_1782),
.B2(n_1755),
.Y(n_3233)
);

INVx2_ASAP7_75t_SL g3234 ( 
.A(n_3151),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_3156),
.B(n_25),
.Y(n_3235)
);

AOI222xp33_ASAP7_75t_L g3236 ( 
.A1(n_3167),
.A2(n_1752),
.B1(n_1749),
.B2(n_1758),
.C1(n_1750),
.C2(n_1747),
.Y(n_3236)
);

AOI22xp33_ASAP7_75t_SL g3237 ( 
.A1(n_3166),
.A2(n_1762),
.B1(n_1764),
.B2(n_1759),
.Y(n_3237)
);

OAI22xp33_ASAP7_75t_L g3238 ( 
.A1(n_3166),
.A2(n_1792),
.B1(n_1818),
.B2(n_1773),
.Y(n_3238)
);

AO21x2_ASAP7_75t_L g3239 ( 
.A1(n_3161),
.A2(n_26),
.B(n_27),
.Y(n_3239)
);

AOI221xp5_ASAP7_75t_L g3240 ( 
.A1(n_3166),
.A2(n_1768),
.B1(n_1771),
.B2(n_1766),
.C(n_1765),
.Y(n_3240)
);

NAND3xp33_ASAP7_75t_L g3241 ( 
.A(n_3166),
.B(n_1778),
.C(n_1776),
.Y(n_3241)
);

AOI221xp5_ASAP7_75t_L g3242 ( 
.A1(n_3166),
.A2(n_1785),
.B1(n_1794),
.B2(n_1783),
.C(n_1780),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3161),
.B(n_1798),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3161),
.B(n_1808),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3136),
.Y(n_3245)
);

AOI21x1_ASAP7_75t_L g3246 ( 
.A1(n_3166),
.A2(n_1823),
.B(n_1813),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3136),
.Y(n_3247)
);

AOI22xp5_ASAP7_75t_SL g3248 ( 
.A1(n_3166),
.A2(n_1825),
.B1(n_1831),
.B2(n_1824),
.Y(n_3248)
);

AOI22xp5_ASAP7_75t_L g3249 ( 
.A1(n_3166),
.A2(n_1838),
.B1(n_1839),
.B2(n_1836),
.Y(n_3249)
);

AOI22xp33_ASAP7_75t_L g3250 ( 
.A1(n_3166),
.A2(n_1842),
.B1(n_1853),
.B2(n_1841),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3136),
.Y(n_3251)
);

OAI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_3166),
.A2(n_1860),
.B1(n_1861),
.B2(n_1855),
.Y(n_3252)
);

AOI22xp33_ASAP7_75t_SL g3253 ( 
.A1(n_3166),
.A2(n_1862),
.B1(n_2408),
.B2(n_1167),
.Y(n_3253)
);

OAI22xp5_ASAP7_75t_L g3254 ( 
.A1(n_3166),
.A2(n_2408),
.B1(n_1822),
.B2(n_1829),
.Y(n_3254)
);

AOI22xp33_ASAP7_75t_L g3255 ( 
.A1(n_3166),
.A2(n_1172),
.B1(n_1175),
.B2(n_1161),
.Y(n_3255)
);

AOI22xp33_ASAP7_75t_L g3256 ( 
.A1(n_3166),
.A2(n_1178),
.B1(n_1187),
.B2(n_1177),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3136),
.Y(n_3257)
);

BUFx5_ASAP7_75t_L g3258 ( 
.A(n_3163),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_3166),
.A2(n_1196),
.B(n_1188),
.Y(n_3259)
);

OR2x2_ASAP7_75t_L g3260 ( 
.A(n_3161),
.B(n_26),
.Y(n_3260)
);

A2O1A1Ixp33_ASAP7_75t_L g3261 ( 
.A1(n_3166),
.A2(n_1204),
.B(n_1209),
.C(n_1197),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3136),
.Y(n_3262)
);

OAI22xp5_ASAP7_75t_SL g3263 ( 
.A1(n_3166),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_3263)
);

BUFx5_ASAP7_75t_L g3264 ( 
.A(n_3163),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3136),
.Y(n_3265)
);

OAI22xp5_ASAP7_75t_L g3266 ( 
.A1(n_3166),
.A2(n_1816),
.B1(n_1820),
.B2(n_1811),
.Y(n_3266)
);

AOI22xp33_ASAP7_75t_L g3267 ( 
.A1(n_3166),
.A2(n_1220),
.B1(n_1226),
.B2(n_1213),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3136),
.Y(n_3268)
);

BUFx6f_ASAP7_75t_L g3269 ( 
.A(n_3151),
.Y(n_3269)
);

AOI22xp33_ASAP7_75t_L g3270 ( 
.A1(n_3166),
.A2(n_1247),
.B1(n_1254),
.B2(n_1239),
.Y(n_3270)
);

AO21x2_ASAP7_75t_L g3271 ( 
.A1(n_3161),
.A2(n_29),
.B(n_30),
.Y(n_3271)
);

OAI211xp5_ASAP7_75t_L g3272 ( 
.A1(n_3169),
.A2(n_34),
.B(n_31),
.C(n_32),
.Y(n_3272)
);

OAI22xp33_ASAP7_75t_L g3273 ( 
.A1(n_3166),
.A2(n_1740),
.B1(n_1741),
.B2(n_1735),
.Y(n_3273)
);

CKINVDCx5p33_ASAP7_75t_R g3274 ( 
.A(n_3138),
.Y(n_3274)
);

BUFx3_ASAP7_75t_L g3275 ( 
.A(n_3141),
.Y(n_3275)
);

AOI22xp33_ASAP7_75t_SL g3276 ( 
.A1(n_3166),
.A2(n_1262),
.B1(n_1267),
.B2(n_1256),
.Y(n_3276)
);

OAI211xp5_ASAP7_75t_L g3277 ( 
.A1(n_3169),
.A2(n_34),
.B(n_31),
.C(n_32),
.Y(n_3277)
);

AOI222xp33_ASAP7_75t_L g3278 ( 
.A1(n_3167),
.A2(n_1319),
.B1(n_1307),
.B2(n_1327),
.C1(n_1318),
.C2(n_1292),
.Y(n_3278)
);

AOI221xp5_ASAP7_75t_L g3279 ( 
.A1(n_3166),
.A2(n_1340),
.B1(n_1355),
.B2(n_1332),
.C(n_1331),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3136),
.Y(n_3280)
);

AOI22xp5_ASAP7_75t_L g3281 ( 
.A1(n_3166),
.A2(n_1359),
.B1(n_1366),
.B2(n_1358),
.Y(n_3281)
);

AOI221xp5_ASAP7_75t_L g3282 ( 
.A1(n_3166),
.A2(n_1377),
.B1(n_1380),
.B2(n_1376),
.C(n_1375),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_3156),
.B(n_35),
.Y(n_3283)
);

AOI22xp33_ASAP7_75t_L g3284 ( 
.A1(n_3166),
.A2(n_1411),
.B1(n_1415),
.B2(n_1398),
.Y(n_3284)
);

OAI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3166),
.A2(n_1706),
.B1(n_1713),
.B2(n_1701),
.Y(n_3285)
);

AOI322xp5_ASAP7_75t_L g3286 ( 
.A1(n_3166),
.A2(n_41),
.A3(n_39),
.B1(n_37),
.B2(n_35),
.C1(n_36),
.C2(n_38),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_3156),
.B(n_41),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_3166),
.A2(n_1436),
.B(n_1430),
.Y(n_3288)
);

HB1xp67_ASAP7_75t_L g3289 ( 
.A(n_3161),
.Y(n_3289)
);

AOI22xp33_ASAP7_75t_L g3290 ( 
.A1(n_3166),
.A2(n_1439),
.B1(n_1444),
.B2(n_1438),
.Y(n_3290)
);

OAI211xp5_ASAP7_75t_L g3291 ( 
.A1(n_3169),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_3182),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3289),
.B(n_3195),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3239),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_3188),
.B(n_42),
.Y(n_3295)
);

OR2x2_ASAP7_75t_L g3296 ( 
.A(n_3208),
.B(n_43),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_3183),
.B(n_44),
.Y(n_3297)
);

AND2x4_ASAP7_75t_L g3298 ( 
.A(n_3275),
.B(n_45),
.Y(n_3298)
);

OR2x2_ASAP7_75t_L g3299 ( 
.A(n_3211),
.B(n_45),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3194),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3193),
.B(n_46),
.Y(n_3301)
);

BUFx3_ASAP7_75t_L g3302 ( 
.A(n_3196),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_3206),
.A2(n_1448),
.B1(n_1450),
.B2(n_1445),
.Y(n_3303)
);

INVx2_ASAP7_75t_SL g3304 ( 
.A(n_3201),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3271),
.Y(n_3305)
);

BUFx6f_ASAP7_75t_L g3306 ( 
.A(n_3269),
.Y(n_3306)
);

AND2x4_ASAP7_75t_L g3307 ( 
.A(n_3234),
.B(n_47),
.Y(n_3307)
);

HB1xp67_ASAP7_75t_L g3308 ( 
.A(n_3245),
.Y(n_3308)
);

NOR2xp67_ASAP7_75t_L g3309 ( 
.A(n_3274),
.B(n_47),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3247),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3199),
.Y(n_3311)
);

INVx3_ASAP7_75t_L g3312 ( 
.A(n_3269),
.Y(n_3312)
);

AND2x2_ASAP7_75t_L g3313 ( 
.A(n_3258),
.B(n_48),
.Y(n_3313)
);

CKINVDCx5p33_ASAP7_75t_R g3314 ( 
.A(n_3220),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3224),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_3204),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_3258),
.B(n_48),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3251),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3258),
.B(n_49),
.Y(n_3319)
);

BUFx4f_ASAP7_75t_L g3320 ( 
.A(n_3212),
.Y(n_3320)
);

OAI221xp5_ASAP7_75t_L g3321 ( 
.A1(n_3216),
.A2(n_1478),
.B1(n_1479),
.B2(n_1474),
.C(n_1460),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3204),
.Y(n_3322)
);

AOI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_3228),
.A2(n_3263),
.B1(n_3252),
.B2(n_3230),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3258),
.B(n_49),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_3257),
.B(n_50),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3264),
.Y(n_3326)
);

AOI221xp5_ASAP7_75t_L g3327 ( 
.A1(n_3233),
.A2(n_1496),
.B1(n_1498),
.B2(n_1491),
.C(n_1487),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3264),
.B(n_51),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3264),
.B(n_51),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3264),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3262),
.Y(n_3331)
);

INVx2_ASAP7_75t_SL g3332 ( 
.A(n_3232),
.Y(n_3332)
);

INVx3_ASAP7_75t_L g3333 ( 
.A(n_3198),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3265),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3235),
.B(n_53),
.Y(n_3335)
);

INVx3_ASAP7_75t_L g3336 ( 
.A(n_3213),
.Y(n_3336)
);

AOI22xp33_ASAP7_75t_L g3337 ( 
.A1(n_3227),
.A2(n_1518),
.B1(n_1540),
.B2(n_1515),
.Y(n_3337)
);

HB1xp67_ASAP7_75t_L g3338 ( 
.A(n_3268),
.Y(n_3338)
);

AOI21x1_ASAP7_75t_L g3339 ( 
.A1(n_3243),
.A2(n_54),
.B(n_57),
.Y(n_3339)
);

OR2x2_ASAP7_75t_L g3340 ( 
.A(n_3280),
.B(n_3260),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3283),
.B(n_58),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_3287),
.B(n_58),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3219),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_3190),
.B(n_59),
.Y(n_3344)
);

OR2x2_ASAP7_75t_L g3345 ( 
.A(n_3244),
.B(n_60),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_3225),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3200),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3221),
.B(n_60),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3184),
.B(n_61),
.Y(n_3349)
);

AND2x4_ASAP7_75t_L g3350 ( 
.A(n_3241),
.B(n_61),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_3249),
.B(n_62),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_3246),
.Y(n_3352)
);

OR2x2_ASAP7_75t_L g3353 ( 
.A(n_3189),
.B(n_62),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3187),
.Y(n_3354)
);

BUFx2_ASAP7_75t_L g3355 ( 
.A(n_3218),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_3281),
.Y(n_3356)
);

OAI22xp5_ASAP7_75t_L g3357 ( 
.A1(n_3231),
.A2(n_1548),
.B1(n_1557),
.B2(n_1552),
.Y(n_3357)
);

HB1xp67_ASAP7_75t_L g3358 ( 
.A(n_3254),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3203),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3186),
.Y(n_3360)
);

BUFx3_ASAP7_75t_L g3361 ( 
.A(n_3181),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3266),
.Y(n_3362)
);

BUFx3_ASAP7_75t_L g3363 ( 
.A(n_3192),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3250),
.B(n_63),
.Y(n_3364)
);

HB1xp67_ASAP7_75t_L g3365 ( 
.A(n_3285),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3248),
.B(n_63),
.Y(n_3366)
);

HB1xp67_ASAP7_75t_L g3367 ( 
.A(n_3185),
.Y(n_3367)
);

AO21x2_ASAP7_75t_L g3368 ( 
.A1(n_3259),
.A2(n_64),
.B(n_66),
.Y(n_3368)
);

INVx1_ASAP7_75t_SL g3369 ( 
.A(n_3253),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3207),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3238),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3273),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3237),
.B(n_66),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3255),
.B(n_67),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3272),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3277),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3256),
.B(n_68),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3291),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3267),
.B(n_68),
.Y(n_3379)
);

INVx3_ASAP7_75t_L g3380 ( 
.A(n_3202),
.Y(n_3380)
);

HB1xp67_ASAP7_75t_L g3381 ( 
.A(n_3288),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_3270),
.B(n_69),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3284),
.B(n_69),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3240),
.B(n_70),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3290),
.B(n_3215),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3214),
.Y(n_3386)
);

HB1xp67_ASAP7_75t_L g3387 ( 
.A(n_3242),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3276),
.B(n_70),
.Y(n_3388)
);

HB1xp67_ASAP7_75t_L g3389 ( 
.A(n_3223),
.Y(n_3389)
);

INVx3_ASAP7_75t_L g3390 ( 
.A(n_3286),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3197),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3205),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_3261),
.B(n_71),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3236),
.B(n_72),
.Y(n_3394)
);

AND2x4_ASAP7_75t_L g3395 ( 
.A(n_3209),
.B(n_73),
.Y(n_3395)
);

AND2x4_ASAP7_75t_SL g3396 ( 
.A(n_3210),
.B(n_73),
.Y(n_3396)
);

BUFx2_ASAP7_75t_L g3397 ( 
.A(n_3279),
.Y(n_3397)
);

OR2x2_ASAP7_75t_L g3398 ( 
.A(n_3226),
.B(n_74),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3191),
.B(n_3282),
.Y(n_3399)
);

BUFx2_ASAP7_75t_L g3400 ( 
.A(n_3222),
.Y(n_3400)
);

OR2x2_ASAP7_75t_L g3401 ( 
.A(n_3278),
.B(n_74),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3217),
.Y(n_3402)
);

NAND2x1_ASAP7_75t_L g3403 ( 
.A(n_3229),
.B(n_75),
.Y(n_3403)
);

INVx2_ASAP7_75t_SL g3404 ( 
.A(n_3275),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3195),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_3274),
.B(n_75),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3195),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3188),
.B(n_76),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3188),
.B(n_77),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3195),
.Y(n_3410)
);

AND2x4_ASAP7_75t_L g3411 ( 
.A(n_3275),
.B(n_77),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3195),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3188),
.B(n_78),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_3275),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3289),
.B(n_79),
.Y(n_3415)
);

BUFx3_ASAP7_75t_L g3416 ( 
.A(n_3275),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3182),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3188),
.B(n_79),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3188),
.B(n_80),
.Y(n_3419)
);

HB1xp67_ASAP7_75t_L g3420 ( 
.A(n_3195),
.Y(n_3420)
);

HB1xp67_ASAP7_75t_L g3421 ( 
.A(n_3195),
.Y(n_3421)
);

INVx5_ASAP7_75t_L g3422 ( 
.A(n_3201),
.Y(n_3422)
);

BUFx3_ASAP7_75t_L g3423 ( 
.A(n_3275),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3289),
.B(n_81),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3206),
.A2(n_1569),
.B1(n_1586),
.B2(n_1547),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3188),
.B(n_81),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3182),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3195),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_SL g3429 ( 
.A1(n_3228),
.A2(n_1600),
.B1(n_1601),
.B2(n_1593),
.Y(n_3429)
);

HB1xp67_ASAP7_75t_L g3430 ( 
.A(n_3195),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3195),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3195),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3195),
.Y(n_3433)
);

AND2x2_ASAP7_75t_L g3434 ( 
.A(n_3188),
.B(n_82),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3188),
.B(n_83),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3182),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3195),
.Y(n_3437)
);

OR2x2_ASAP7_75t_L g3438 ( 
.A(n_3289),
.B(n_83),
.Y(n_3438)
);

NAND2x1p5_ASAP7_75t_L g3439 ( 
.A(n_3269),
.B(n_84),
.Y(n_3439)
);

OR2x2_ASAP7_75t_L g3440 ( 
.A(n_3289),
.B(n_85),
.Y(n_3440)
);

AO21x2_ASAP7_75t_L g3441 ( 
.A1(n_3182),
.A2(n_85),
.B(n_86),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3195),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3289),
.B(n_87),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3188),
.B(n_87),
.Y(n_3444)
);

OA21x2_ASAP7_75t_L g3445 ( 
.A1(n_3194),
.A2(n_1610),
.B(n_1609),
.Y(n_3445)
);

AOI221xp5_ASAP7_75t_L g3446 ( 
.A1(n_3230),
.A2(n_1627),
.B1(n_1630),
.B2(n_1623),
.C(n_1613),
.Y(n_3446)
);

OAI221xp5_ASAP7_75t_L g3447 ( 
.A1(n_3303),
.A2(n_1669),
.B1(n_1680),
.B2(n_1666),
.C(n_1659),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3416),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3422),
.B(n_88),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3423),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3422),
.Y(n_3451)
);

OAI321xp33_ASAP7_75t_L g3452 ( 
.A1(n_3425),
.A2(n_93),
.A3(n_95),
.B1(n_90),
.B2(n_91),
.C(n_94),
.Y(n_3452)
);

OAI221xp5_ASAP7_75t_L g3453 ( 
.A1(n_3320),
.A2(n_1726),
.B1(n_1728),
.B2(n_1696),
.C(n_1689),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3381),
.A2(n_1732),
.B(n_1731),
.Y(n_3454)
);

INVx1_ASAP7_75t_SL g3455 ( 
.A(n_3302),
.Y(n_3455)
);

OAI221xp5_ASAP7_75t_L g3456 ( 
.A1(n_3389),
.A2(n_1781),
.B1(n_1788),
.B2(n_1756),
.C(n_1753),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3390),
.A2(n_1854),
.B1(n_1805),
.B2(n_93),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3414),
.B(n_90),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3332),
.B(n_91),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3308),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3358),
.B(n_94),
.Y(n_3461)
);

OAI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3349),
.A2(n_3323),
.B(n_3309),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3338),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3300),
.Y(n_3464)
);

INVxp67_ASAP7_75t_SL g3465 ( 
.A(n_3445),
.Y(n_3465)
);

INVx2_ASAP7_75t_SL g3466 ( 
.A(n_3314),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_SL g3467 ( 
.A(n_3304),
.B(n_95),
.Y(n_3467)
);

OR2x2_ASAP7_75t_L g3468 ( 
.A(n_3340),
.B(n_96),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3404),
.B(n_3312),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3310),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_L g3471 ( 
.A1(n_3361),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3318),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3331),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3420),
.B(n_98),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_L g3475 ( 
.A(n_3365),
.B(n_99),
.Y(n_3475)
);

OAI211xp5_ASAP7_75t_L g3476 ( 
.A1(n_3375),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_3476)
);

OA21x2_ASAP7_75t_L g3477 ( 
.A1(n_3294),
.A2(n_3305),
.B(n_3292),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3334),
.Y(n_3478)
);

OAI221xp5_ASAP7_75t_L g3479 ( 
.A1(n_3316),
.A2(n_3322),
.B1(n_3399),
.B2(n_3394),
.C(n_3352),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3421),
.Y(n_3480)
);

AO21x2_ASAP7_75t_L g3481 ( 
.A1(n_3415),
.A2(n_101),
.B(n_103),
.Y(n_3481)
);

OAI21xp33_ASAP7_75t_L g3482 ( 
.A1(n_3376),
.A2(n_3378),
.B(n_3293),
.Y(n_3482)
);

OR2x2_ASAP7_75t_L g3483 ( 
.A(n_3405),
.B(n_103),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3430),
.B(n_104),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3407),
.Y(n_3485)
);

AND2x2_ASAP7_75t_L g3486 ( 
.A(n_3295),
.B(n_104),
.Y(n_3486)
);

OAI22xp5_ASAP7_75t_L g3487 ( 
.A1(n_3438),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_3487)
);

BUFx2_ASAP7_75t_L g3488 ( 
.A(n_3306),
.Y(n_3488)
);

BUFx2_ASAP7_75t_L g3489 ( 
.A(n_3306),
.Y(n_3489)
);

OAI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3440),
.A2(n_108),
.B1(n_105),
.B2(n_106),
.Y(n_3490)
);

AOI221xp5_ASAP7_75t_L g3491 ( 
.A1(n_3387),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.C(n_111),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3336),
.B(n_109),
.Y(n_3492)
);

BUFx3_ASAP7_75t_L g3493 ( 
.A(n_3298),
.Y(n_3493)
);

OAI222xp33_ASAP7_75t_L g3494 ( 
.A1(n_3315),
.A2(n_136),
.B1(n_118),
.B2(n_145),
.C1(n_127),
.C2(n_110),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_L g3495 ( 
.A(n_3355),
.B(n_111),
.Y(n_3495)
);

OAI221xp5_ASAP7_75t_L g3496 ( 
.A1(n_3363),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.C(n_115),
.Y(n_3496)
);

OAI211xp5_ASAP7_75t_L g3497 ( 
.A1(n_3408),
.A2(n_3409),
.B(n_3418),
.C(n_3413),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_3419),
.B(n_3426),
.Y(n_3498)
);

NAND3xp33_ASAP7_75t_SL g3499 ( 
.A(n_3400),
.B(n_113),
.C(n_114),
.Y(n_3499)
);

OAI221xp5_ASAP7_75t_L g3500 ( 
.A1(n_3403),
.A2(n_119),
.B1(n_116),
.B2(n_117),
.C(n_120),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3441),
.Y(n_3501)
);

OAI33xp33_ASAP7_75t_L g3502 ( 
.A1(n_3410),
.A2(n_122),
.A3(n_124),
.B1(n_116),
.B2(n_119),
.B3(n_123),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3412),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3397),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3428),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3431),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3434),
.B(n_125),
.Y(n_3507)
);

OAI21x1_ASAP7_75t_L g3508 ( 
.A1(n_3417),
.A2(n_125),
.B(n_126),
.Y(n_3508)
);

OA21x2_ASAP7_75t_L g3509 ( 
.A1(n_3427),
.A2(n_127),
.B(n_128),
.Y(n_3509)
);

CKINVDCx5p33_ASAP7_75t_R g3510 ( 
.A(n_3356),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3432),
.B(n_3433),
.Y(n_3511)
);

OAI21xp33_ASAP7_75t_L g3512 ( 
.A1(n_3437),
.A2(n_129),
.B(n_130),
.Y(n_3512)
);

OR2x6_ASAP7_75t_L g3513 ( 
.A(n_3439),
.B(n_129),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_3435),
.B(n_130),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3444),
.B(n_131),
.Y(n_3515)
);

OAI211xp5_ASAP7_75t_L g3516 ( 
.A1(n_3406),
.A2(n_134),
.B(n_131),
.C(n_132),
.Y(n_3516)
);

OAI33xp33_ASAP7_75t_L g3517 ( 
.A1(n_3442),
.A2(n_137),
.A3(n_139),
.B1(n_134),
.B2(n_135),
.B3(n_138),
.Y(n_3517)
);

AOI221xp5_ASAP7_75t_L g3518 ( 
.A1(n_3391),
.A2(n_143),
.B1(n_140),
.B2(n_141),
.C(n_144),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3313),
.B(n_140),
.Y(n_3519)
);

OAI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3317),
.A2(n_3324),
.B1(n_3328),
.B2(n_3319),
.Y(n_3520)
);

OAI22xp5_ASAP7_75t_L g3521 ( 
.A1(n_3329),
.A2(n_145),
.B1(n_141),
.B2(n_143),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3343),
.B(n_146),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_3362),
.B(n_146),
.Y(n_3523)
);

OAI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3296),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_3524)
);

OAI31xp33_ASAP7_75t_L g3525 ( 
.A1(n_3369),
.A2(n_3348),
.A3(n_3350),
.B(n_3398),
.Y(n_3525)
);

OAI221xp5_ASAP7_75t_L g3526 ( 
.A1(n_3353),
.A2(n_150),
.B1(n_147),
.B2(n_148),
.C(n_152),
.Y(n_3526)
);

INVx1_ASAP7_75t_SL g3527 ( 
.A(n_3366),
.Y(n_3527)
);

AOI22xp33_ASAP7_75t_L g3528 ( 
.A1(n_3370),
.A2(n_3392),
.B1(n_3436),
.B2(n_3380),
.Y(n_3528)
);

OA21x2_ASAP7_75t_L g3529 ( 
.A1(n_3326),
.A2(n_152),
.B(n_153),
.Y(n_3529)
);

OR2x2_ASAP7_75t_L g3530 ( 
.A(n_3299),
.B(n_154),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3325),
.B(n_3341),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3424),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3443),
.Y(n_3533)
);

INVx3_ASAP7_75t_L g3534 ( 
.A(n_3411),
.Y(n_3534)
);

AOI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_3368),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_3535)
);

NAND3xp33_ASAP7_75t_L g3536 ( 
.A(n_3384),
.B(n_155),
.C(n_156),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_3346),
.Y(n_3537)
);

AOI221xp5_ASAP7_75t_L g3538 ( 
.A1(n_3360),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.C(n_160),
.Y(n_3538)
);

AOI221xp5_ASAP7_75t_L g3539 ( 
.A1(n_3359),
.A2(n_161),
.B1(n_157),
.B2(n_158),
.C(n_162),
.Y(n_3539)
);

BUFx3_ASAP7_75t_L g3540 ( 
.A(n_3344),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3333),
.A2(n_164),
.B1(n_161),
.B2(n_163),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3311),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3297),
.B(n_164),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_3301),
.B(n_165),
.Y(n_3544)
);

AND2x6_ASAP7_75t_L g3545 ( 
.A(n_3342),
.B(n_165),
.Y(n_3545)
);

OAI33xp33_ASAP7_75t_L g3546 ( 
.A1(n_3371),
.A2(n_168),
.A3(n_170),
.B1(n_166),
.B2(n_167),
.B3(n_169),
.Y(n_3546)
);

AO21x2_ASAP7_75t_L g3547 ( 
.A1(n_3335),
.A2(n_167),
.B(n_168),
.Y(n_3547)
);

AOI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_3385),
.A2(n_169),
.B(n_170),
.Y(n_3548)
);

AND2x4_ASAP7_75t_L g3549 ( 
.A(n_3307),
.B(n_171),
.Y(n_3549)
);

BUFx3_ASAP7_75t_L g3550 ( 
.A(n_3354),
.Y(n_3550)
);

AOI222xp33_ASAP7_75t_SL g3551 ( 
.A1(n_3347),
.A2(n_175),
.B1(n_177),
.B2(n_172),
.C1(n_174),
.C2(n_176),
.Y(n_3551)
);

INVxp67_ASAP7_75t_L g3552 ( 
.A(n_3367),
.Y(n_3552)
);

AOI221xp5_ASAP7_75t_L g3553 ( 
.A1(n_3351),
.A2(n_175),
.B1(n_172),
.B2(n_174),
.C(n_176),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3372),
.B(n_3386),
.Y(n_3554)
);

AND2x4_ASAP7_75t_L g3555 ( 
.A(n_3345),
.B(n_178),
.Y(n_3555)
);

INVxp67_ASAP7_75t_L g3556 ( 
.A(n_3402),
.Y(n_3556)
);

OAI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_3337),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_3557)
);

AOI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_3395),
.A2(n_183),
.B1(n_179),
.B2(n_182),
.Y(n_3558)
);

INVx4_ASAP7_75t_L g3559 ( 
.A(n_3373),
.Y(n_3559)
);

BUFx2_ASAP7_75t_L g3560 ( 
.A(n_3330),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3339),
.B(n_184),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3374),
.Y(n_3562)
);

OA21x2_ASAP7_75t_L g3563 ( 
.A1(n_3388),
.A2(n_184),
.B(n_186),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_3401),
.B(n_186),
.Y(n_3564)
);

HB1xp67_ASAP7_75t_L g3565 ( 
.A(n_3364),
.Y(n_3565)
);

AND2x4_ASAP7_75t_L g3566 ( 
.A(n_3377),
.B(n_187),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3379),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_3382),
.Y(n_3568)
);

INVx3_ASAP7_75t_L g3569 ( 
.A(n_3393),
.Y(n_3569)
);

AOI221xp5_ASAP7_75t_L g3570 ( 
.A1(n_3383),
.A2(n_190),
.B1(n_187),
.B2(n_188),
.C(n_191),
.Y(n_3570)
);

OAI33xp33_ASAP7_75t_L g3571 ( 
.A1(n_3357),
.A2(n_193),
.A3(n_195),
.B1(n_191),
.B2(n_192),
.B3(n_194),
.Y(n_3571)
);

AOI21xp33_ASAP7_75t_L g3572 ( 
.A1(n_3429),
.A2(n_194),
.B(n_196),
.Y(n_3572)
);

AOI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_3396),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_3573)
);

OA21x2_ASAP7_75t_L g3574 ( 
.A1(n_3327),
.A2(n_197),
.B(n_198),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3321),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3446),
.B(n_199),
.Y(n_3576)
);

AOI221xp5_ASAP7_75t_L g3577 ( 
.A1(n_3390),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3416),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3422),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_3390),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3308),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3308),
.Y(n_3582)
);

AOI22xp33_ASAP7_75t_SL g3583 ( 
.A1(n_3390),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_3583)
);

NOR3xp33_ASAP7_75t_SL g3584 ( 
.A(n_3314),
.B(n_206),
.C(n_207),
.Y(n_3584)
);

OAI221xp5_ASAP7_75t_L g3585 ( 
.A1(n_3303),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.C(n_212),
.Y(n_3585)
);

AOI22xp33_ASAP7_75t_L g3586 ( 
.A1(n_3390),
.A2(n_213),
.B1(n_208),
.B2(n_212),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3308),
.Y(n_3587)
);

AOI33xp33_ASAP7_75t_L g3588 ( 
.A1(n_3375),
.A2(n_216),
.A3(n_218),
.B1(n_213),
.B2(n_215),
.B3(n_217),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3422),
.B(n_216),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3422),
.B(n_218),
.Y(n_3590)
);

OAI321xp33_ASAP7_75t_L g3591 ( 
.A1(n_3303),
.A2(n_221),
.A3(n_223),
.B1(n_219),
.B2(n_220),
.C(n_222),
.Y(n_3591)
);

OAI22xp33_ASAP7_75t_L g3592 ( 
.A1(n_3390),
.A2(n_229),
.B1(n_237),
.B2(n_219),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3422),
.B(n_220),
.Y(n_3593)
);

BUFx3_ASAP7_75t_L g3594 ( 
.A(n_3302),
.Y(n_3594)
);

OAI22xp33_ASAP7_75t_L g3595 ( 
.A1(n_3390),
.A2(n_231),
.B1(n_240),
.B2(n_221),
.Y(n_3595)
);

OAI33xp33_ASAP7_75t_L g3596 ( 
.A1(n_3375),
.A2(n_225),
.A3(n_227),
.B1(n_222),
.B2(n_224),
.B3(n_226),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3308),
.Y(n_3597)
);

AOI22xp33_ASAP7_75t_SL g3598 ( 
.A1(n_3390),
.A2(n_230),
.B1(n_227),
.B2(n_229),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3416),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3416),
.Y(n_3600)
);

AOI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3390),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_3601)
);

HB1xp67_ASAP7_75t_L g3602 ( 
.A(n_3308),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3308),
.Y(n_3603)
);

AOI211xp5_ASAP7_75t_L g3604 ( 
.A1(n_3375),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_3604)
);

AOI221xp5_ASAP7_75t_L g3605 ( 
.A1(n_3390),
.A2(n_236),
.B1(n_233),
.B2(n_234),
.C(n_237),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3308),
.Y(n_3606)
);

AND2x2_ASAP7_75t_L g3607 ( 
.A(n_3422),
.B(n_236),
.Y(n_3607)
);

NAND3xp33_ASAP7_75t_L g3608 ( 
.A(n_3389),
.B(n_239),
.C(n_240),
.Y(n_3608)
);

OAI33xp33_ASAP7_75t_L g3609 ( 
.A1(n_3375),
.A2(n_243),
.A3(n_246),
.B1(n_239),
.B2(n_241),
.B3(n_244),
.Y(n_3609)
);

AOI221xp5_ASAP7_75t_L g3610 ( 
.A1(n_3390),
.A2(n_247),
.B1(n_243),
.B2(n_244),
.C(n_248),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3308),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3358),
.B(n_247),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3308),
.Y(n_3613)
);

AND2x2_ASAP7_75t_L g3614 ( 
.A(n_3422),
.B(n_249),
.Y(n_3614)
);

OAI221xp5_ASAP7_75t_L g3615 ( 
.A1(n_3303),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.C(n_252),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_SL g3616 ( 
.A1(n_3390),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3422),
.B(n_253),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3422),
.B(n_253),
.Y(n_3618)
);

AOI22xp5_ASAP7_75t_L g3619 ( 
.A1(n_3389),
.A2(n_257),
.B1(n_254),
.B2(n_256),
.Y(n_3619)
);

INVx3_ASAP7_75t_L g3620 ( 
.A(n_3302),
.Y(n_3620)
);

INVxp33_ASAP7_75t_L g3621 ( 
.A(n_3302),
.Y(n_3621)
);

INVx1_ASAP7_75t_SL g3622 ( 
.A(n_3302),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3308),
.Y(n_3623)
);

AOI322xp5_ASAP7_75t_L g3624 ( 
.A1(n_3390),
.A2(n_261),
.A3(n_260),
.B1(n_257),
.B2(n_254),
.C1(n_256),
.C2(n_258),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_3416),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_3422),
.B(n_258),
.Y(n_3626)
);

AOI22xp33_ASAP7_75t_L g3627 ( 
.A1(n_3390),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_3627)
);

HB1xp67_ASAP7_75t_L g3628 ( 
.A(n_3308),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3416),
.Y(n_3629)
);

NAND2xp33_ASAP7_75t_SL g3630 ( 
.A(n_3304),
.B(n_262),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3308),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3390),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3308),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_3416),
.Y(n_3634)
);

AOI22xp33_ASAP7_75t_L g3635 ( 
.A1(n_3390),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3308),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3475),
.B(n_267),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_3621),
.B(n_268),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3465),
.B(n_272),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3602),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3540),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3498),
.B(n_272),
.Y(n_3642)
);

OR2x2_ASAP7_75t_L g3643 ( 
.A(n_3511),
.B(n_3480),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3510),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3628),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3469),
.B(n_273),
.Y(n_3646)
);

HB1xp67_ASAP7_75t_L g3647 ( 
.A(n_3448),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3464),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3537),
.A2(n_273),
.B(n_274),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3488),
.B(n_275),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3450),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3547),
.B(n_275),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3578),
.Y(n_3653)
);

OR2x2_ASAP7_75t_L g3654 ( 
.A(n_3468),
.B(n_276),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3489),
.B(n_3599),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3600),
.B(n_276),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3625),
.B(n_277),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3629),
.B(n_277),
.Y(n_3658)
);

INVxp67_ASAP7_75t_L g3659 ( 
.A(n_3594),
.Y(n_3659)
);

INVxp67_ASAP7_75t_SL g3660 ( 
.A(n_3620),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3481),
.B(n_278),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3523),
.B(n_278),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_3634),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3470),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3451),
.B(n_3455),
.Y(n_3665)
);

AND2x4_ASAP7_75t_L g3666 ( 
.A(n_3493),
.B(n_280),
.Y(n_3666)
);

BUFx3_ASAP7_75t_L g3667 ( 
.A(n_3545),
.Y(n_3667)
);

AND2x2_ASAP7_75t_L g3668 ( 
.A(n_3622),
.B(n_3534),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3466),
.B(n_3458),
.Y(n_3669)
);

HB1xp67_ASAP7_75t_L g3670 ( 
.A(n_3531),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3529),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3472),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3473),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_3459),
.B(n_280),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3550),
.Y(n_3675)
);

NOR2xp67_ASAP7_75t_L g3676 ( 
.A(n_3559),
.B(n_281),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_3589),
.B(n_281),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3590),
.B(n_282),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3478),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3593),
.B(n_282),
.Y(n_3680)
);

INVx4_ASAP7_75t_L g3681 ( 
.A(n_3607),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3460),
.Y(n_3682)
);

HB1xp67_ASAP7_75t_L g3683 ( 
.A(n_3532),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3509),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3614),
.B(n_283),
.Y(n_3685)
);

HB1xp67_ASAP7_75t_L g3686 ( 
.A(n_3533),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3617),
.B(n_283),
.Y(n_3687)
);

HB1xp67_ASAP7_75t_L g3688 ( 
.A(n_3483),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3463),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3581),
.Y(n_3690)
);

INVx3_ASAP7_75t_L g3691 ( 
.A(n_3549),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3626),
.B(n_284),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_SL g3693 ( 
.A(n_3520),
.B(n_285),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3582),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_3497),
.B(n_286),
.Y(n_3695)
);

AND2x2_ASAP7_75t_L g3696 ( 
.A(n_3482),
.B(n_286),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3552),
.B(n_287),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3587),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3597),
.Y(n_3699)
);

INVxp67_ASAP7_75t_SL g3700 ( 
.A(n_3454),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3603),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3606),
.B(n_288),
.Y(n_3702)
);

AND2x4_ASAP7_75t_L g3703 ( 
.A(n_3522),
.B(n_289),
.Y(n_3703)
);

OR2x2_ASAP7_75t_L g3704 ( 
.A(n_3611),
.B(n_3613),
.Y(n_3704)
);

NAND2x1_ASAP7_75t_L g3705 ( 
.A(n_3623),
.B(n_289),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3631),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3633),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3636),
.B(n_290),
.Y(n_3708)
);

INVx3_ASAP7_75t_L g3709 ( 
.A(n_3513),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3561),
.B(n_3495),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3485),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3503),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3505),
.B(n_290),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3506),
.B(n_291),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3563),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3474),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3484),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3560),
.B(n_291),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3486),
.B(n_292),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3461),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3555),
.Y(n_3721)
);

AND2x4_ASAP7_75t_L g3722 ( 
.A(n_3543),
.B(n_293),
.Y(n_3722)
);

INVx3_ASAP7_75t_L g3723 ( 
.A(n_3513),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3507),
.B(n_294),
.Y(n_3724)
);

INVxp67_ASAP7_75t_L g3725 ( 
.A(n_3545),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3612),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3514),
.B(n_294),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3492),
.B(n_295),
.Y(n_3728)
);

AND2x4_ASAP7_75t_L g3729 ( 
.A(n_3544),
.B(n_295),
.Y(n_3729)
);

BUFx2_ASAP7_75t_L g3730 ( 
.A(n_3630),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3477),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3515),
.B(n_296),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3501),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3519),
.B(n_296),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3527),
.B(n_297),
.Y(n_3735)
);

INVx1_ASAP7_75t_SL g3736 ( 
.A(n_3545),
.Y(n_3736)
);

INVx1_ASAP7_75t_SL g3737 ( 
.A(n_3530),
.Y(n_3737)
);

AND2x2_ASAP7_75t_L g3738 ( 
.A(n_3618),
.B(n_297),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3556),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3565),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3535),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3467),
.B(n_299),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3508),
.Y(n_3743)
);

AND2x4_ASAP7_75t_L g3744 ( 
.A(n_3462),
.B(n_299),
.Y(n_3744)
);

INVx2_ASAP7_75t_SL g3745 ( 
.A(n_3449),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3554),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3567),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3542),
.Y(n_3748)
);

OR2x2_ASAP7_75t_L g3749 ( 
.A(n_3569),
.B(n_300),
.Y(n_3749)
);

NOR2xp33_ASAP7_75t_L g3750 ( 
.A(n_3536),
.B(n_300),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3457),
.B(n_301),
.Y(n_3751)
);

AND2x2_ASAP7_75t_L g3752 ( 
.A(n_3584),
.B(n_301),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3574),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3619),
.B(n_3548),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3541),
.B(n_302),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3574),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3524),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3562),
.B(n_302),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3592),
.B(n_303),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3568),
.Y(n_3760)
);

OR2x2_ASAP7_75t_L g3761 ( 
.A(n_3487),
.B(n_303),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3596),
.B(n_304),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3566),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3512),
.B(n_304),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3490),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3608),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3588),
.Y(n_3767)
);

AND2x2_ASAP7_75t_L g3768 ( 
.A(n_3575),
.B(n_305),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3576),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_3525),
.B(n_305),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3660),
.B(n_3668),
.Y(n_3771)
);

AOI22xp33_ASAP7_75t_L g3772 ( 
.A1(n_3741),
.A2(n_3479),
.B1(n_3546),
.B2(n_3609),
.Y(n_3772)
);

OA21x2_ASAP7_75t_L g3773 ( 
.A1(n_3731),
.A2(n_3528),
.B(n_3577),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3667),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3665),
.B(n_3598),
.Y(n_3775)
);

OAI22xp5_ASAP7_75t_L g3776 ( 
.A1(n_3730),
.A2(n_3604),
.B1(n_3616),
.B2(n_3583),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3688),
.Y(n_3777)
);

AOI33xp33_ASAP7_75t_L g3778 ( 
.A1(n_3740),
.A2(n_3586),
.A3(n_3601),
.B1(n_3632),
.B2(n_3627),
.B3(n_3580),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3670),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3669),
.B(n_3579),
.Y(n_3780)
);

INVxp67_ASAP7_75t_SL g3781 ( 
.A(n_3676),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3659),
.B(n_3564),
.Y(n_3782)
);

AND2x2_ASAP7_75t_SL g3783 ( 
.A(n_3730),
.B(n_3605),
.Y(n_3783)
);

AND2x4_ASAP7_75t_L g3784 ( 
.A(n_3655),
.B(n_3558),
.Y(n_3784)
);

NOR2xp67_ASAP7_75t_L g3785 ( 
.A(n_3681),
.B(n_3499),
.Y(n_3785)
);

OAI33xp33_ASAP7_75t_L g3786 ( 
.A1(n_3640),
.A2(n_3595),
.A3(n_3521),
.B1(n_3557),
.B2(n_3551),
.B3(n_3624),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3683),
.Y(n_3787)
);

AND2x4_ASAP7_75t_SL g3788 ( 
.A(n_3644),
.B(n_3647),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3686),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3697),
.Y(n_3790)
);

OR2x2_ASAP7_75t_SL g3791 ( 
.A(n_3641),
.B(n_3516),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3709),
.Y(n_3792)
);

OAI31xp33_ASAP7_75t_L g3793 ( 
.A1(n_3715),
.A2(n_3476),
.A3(n_3494),
.B(n_3526),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3695),
.A2(n_3635),
.B1(n_3610),
.B2(n_3496),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3737),
.B(n_3553),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3642),
.Y(n_3796)
);

NAND3xp33_ASAP7_75t_L g3797 ( 
.A(n_3675),
.B(n_3491),
.C(n_3538),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3723),
.Y(n_3798)
);

OAI31xp33_ASAP7_75t_L g3799 ( 
.A1(n_3754),
.A2(n_3500),
.A3(n_3456),
.B(n_3585),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_SL g3800 ( 
.A(n_3736),
.B(n_3502),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3705),
.Y(n_3801)
);

AND2x2_ASAP7_75t_L g3802 ( 
.A(n_3646),
.B(n_3471),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3718),
.B(n_3570),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3735),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3702),
.B(n_3504),
.Y(n_3805)
);

OAI31xp33_ASAP7_75t_L g3806 ( 
.A1(n_3753),
.A2(n_3615),
.A3(n_3572),
.B(n_3573),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3708),
.B(n_3518),
.Y(n_3807)
);

AO22x1_ASAP7_75t_L g3808 ( 
.A1(n_3744),
.A2(n_3517),
.B1(n_3571),
.B2(n_3452),
.Y(n_3808)
);

OAI22xp5_ASAP7_75t_L g3809 ( 
.A1(n_3765),
.A2(n_3539),
.B1(n_3447),
.B2(n_3453),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3700),
.B(n_306),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3747),
.Y(n_3811)
);

OAI221xp5_ASAP7_75t_L g3812 ( 
.A1(n_3756),
.A2(n_3591),
.B1(n_308),
.B2(n_306),
.C(n_307),
.Y(n_3812)
);

NAND4xp25_ASAP7_75t_L g3813 ( 
.A(n_3645),
.B(n_309),
.C(n_307),
.D(n_308),
.Y(n_3813)
);

AND2x2_ASAP7_75t_L g3814 ( 
.A(n_3691),
.B(n_310),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3650),
.B(n_310),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3654),
.Y(n_3816)
);

OR2x2_ASAP7_75t_L g3817 ( 
.A(n_3704),
.B(n_311),
.Y(n_3817)
);

OAI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3693),
.A2(n_3710),
.B(n_3770),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3722),
.Y(n_3819)
);

INVxp67_ASAP7_75t_L g3820 ( 
.A(n_3762),
.Y(n_3820)
);

OR2x2_ASAP7_75t_L g3821 ( 
.A(n_3643),
.B(n_312),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3639),
.Y(n_3822)
);

INVx3_ASAP7_75t_L g3823 ( 
.A(n_3666),
.Y(n_3823)
);

AOI22xp5_ASAP7_75t_L g3824 ( 
.A1(n_3769),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.Y(n_3824)
);

AND2x4_ASAP7_75t_L g3825 ( 
.A(n_3651),
.B(n_313),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3653),
.B(n_316),
.Y(n_3826)
);

INVx1_ASAP7_75t_SL g3827 ( 
.A(n_3719),
.Y(n_3827)
);

OAI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3739),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3663),
.B(n_317),
.Y(n_3829)
);

OR2x2_ASAP7_75t_L g3830 ( 
.A(n_3716),
.B(n_318),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3760),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3696),
.B(n_320),
.Y(n_3832)
);

NAND4xp25_ASAP7_75t_L g3833 ( 
.A(n_3682),
.B(n_322),
.C(n_320),
.D(n_321),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3713),
.B(n_321),
.Y(n_3834)
);

OR2x2_ASAP7_75t_L g3835 ( 
.A(n_3717),
.B(n_322),
.Y(n_3835)
);

OAI22xp5_ASAP7_75t_L g3836 ( 
.A1(n_3757),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3714),
.B(n_324),
.Y(n_3837)
);

NAND2x1_ASAP7_75t_L g3838 ( 
.A(n_3671),
.B(n_325),
.Y(n_3838)
);

NAND3xp33_ASAP7_75t_L g3839 ( 
.A(n_3766),
.B(n_327),
.C(n_328),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3729),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3767),
.B(n_327),
.Y(n_3841)
);

AOI22xp33_ASAP7_75t_L g3842 ( 
.A1(n_3684),
.A2(n_331),
.B1(n_328),
.B2(n_329),
.Y(n_3842)
);

AOI33xp33_ASAP7_75t_L g3843 ( 
.A1(n_3689),
.A2(n_359),
.A3(n_341),
.B1(n_369),
.B2(n_351),
.B3(n_332),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3721),
.B(n_332),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_SL g3845 ( 
.A1(n_3750),
.A2(n_333),
.B(n_334),
.Y(n_3845)
);

AND2x2_ASAP7_75t_L g3846 ( 
.A(n_3638),
.B(n_3690),
.Y(n_3846)
);

AOI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_3745),
.A2(n_336),
.B1(n_333),
.B2(n_334),
.Y(n_3847)
);

OAI322xp33_ASAP7_75t_L g3848 ( 
.A1(n_3694),
.A2(n_343),
.A3(n_342),
.B1(n_339),
.B2(n_337),
.C1(n_338),
.C2(n_340),
.Y(n_3848)
);

XOR2xp5_ASAP7_75t_L g3849 ( 
.A(n_3734),
.B(n_337),
.Y(n_3849)
);

INVx1_ASAP7_75t_SL g3850 ( 
.A(n_3724),
.Y(n_3850)
);

NOR3xp33_ASAP7_75t_L g3851 ( 
.A(n_3725),
.B(n_338),
.C(n_339),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3749),
.Y(n_3852)
);

NAND3xp33_ASAP7_75t_L g3853 ( 
.A(n_3720),
.B(n_3726),
.C(n_3699),
.Y(n_3853)
);

NAND2x1p5_ASAP7_75t_SL g3854 ( 
.A(n_3733),
.B(n_340),
.Y(n_3854)
);

OR2x2_ASAP7_75t_L g3855 ( 
.A(n_3698),
.B(n_342),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3701),
.B(n_3706),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3758),
.B(n_344),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3763),
.B(n_344),
.Y(n_3858)
);

OR2x2_ASAP7_75t_L g3859 ( 
.A(n_3707),
.B(n_345),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3827),
.B(n_3727),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3810),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3841),
.Y(n_3862)
);

INVxp67_ASAP7_75t_SL g3863 ( 
.A(n_3771),
.Y(n_3863)
);

AND2x2_ASAP7_75t_L g3864 ( 
.A(n_3788),
.B(n_3780),
.Y(n_3864)
);

OR2x2_ASAP7_75t_L g3865 ( 
.A(n_3850),
.B(n_3711),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3821),
.Y(n_3866)
);

OR2x2_ASAP7_75t_L g3867 ( 
.A(n_3817),
.B(n_3712),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3834),
.Y(n_3868)
);

OR2x2_ASAP7_75t_L g3869 ( 
.A(n_3779),
.B(n_3648),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3837),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3808),
.B(n_3732),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3783),
.B(n_3661),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3830),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3801),
.B(n_3664),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3846),
.B(n_3672),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3804),
.B(n_3652),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3807),
.B(n_3746),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3835),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3823),
.B(n_3673),
.Y(n_3879)
);

AO21x1_ASAP7_75t_L g3880 ( 
.A1(n_3776),
.A2(n_3800),
.B(n_3793),
.Y(n_3880)
);

BUFx2_ASAP7_75t_L g3881 ( 
.A(n_3782),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3815),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3777),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3855),
.Y(n_3884)
);

HB1xp67_ASAP7_75t_L g3885 ( 
.A(n_3785),
.Y(n_3885)
);

AND2x4_ASAP7_75t_L g3886 ( 
.A(n_3774),
.B(n_3656),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3859),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3856),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3816),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3822),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3826),
.B(n_3677),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3825),
.Y(n_3892)
);

NOR2xp33_ASAP7_75t_SL g3893 ( 
.A(n_3781),
.B(n_3678),
.Y(n_3893)
);

OR2x2_ASAP7_75t_L g3894 ( 
.A(n_3791),
.B(n_3679),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3792),
.B(n_3657),
.Y(n_3895)
);

INVx2_ASAP7_75t_L g3896 ( 
.A(n_3844),
.Y(n_3896)
);

OR2x2_ASAP7_75t_L g3897 ( 
.A(n_3787),
.B(n_3637),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3829),
.B(n_3680),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3838),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3775),
.B(n_3685),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3789),
.B(n_3798),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3857),
.Y(n_3902)
);

OR2x2_ASAP7_75t_L g3903 ( 
.A(n_3820),
.B(n_3728),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3814),
.B(n_3658),
.Y(n_3904)
);

NOR2xp33_ASAP7_75t_L g3905 ( 
.A(n_3786),
.B(n_3858),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3851),
.B(n_3687),
.Y(n_3906)
);

NOR2xp33_ASAP7_75t_L g3907 ( 
.A(n_3796),
.B(n_3662),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3784),
.B(n_3674),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3832),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3790),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3852),
.B(n_3692),
.Y(n_3911)
);

INVx3_ASAP7_75t_L g3912 ( 
.A(n_3819),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3843),
.Y(n_3913)
);

INVxp67_ASAP7_75t_L g3914 ( 
.A(n_3893),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3881),
.Y(n_3915)
);

INVxp67_ASAP7_75t_SL g3916 ( 
.A(n_3880),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3864),
.B(n_3818),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3863),
.B(n_3840),
.Y(n_3918)
);

OAI33xp33_ASAP7_75t_L g3919 ( 
.A1(n_3894),
.A2(n_3831),
.A3(n_3811),
.B1(n_3795),
.B2(n_3853),
.B3(n_3794),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3903),
.Y(n_3920)
);

HB1xp67_ASAP7_75t_L g3921 ( 
.A(n_3885),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3908),
.B(n_3802),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3860),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3868),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3875),
.B(n_3805),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3870),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3882),
.B(n_3778),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3901),
.B(n_3752),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3904),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3867),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3879),
.B(n_3824),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3895),
.Y(n_3932)
);

OAI221xp5_ASAP7_75t_L g3933 ( 
.A1(n_3872),
.A2(n_3772),
.B1(n_3806),
.B2(n_3773),
.C(n_3812),
.Y(n_3933)
);

AND2x2_ASAP7_75t_L g3934 ( 
.A(n_3888),
.B(n_3803),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3874),
.B(n_3742),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3886),
.B(n_3738),
.Y(n_3936)
);

OR2x2_ASAP7_75t_L g3937 ( 
.A(n_3865),
.B(n_3813),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3897),
.B(n_3799),
.Y(n_3938)
);

INVx1_ASAP7_75t_SL g3939 ( 
.A(n_3900),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3866),
.B(n_3842),
.Y(n_3940)
);

OR2x2_ASAP7_75t_L g3941 ( 
.A(n_3869),
.B(n_3833),
.Y(n_3941)
);

OAI21xp33_ASAP7_75t_SL g3942 ( 
.A1(n_3905),
.A2(n_3845),
.B(n_3847),
.Y(n_3942)
);

INVxp67_ASAP7_75t_L g3943 ( 
.A(n_3899),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3907),
.B(n_3836),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_SL g3945 ( 
.A1(n_3871),
.A2(n_3773),
.B1(n_3797),
.B2(n_3751),
.Y(n_3945)
);

OR2x6_ASAP7_75t_L g3946 ( 
.A(n_3912),
.B(n_3768),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3883),
.B(n_3913),
.Y(n_3947)
);

INVx1_ASAP7_75t_SL g3948 ( 
.A(n_3891),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3890),
.B(n_3809),
.Y(n_3949)
);

INVx2_ASAP7_75t_SL g3950 ( 
.A(n_3911),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3862),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3877),
.B(n_3854),
.Y(n_3952)
);

OR2x2_ASAP7_75t_L g3953 ( 
.A(n_3910),
.B(n_3839),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_SL g3954 ( 
.A(n_3916),
.B(n_3906),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3921),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3918),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3925),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3922),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3939),
.B(n_3873),
.Y(n_3959)
);

OR2x2_ASAP7_75t_L g3960 ( 
.A(n_3929),
.B(n_3915),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3917),
.B(n_3884),
.Y(n_3961)
);

HB1xp67_ASAP7_75t_L g3962 ( 
.A(n_3914),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3928),
.B(n_3887),
.Y(n_3963)
);

OR2x2_ASAP7_75t_L g3964 ( 
.A(n_3948),
.B(n_3950),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3946),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3938),
.B(n_3878),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3934),
.B(n_3902),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3935),
.B(n_3861),
.Y(n_3968)
);

AND4x1_ASAP7_75t_L g3969 ( 
.A(n_3919),
.B(n_3909),
.C(n_3889),
.D(n_3876),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3949),
.Y(n_3970)
);

NAND2x1p5_ASAP7_75t_L g3971 ( 
.A(n_3932),
.B(n_3920),
.Y(n_3971)
);

OAI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3942),
.A2(n_3898),
.B(n_3759),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3936),
.B(n_3896),
.Y(n_3973)
);

NAND2x1p5_ASAP7_75t_L g3974 ( 
.A(n_3930),
.B(n_3764),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3952),
.B(n_3892),
.Y(n_3975)
);

OAI31xp33_ASAP7_75t_L g3976 ( 
.A1(n_3933),
.A2(n_3761),
.A3(n_3755),
.B(n_3828),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3923),
.B(n_3703),
.Y(n_3977)
);

OR2x2_ASAP7_75t_L g3978 ( 
.A(n_3937),
.B(n_3748),
.Y(n_3978)
);

OAI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3945),
.A2(n_3849),
.B(n_3649),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3947),
.B(n_3743),
.Y(n_3980)
);

XNOR2xp5_ASAP7_75t_L g3981 ( 
.A(n_3946),
.B(n_3848),
.Y(n_3981)
);

AND2x2_ASAP7_75t_L g3982 ( 
.A(n_3924),
.B(n_345),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3931),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3926),
.B(n_346),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3941),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3943),
.B(n_347),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3940),
.Y(n_3987)
);

OR2x2_ASAP7_75t_L g3988 ( 
.A(n_3953),
.B(n_350),
.Y(n_3988)
);

OR2x2_ASAP7_75t_L g3989 ( 
.A(n_3951),
.B(n_352),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3944),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3927),
.B(n_352),
.Y(n_3991)
);

OR2x2_ASAP7_75t_L g3992 ( 
.A(n_3939),
.B(n_353),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3917),
.B(n_353),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3946),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3961),
.B(n_354),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_SL g3996 ( 
.A1(n_3980),
.A2(n_3979),
.B1(n_3963),
.B2(n_3987),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3970),
.B(n_355),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3993),
.B(n_355),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3957),
.B(n_356),
.Y(n_3999)
);

BUFx2_ASAP7_75t_L g4000 ( 
.A(n_3971),
.Y(n_4000)
);

AND2x2_ASAP7_75t_L g4001 ( 
.A(n_3956),
.B(n_357),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3983),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3974),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3968),
.B(n_357),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3966),
.Y(n_4005)
);

NAND3xp33_ASAP7_75t_L g4006 ( 
.A(n_3969),
.B(n_358),
.C(n_360),
.Y(n_4006)
);

AOI22xp33_ASAP7_75t_SL g4007 ( 
.A1(n_3975),
.A2(n_361),
.B1(n_358),
.B2(n_360),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_L g4008 ( 
.A(n_3990),
.B(n_361),
.Y(n_4008)
);

INVx2_ASAP7_75t_L g4009 ( 
.A(n_3992),
.Y(n_4009)
);

INVx1_ASAP7_75t_SL g4010 ( 
.A(n_3964),
.Y(n_4010)
);

OR2x2_ASAP7_75t_L g4011 ( 
.A(n_3967),
.B(n_3960),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3962),
.B(n_362),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3977),
.Y(n_4013)
);

AND2x4_ASAP7_75t_L g4014 ( 
.A(n_3965),
.B(n_364),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3958),
.B(n_366),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3954),
.A2(n_368),
.B(n_367),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3988),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_SL g4018 ( 
.A1(n_3991),
.A2(n_3972),
.B1(n_3959),
.B2(n_3994),
.Y(n_4018)
);

AOI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_3981),
.A2(n_377),
.B1(n_385),
.B2(n_366),
.Y(n_4019)
);

AOI221x1_ASAP7_75t_SL g4020 ( 
.A1(n_3955),
.A2(n_3973),
.B1(n_3985),
.B2(n_3986),
.C(n_3978),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3982),
.B(n_368),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3984),
.B(n_369),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_3989),
.B(n_370),
.Y(n_4023)
);

INVx3_ASAP7_75t_SL g4024 ( 
.A(n_3976),
.Y(n_4024)
);

XOR2xp5_ASAP7_75t_L g4025 ( 
.A(n_3981),
.B(n_370),
.Y(n_4025)
);

NAND3xp33_ASAP7_75t_L g4026 ( 
.A(n_3969),
.B(n_371),
.C(n_373),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3961),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_3961),
.B(n_371),
.Y(n_4028)
);

OR2x2_ASAP7_75t_L g4029 ( 
.A(n_3971),
.B(n_373),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3971),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3961),
.Y(n_4031)
);

OAI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_3954),
.A2(n_374),
.B(n_376),
.Y(n_4032)
);

AND2x4_ASAP7_75t_SL g4033 ( 
.A(n_3962),
.B(n_376),
.Y(n_4033)
);

AOI22x1_ASAP7_75t_L g4034 ( 
.A1(n_3962),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3970),
.B(n_378),
.Y(n_4035)
);

NOR2x1_ASAP7_75t_L g4036 ( 
.A(n_3964),
.B(n_380),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3970),
.B(n_381),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_3961),
.B(n_381),
.Y(n_4038)
);

NAND2x1p5_ASAP7_75t_L g4039 ( 
.A(n_3964),
.B(n_382),
.Y(n_4039)
);

INVx2_ASAP7_75t_SL g4040 ( 
.A(n_3971),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3970),
.B(n_382),
.Y(n_4041)
);

OR2x2_ASAP7_75t_L g4042 ( 
.A(n_3971),
.B(n_383),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3970),
.B(n_383),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_3961),
.B(n_384),
.Y(n_4044)
);

NOR2xp33_ASAP7_75t_L g4045 ( 
.A(n_4000),
.B(n_384),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_4011),
.Y(n_4046)
);

AOI22xp5_ASAP7_75t_L g4047 ( 
.A1(n_4006),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_4039),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3995),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_4040),
.B(n_386),
.Y(n_4050)
);

O2A1O1Ixp33_ASAP7_75t_L g4051 ( 
.A1(n_4026),
.A2(n_4024),
.B(n_4032),
.C(n_4030),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_4028),
.B(n_387),
.Y(n_4052)
);

OA21x2_ASAP7_75t_L g4053 ( 
.A1(n_4016),
.A2(n_388),
.B(n_389),
.Y(n_4053)
);

OAI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_4010),
.A2(n_392),
.B1(n_389),
.B2(n_391),
.Y(n_4054)
);

O2A1O1Ixp33_ASAP7_75t_L g4055 ( 
.A1(n_4003),
.A2(n_395),
.B(n_393),
.C(n_394),
.Y(n_4055)
);

INVx1_ASAP7_75t_SL g4056 ( 
.A(n_4029),
.Y(n_4056)
);

OR2x2_ASAP7_75t_L g4057 ( 
.A(n_4027),
.B(n_395),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_4038),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_4031),
.B(n_396),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_4005),
.B(n_397),
.Y(n_4060)
);

AOI21xp5_ASAP7_75t_L g4061 ( 
.A1(n_4044),
.A2(n_398),
.B(n_399),
.Y(n_4061)
);

AOI21xp33_ASAP7_75t_L g4062 ( 
.A1(n_4036),
.A2(n_398),
.B(n_399),
.Y(n_4062)
);

HB1xp67_ASAP7_75t_L g4063 ( 
.A(n_4004),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_4033),
.B(n_400),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_4013),
.B(n_402),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3996),
.B(n_403),
.Y(n_4066)
);

INVx2_ASAP7_75t_SL g4067 ( 
.A(n_4042),
.Y(n_4067)
);

OAI21xp33_ASAP7_75t_L g4068 ( 
.A1(n_4018),
.A2(n_404),
.B(n_405),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_4025),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_4012),
.B(n_406),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3998),
.Y(n_4071)
);

OAI21xp5_ASAP7_75t_L g4072 ( 
.A1(n_4002),
.A2(n_407),
.B(n_408),
.Y(n_4072)
);

NOR4xp25_ASAP7_75t_L g4073 ( 
.A(n_4017),
.B(n_410),
.C(n_408),
.D(n_409),
.Y(n_4073)
);

OAI211xp5_ASAP7_75t_L g4074 ( 
.A1(n_3999),
.A2(n_413),
.B(n_409),
.C(n_412),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_4007),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_4075)
);

OR2x2_ASAP7_75t_L g4076 ( 
.A(n_3997),
.B(n_414),
.Y(n_4076)
);

INVx1_ASAP7_75t_SL g4077 ( 
.A(n_4023),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4021),
.Y(n_4078)
);

OAI31xp33_ASAP7_75t_L g4079 ( 
.A1(n_4008),
.A2(n_417),
.A3(n_415),
.B(n_416),
.Y(n_4079)
);

AOI211xp5_ASAP7_75t_SL g4080 ( 
.A1(n_4035),
.A2(n_419),
.B(n_417),
.C(n_418),
.Y(n_4080)
);

AOI32xp33_ASAP7_75t_L g4081 ( 
.A1(n_4009),
.A2(n_420),
.A3(n_418),
.B1(n_419),
.B2(n_421),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_4022),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_4019),
.B(n_420),
.Y(n_4083)
);

OAI22xp33_ASAP7_75t_L g4084 ( 
.A1(n_4037),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_4084)
);

INVx2_ASAP7_75t_SL g4085 ( 
.A(n_4001),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_4015),
.B(n_422),
.Y(n_4086)
);

AOI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_4041),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_4087)
);

OAI22xp33_ASAP7_75t_L g4088 ( 
.A1(n_4043),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_4088)
);

AOI21xp33_ASAP7_75t_SL g4089 ( 
.A1(n_4034),
.A2(n_427),
.B(n_428),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_4014),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_4020),
.B(n_429),
.Y(n_4091)
);

AOI21xp33_ASAP7_75t_L g4092 ( 
.A1(n_4006),
.A2(n_429),
.B(n_430),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4011),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_4011),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4011),
.Y(n_4095)
);

AOI22xp5_ASAP7_75t_L g4096 ( 
.A1(n_4006),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_4096)
);

AOI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_4006),
.A2(n_431),
.B(n_432),
.Y(n_4097)
);

AOI21xp5_ASAP7_75t_SL g4098 ( 
.A1(n_4040),
.A2(n_434),
.B(n_435),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_4000),
.B(n_434),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_4000),
.B(n_435),
.Y(n_4100)
);

AOI21xp5_ASAP7_75t_L g4101 ( 
.A1(n_4006),
.A2(n_436),
.B(n_437),
.Y(n_4101)
);

OAI31xp33_ASAP7_75t_L g4102 ( 
.A1(n_4006),
.A2(n_439),
.A3(n_436),
.B(n_438),
.Y(n_4102)
);

AOI222xp33_ASAP7_75t_L g4103 ( 
.A1(n_4006),
.A2(n_441),
.B1(n_443),
.B2(n_439),
.C1(n_440),
.C2(n_442),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_4000),
.B(n_440),
.Y(n_4104)
);

AOI32xp33_ASAP7_75t_L g4105 ( 
.A1(n_3996),
.A2(n_445),
.A3(n_441),
.B1(n_442),
.B2(n_446),
.Y(n_4105)
);

AOI321xp33_ASAP7_75t_L g4106 ( 
.A1(n_4003),
.A2(n_451),
.A3(n_453),
.B1(n_448),
.B2(n_450),
.C(n_452),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_4000),
.B(n_448),
.Y(n_4107)
);

INVxp67_ASAP7_75t_L g4108 ( 
.A(n_4000),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_4011),
.Y(n_4109)
);

HB1xp67_ASAP7_75t_L g4110 ( 
.A(n_4000),
.Y(n_4110)
);

OAI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_4006),
.A2(n_450),
.B(n_452),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4011),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_4039),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4000),
.B(n_453),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4011),
.Y(n_4115)
);

AOI32xp33_ASAP7_75t_L g4116 ( 
.A1(n_3996),
.A2(n_456),
.A3(n_454),
.B1(n_455),
.B2(n_457),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_4000),
.B(n_455),
.Y(n_4117)
);

INVxp67_ASAP7_75t_SL g4118 ( 
.A(n_4000),
.Y(n_4118)
);

AOI21xp33_ASAP7_75t_SL g4119 ( 
.A1(n_4040),
.A2(n_456),
.B(n_458),
.Y(n_4119)
);

OAI221xp5_ASAP7_75t_L g4120 ( 
.A1(n_4006),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.C(n_461),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_4011),
.Y(n_4121)
);

OAI21xp33_ASAP7_75t_SL g4122 ( 
.A1(n_4040),
.A2(n_459),
.B(n_462),
.Y(n_4122)
);

OAI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_4006),
.A2(n_465),
.B1(n_462),
.B2(n_463),
.Y(n_4123)
);

NOR2xp33_ASAP7_75t_L g4124 ( 
.A(n_4000),
.B(n_463),
.Y(n_4124)
);

OR2x2_ASAP7_75t_L g4125 ( 
.A(n_4011),
.B(n_465),
.Y(n_4125)
);

O2A1O1Ixp33_ASAP7_75t_L g4126 ( 
.A1(n_4006),
.A2(n_468),
.B(n_466),
.C(n_467),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4011),
.Y(n_4127)
);

XOR2x2_ASAP7_75t_L g4128 ( 
.A(n_4063),
.B(n_4080),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_SL g4129 ( 
.A(n_4122),
.B(n_466),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_4125),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_4110),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_4118),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4086),
.Y(n_4133)
);

OR2x2_ASAP7_75t_L g4134 ( 
.A(n_4046),
.B(n_467),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4073),
.B(n_469),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_4070),
.B(n_469),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_4053),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4093),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4094),
.Y(n_4139)
);

OR2x2_ASAP7_75t_L g4140 ( 
.A(n_4095),
.B(n_470),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4109),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4112),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4115),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4121),
.Y(n_4144)
);

OR2x2_ASAP7_75t_L g4145 ( 
.A(n_4127),
.B(n_470),
.Y(n_4145)
);

NOR2xp33_ASAP7_75t_L g4146 ( 
.A(n_4119),
.B(n_471),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4052),
.Y(n_4147)
);

OR2x2_ASAP7_75t_L g4148 ( 
.A(n_4056),
.B(n_471),
.Y(n_4148)
);

NOR2xp33_ASAP7_75t_L g4149 ( 
.A(n_4089),
.B(n_472),
.Y(n_4149)
);

OR2x2_ASAP7_75t_L g4150 ( 
.A(n_4108),
.B(n_472),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4050),
.B(n_4067),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4045),
.B(n_473),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4106),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4066),
.Y(n_4154)
);

AOI21xp33_ASAP7_75t_SL g4155 ( 
.A1(n_4051),
.A2(n_474),
.B(n_476),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4065),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_4098),
.B(n_4068),
.Y(n_4157)
);

AOI321xp33_ASAP7_75t_L g4158 ( 
.A1(n_4049),
.A2(n_478),
.A3(n_480),
.B1(n_476),
.B2(n_477),
.C(n_479),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_4124),
.B(n_478),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_4059),
.B(n_481),
.Y(n_4160)
);

OR2x2_ASAP7_75t_L g4161 ( 
.A(n_4099),
.B(n_482),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4060),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_4048),
.B(n_482),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_4113),
.B(n_483),
.Y(n_4164)
);

OR2x2_ASAP7_75t_L g4165 ( 
.A(n_4100),
.B(n_484),
.Y(n_4165)
);

INVxp33_ASAP7_75t_L g4166 ( 
.A(n_4053),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_4085),
.B(n_484),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_4077),
.B(n_485),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4057),
.Y(n_4169)
);

OAI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_4104),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_4058),
.B(n_487),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_4076),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4064),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4090),
.Y(n_4174)
);

OR2x2_ASAP7_75t_L g4175 ( 
.A(n_4107),
.B(n_4114),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_4061),
.B(n_489),
.Y(n_4176)
);

INVx1_ASAP7_75t_SL g4177 ( 
.A(n_4117),
.Y(n_4177)
);

INVx2_ASAP7_75t_SL g4178 ( 
.A(n_4091),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4071),
.Y(n_4179)
);

INVx1_ASAP7_75t_SL g4180 ( 
.A(n_4078),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_4111),
.B(n_490),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4082),
.Y(n_4182)
);

INVx1_ASAP7_75t_SL g4183 ( 
.A(n_4062),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4074),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4069),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_L g4186 ( 
.A(n_4120),
.B(n_490),
.Y(n_4186)
);

INVx1_ASAP7_75t_SL g4187 ( 
.A(n_4083),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4105),
.B(n_491),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4116),
.B(n_491),
.Y(n_4189)
);

OAI321xp33_ASAP7_75t_L g4190 ( 
.A1(n_4123),
.A2(n_494),
.A3(n_496),
.B1(n_492),
.B2(n_493),
.C(n_495),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4055),
.Y(n_4191)
);

OR2x2_ASAP7_75t_L g4192 ( 
.A(n_4054),
.B(n_494),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_4072),
.B(n_495),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4087),
.Y(n_4194)
);

NOR2xp33_ASAP7_75t_L g4195 ( 
.A(n_4075),
.B(n_496),
.Y(n_4195)
);

INVxp67_ASAP7_75t_L g4196 ( 
.A(n_4103),
.Y(n_4196)
);

OAI21xp5_ASAP7_75t_SL g4197 ( 
.A1(n_4102),
.A2(n_497),
.B(n_498),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4047),
.Y(n_4198)
);

INVx3_ASAP7_75t_L g4199 ( 
.A(n_4081),
.Y(n_4199)
);

INVx2_ASAP7_75t_L g4200 ( 
.A(n_4096),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4097),
.B(n_497),
.Y(n_4201)
);

OR2x2_ASAP7_75t_L g4202 ( 
.A(n_4101),
.B(n_498),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4126),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_4079),
.B(n_499),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_4084),
.Y(n_4205)
);

OR2x2_ASAP7_75t_L g4206 ( 
.A(n_4092),
.B(n_499),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_SL g4207 ( 
.A(n_4088),
.B(n_500),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4063),
.Y(n_4208)
);

INVx2_ASAP7_75t_SL g4209 ( 
.A(n_4110),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4063),
.B(n_500),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4137),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4128),
.Y(n_4212)
);

AOI31xp33_ASAP7_75t_L g4213 ( 
.A1(n_4209),
.A2(n_503),
.A3(n_501),
.B(n_502),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4160),
.Y(n_4214)
);

OAI31xp33_ASAP7_75t_L g4215 ( 
.A1(n_4166),
.A2(n_4157),
.A3(n_4154),
.B(n_4153),
.Y(n_4215)
);

AOI21xp33_ASAP7_75t_L g4216 ( 
.A1(n_4177),
.A2(n_501),
.B(n_502),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4132),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_4151),
.Y(n_4218)
);

NOR2xp33_ASAP7_75t_L g4219 ( 
.A(n_4129),
.B(n_503),
.Y(n_4219)
);

AOI222xp33_ASAP7_75t_L g4220 ( 
.A1(n_4183),
.A2(n_506),
.B1(n_508),
.B2(n_504),
.C1(n_505),
.C2(n_507),
.Y(n_4220)
);

XNOR2xp5_ASAP7_75t_L g4221 ( 
.A(n_4133),
.B(n_506),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4152),
.B(n_504),
.Y(n_4222)
);

OAI21xp33_ASAP7_75t_L g4223 ( 
.A1(n_4131),
.A2(n_4208),
.B(n_4180),
.Y(n_4223)
);

AOI211xp5_ASAP7_75t_SL g4224 ( 
.A1(n_4138),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_4139),
.B(n_509),
.Y(n_4225)
);

OAI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_4141),
.A2(n_4142),
.B1(n_4144),
.B2(n_4143),
.Y(n_4226)
);

AOI22xp33_ASAP7_75t_L g4227 ( 
.A1(n_4178),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4135),
.Y(n_4228)
);

XOR2x2_ASAP7_75t_L g4229 ( 
.A(n_4207),
.B(n_511),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_4174),
.Y(n_4230)
);

OAI221xp5_ASAP7_75t_L g4231 ( 
.A1(n_4197),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.C(n_515),
.Y(n_4231)
);

AOI21xp33_ASAP7_75t_SL g4232 ( 
.A1(n_4149),
.A2(n_4146),
.B(n_4210),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4179),
.B(n_513),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4136),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4158),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_4159),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_4162),
.B(n_514),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_4148),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4134),
.Y(n_4239)
);

HB1xp67_ASAP7_75t_L g4240 ( 
.A(n_4130),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4140),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4145),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_4161),
.Y(n_4243)
);

A2O1A1Ixp33_ASAP7_75t_L g4244 ( 
.A1(n_4195),
.A2(n_4186),
.B(n_4196),
.C(n_4182),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4176),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4165),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4150),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4169),
.B(n_516),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_4175),
.Y(n_4249)
);

INVx1_ASAP7_75t_SL g4250 ( 
.A(n_4163),
.Y(n_4250)
);

AOI22xp5_ASAP7_75t_L g4251 ( 
.A1(n_4173),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_4251)
);

NAND3xp33_ASAP7_75t_L g4252 ( 
.A(n_4155),
.B(n_519),
.C(n_518),
.Y(n_4252)
);

AOI221xp5_ASAP7_75t_L g4253 ( 
.A1(n_4203),
.A2(n_520),
.B1(n_517),
.B2(n_519),
.C(n_521),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_SL g4254 ( 
.A(n_4190),
.B(n_522),
.Y(n_4254)
);

OAI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_4168),
.A2(n_522),
.B(n_523),
.Y(n_4255)
);

AOI21xp33_ASAP7_75t_SL g4256 ( 
.A1(n_4184),
.A2(n_523),
.B(n_524),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4164),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4187),
.B(n_525),
.Y(n_4258)
);

NAND2xp33_ASAP7_75t_SL g4259 ( 
.A(n_4188),
.B(n_525),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4172),
.Y(n_4260)
);

INVx1_ASAP7_75t_SL g4261 ( 
.A(n_4181),
.Y(n_4261)
);

NOR2xp33_ASAP7_75t_L g4262 ( 
.A(n_4191),
.B(n_526),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4156),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_4193),
.B(n_4147),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4167),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_4201),
.B(n_4199),
.Y(n_4266)
);

XNOR2x1_ASAP7_75t_L g4267 ( 
.A(n_4202),
.B(n_526),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4171),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4205),
.B(n_527),
.Y(n_4269)
);

OR2x2_ASAP7_75t_L g4270 ( 
.A(n_4189),
.B(n_527),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4204),
.Y(n_4271)
);

AOI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_4170),
.A2(n_528),
.B(n_529),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4198),
.B(n_529),
.Y(n_4273)
);

INVxp67_ASAP7_75t_L g4274 ( 
.A(n_4192),
.Y(n_4274)
);

AOI221xp5_ASAP7_75t_L g4275 ( 
.A1(n_4200),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.C(n_535),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4194),
.B(n_530),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4206),
.B(n_532),
.Y(n_4277)
);

XNOR2x1_ASAP7_75t_L g4278 ( 
.A(n_4185),
.B(n_535),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4137),
.Y(n_4279)
);

AOI211xp5_ASAP7_75t_L g4280 ( 
.A1(n_4208),
.A2(n_539),
.B(n_536),
.C(n_537),
.Y(n_4280)
);

NOR2xp33_ASAP7_75t_L g4281 ( 
.A(n_4166),
.B(n_537),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_4209),
.A2(n_539),
.B(n_541),
.Y(n_4282)
);

XNOR2x1_ASAP7_75t_L g4283 ( 
.A(n_4128),
.B(n_541),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4209),
.B(n_542),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4137),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4137),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4209),
.B(n_542),
.Y(n_4287)
);

OAI21xp33_ASAP7_75t_L g4288 ( 
.A1(n_4209),
.A2(n_543),
.B(n_544),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4137),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4209),
.B(n_545),
.Y(n_4290)
);

HB1xp67_ASAP7_75t_L g4291 ( 
.A(n_4137),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_4209),
.B(n_545),
.Y(n_4292)
);

OR2x2_ASAP7_75t_L g4293 ( 
.A(n_4209),
.B(n_546),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4137),
.Y(n_4294)
);

A2O1A1Ixp33_ASAP7_75t_L g4295 ( 
.A1(n_4178),
.A2(n_555),
.B(n_563),
.C(n_546),
.Y(n_4295)
);

AOI211xp5_ASAP7_75t_L g4296 ( 
.A1(n_4226),
.A2(n_549),
.B(n_547),
.C(n_548),
.Y(n_4296)
);

XNOR2x1_ASAP7_75t_L g4297 ( 
.A(n_4283),
.B(n_547),
.Y(n_4297)
);

AOI221xp5_ASAP7_75t_L g4298 ( 
.A1(n_4291),
.A2(n_551),
.B1(n_548),
.B2(n_549),
.C(n_552),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4224),
.B(n_553),
.Y(n_4299)
);

OAI221xp5_ASAP7_75t_L g4300 ( 
.A1(n_4215),
.A2(n_554),
.B1(n_552),
.B2(n_553),
.C(n_556),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4249),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4240),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4213),
.Y(n_4303)
);

XNOR2xp5_ASAP7_75t_L g4304 ( 
.A(n_4278),
.B(n_556),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4235),
.B(n_558),
.Y(n_4305)
);

OAI21xp33_ASAP7_75t_L g4306 ( 
.A1(n_4223),
.A2(n_557),
.B(n_558),
.Y(n_4306)
);

INVx3_ASAP7_75t_L g4307 ( 
.A(n_4218),
.Y(n_4307)
);

OR2x2_ASAP7_75t_L g4308 ( 
.A(n_4293),
.B(n_557),
.Y(n_4308)
);

AOI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_4282),
.A2(n_559),
.B(n_560),
.Y(n_4309)
);

AOI21xp33_ASAP7_75t_L g4310 ( 
.A1(n_4211),
.A2(n_559),
.B(n_560),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4279),
.Y(n_4311)
);

XNOR2x1_ASAP7_75t_L g4312 ( 
.A(n_4267),
.B(n_561),
.Y(n_4312)
);

XOR2xp5_ASAP7_75t_SL g4313 ( 
.A(n_4284),
.B(n_561),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_4285),
.Y(n_4314)
);

INVxp67_ASAP7_75t_L g4315 ( 
.A(n_4281),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4286),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4289),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4294),
.Y(n_4318)
);

NOR2xp33_ASAP7_75t_L g4319 ( 
.A(n_4230),
.B(n_562),
.Y(n_4319)
);

AO21x1_ASAP7_75t_L g4320 ( 
.A1(n_4290),
.A2(n_562),
.B(n_563),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4233),
.B(n_565),
.Y(n_4321)
);

OR2x2_ASAP7_75t_L g4322 ( 
.A(n_4292),
.B(n_564),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_SL g4323 ( 
.A(n_4256),
.B(n_565),
.Y(n_4323)
);

OAI221xp5_ASAP7_75t_L g4324 ( 
.A1(n_4212),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.C(n_569),
.Y(n_4324)
);

OR2x2_ASAP7_75t_L g4325 ( 
.A(n_4260),
.B(n_567),
.Y(n_4325)
);

OAI22xp5_ASAP7_75t_L g4326 ( 
.A1(n_4217),
.A2(n_570),
.B1(n_568),
.B2(n_569),
.Y(n_4326)
);

OAI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_4263),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_4327)
);

AND2x2_ASAP7_75t_L g4328 ( 
.A(n_4287),
.B(n_571),
.Y(n_4328)
);

XNOR2xp5_ASAP7_75t_L g4329 ( 
.A(n_4221),
.B(n_4229),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4225),
.B(n_573),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4222),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4220),
.B(n_572),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4214),
.Y(n_4333)
);

INVx2_ASAP7_75t_L g4334 ( 
.A(n_4243),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4236),
.Y(n_4335)
);

INVx1_ASAP7_75t_SL g4336 ( 
.A(n_4270),
.Y(n_4336)
);

NOR2xp33_ASAP7_75t_L g4337 ( 
.A(n_4261),
.B(n_574),
.Y(n_4337)
);

OAI322xp33_ASAP7_75t_L g4338 ( 
.A1(n_4228),
.A2(n_581),
.A3(n_580),
.B1(n_577),
.B2(n_575),
.C1(n_576),
.C2(n_579),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4238),
.Y(n_4339)
);

OR2x2_ASAP7_75t_L g4340 ( 
.A(n_4237),
.B(n_576),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4250),
.B(n_580),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_4254),
.A2(n_4288),
.B(n_4295),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4264),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4258),
.A2(n_579),
.B(n_581),
.Y(n_4344)
);

AOI21xp5_ASAP7_75t_L g4345 ( 
.A1(n_4231),
.A2(n_582),
.B(n_583),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_4246),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_L g4347 ( 
.A(n_4219),
.B(n_585),
.Y(n_4347)
);

O2A1O1Ixp33_ASAP7_75t_SL g4348 ( 
.A1(n_4244),
.A2(n_4280),
.B(n_4216),
.C(n_4248),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4239),
.Y(n_4349)
);

INVxp67_ASAP7_75t_SL g4350 ( 
.A(n_4266),
.Y(n_4350)
);

INVxp67_ASAP7_75t_L g4351 ( 
.A(n_4262),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4241),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4245),
.B(n_586),
.Y(n_4353)
);

OAI21xp33_ASAP7_75t_L g4354 ( 
.A1(n_4271),
.A2(n_582),
.B(n_586),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4242),
.Y(n_4355)
);

OAI211xp5_ASAP7_75t_SL g4356 ( 
.A1(n_4274),
.A2(n_590),
.B(n_587),
.C(n_589),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4257),
.Y(n_4357)
);

AOI22xp5_ASAP7_75t_L g4358 ( 
.A1(n_4265),
.A2(n_592),
.B1(n_589),
.B2(n_591),
.Y(n_4358)
);

NAND2x1_ASAP7_75t_L g4359 ( 
.A(n_4247),
.B(n_592),
.Y(n_4359)
);

OR2x2_ASAP7_75t_L g4360 ( 
.A(n_4252),
.B(n_593),
.Y(n_4360)
);

XOR2x2_ASAP7_75t_L g4361 ( 
.A(n_4269),
.B(n_593),
.Y(n_4361)
);

AOI221xp5_ASAP7_75t_L g4362 ( 
.A1(n_4232),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.C(n_597),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_4277),
.B(n_595),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4276),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4234),
.Y(n_4365)
);

XNOR2x1_ASAP7_75t_L g4366 ( 
.A(n_4255),
.B(n_594),
.Y(n_4366)
);

NAND5xp2_ASAP7_75t_L g4367 ( 
.A(n_4268),
.B(n_601),
.C(n_596),
.D(n_597),
.E(n_603),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4273),
.Y(n_4368)
);

OR2x2_ASAP7_75t_L g4369 ( 
.A(n_4227),
.B(n_4272),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_4251),
.B(n_603),
.Y(n_4370)
);

AND2x2_ASAP7_75t_L g4371 ( 
.A(n_4253),
.B(n_601),
.Y(n_4371)
);

CKINVDCx20_ASAP7_75t_R g4372 ( 
.A(n_4329),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4350),
.B(n_4275),
.Y(n_4373)
);

NAND4xp75_ASAP7_75t_L g4374 ( 
.A(n_4302),
.B(n_4259),
.C(n_606),
.D(n_604),
.Y(n_4374)
);

NOR2xp67_ASAP7_75t_L g4375 ( 
.A(n_4307),
.B(n_605),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4307),
.Y(n_4376)
);

AO22x1_ASAP7_75t_L g4377 ( 
.A1(n_4311),
.A2(n_4314),
.B1(n_4317),
.B2(n_4316),
.Y(n_4377)
);

NOR2x1_ASAP7_75t_L g4378 ( 
.A(n_4318),
.B(n_609),
.Y(n_4378)
);

NOR2x1_ASAP7_75t_L g4379 ( 
.A(n_4301),
.B(n_4343),
.Y(n_4379)
);

NAND5xp2_ASAP7_75t_L g4380 ( 
.A(n_4342),
.B(n_611),
.C(n_609),
.D(n_610),
.E(n_612),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4320),
.Y(n_4381)
);

NOR3xp33_ASAP7_75t_L g4382 ( 
.A(n_4300),
.B(n_610),
.C(n_611),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4359),
.Y(n_4383)
);

NOR3xp33_ASAP7_75t_L g4384 ( 
.A(n_4339),
.B(n_612),
.C(n_613),
.Y(n_4384)
);

NAND5xp2_ASAP7_75t_SL g4385 ( 
.A(n_4332),
.B(n_618),
.C(n_614),
.D(n_615),
.E(n_619),
.Y(n_4385)
);

NAND4xp75_ASAP7_75t_L g4386 ( 
.A(n_4349),
.B(n_620),
.C(n_615),
.D(n_618),
.Y(n_4386)
);

NOR3xp33_ASAP7_75t_L g4387 ( 
.A(n_4352),
.B(n_620),
.C(n_621),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4328),
.Y(n_4388)
);

NAND4xp25_ASAP7_75t_L g4389 ( 
.A(n_4355),
.B(n_623),
.C(n_621),
.D(n_622),
.Y(n_4389)
);

OAI211xp5_ASAP7_75t_SL g4390 ( 
.A1(n_4333),
.A2(n_625),
.B(n_622),
.C(n_624),
.Y(n_4390)
);

O2A1O1Ixp33_ASAP7_75t_L g4391 ( 
.A1(n_4335),
.A2(n_628),
.B(n_625),
.C(n_626),
.Y(n_4391)
);

NOR2xp33_ASAP7_75t_L g4392 ( 
.A(n_4367),
.B(n_628),
.Y(n_4392)
);

NOR2xp33_ASAP7_75t_L g4393 ( 
.A(n_4334),
.B(n_629),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4308),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4304),
.Y(n_4395)
);

NOR3xp33_ASAP7_75t_SL g4396 ( 
.A(n_4305),
.B(n_629),
.C(n_630),
.Y(n_4396)
);

INVx1_ASAP7_75t_SL g4397 ( 
.A(n_4297),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4299),
.Y(n_4398)
);

OAI22xp5_ASAP7_75t_L g4399 ( 
.A1(n_4357),
.A2(n_633),
.B1(n_631),
.B2(n_632),
.Y(n_4399)
);

NAND3xp33_ASAP7_75t_L g4400 ( 
.A(n_4319),
.B(n_631),
.C(n_634),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_SL g4401 ( 
.A(n_4346),
.B(n_634),
.Y(n_4401)
);

AO22x2_ASAP7_75t_L g4402 ( 
.A1(n_4312),
.A2(n_638),
.B1(n_635),
.B2(n_637),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4363),
.Y(n_4403)
);

AOI31xp33_ASAP7_75t_L g4404 ( 
.A1(n_4296),
.A2(n_639),
.A3(n_635),
.B(n_638),
.Y(n_4404)
);

INVxp67_ASAP7_75t_L g4405 ( 
.A(n_4337),
.Y(n_4405)
);

AOI211xp5_ASAP7_75t_L g4406 ( 
.A1(n_4306),
.A2(n_641),
.B(n_642),
.C(n_640),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4321),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4330),
.Y(n_4408)
);

NOR3xp33_ASAP7_75t_L g4409 ( 
.A(n_4365),
.B(n_639),
.C(n_640),
.Y(n_4409)
);

NOR2x1_ASAP7_75t_L g4410 ( 
.A(n_4338),
.B(n_641),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4325),
.Y(n_4411)
);

NAND5xp2_ASAP7_75t_L g4412 ( 
.A(n_4303),
.B(n_645),
.C(n_643),
.D(n_644),
.E(n_646),
.Y(n_4412)
);

NOR2x1_ASAP7_75t_L g4413 ( 
.A(n_4324),
.B(n_643),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4371),
.B(n_644),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4331),
.A2(n_649),
.B1(n_645),
.B2(n_648),
.Y(n_4415)
);

AND5x1_ASAP7_75t_L g4416 ( 
.A(n_4348),
.B(n_651),
.C(n_648),
.D(n_650),
.E(n_652),
.Y(n_4416)
);

NOR3xp33_ASAP7_75t_L g4417 ( 
.A(n_4341),
.B(n_650),
.C(n_651),
.Y(n_4417)
);

AOI22xp5_ASAP7_75t_L g4418 ( 
.A1(n_4370),
.A2(n_656),
.B1(n_653),
.B2(n_654),
.Y(n_4418)
);

NOR3xp33_ASAP7_75t_L g4419 ( 
.A(n_4336),
.B(n_653),
.C(n_654),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4361),
.Y(n_4420)
);

NOR3xp33_ASAP7_75t_L g4421 ( 
.A(n_4315),
.B(n_657),
.C(n_658),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4340),
.Y(n_4422)
);

NOR3xp33_ASAP7_75t_L g4423 ( 
.A(n_4368),
.B(n_657),
.C(n_658),
.Y(n_4423)
);

NOR2xp33_ASAP7_75t_L g4424 ( 
.A(n_4356),
.B(n_659),
.Y(n_4424)
);

NOR3x1_ASAP7_75t_L g4425 ( 
.A(n_4347),
.B(n_4353),
.C(n_4323),
.Y(n_4425)
);

HB1xp67_ASAP7_75t_L g4426 ( 
.A(n_4313),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4379),
.B(n_4309),
.Y(n_4427)
);

AOI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4377),
.A2(n_4354),
.B(n_4310),
.Y(n_4428)
);

HB1xp67_ASAP7_75t_L g4429 ( 
.A(n_4375),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_4381),
.B(n_4364),
.Y(n_4430)
);

OAI211xp5_ASAP7_75t_SL g4431 ( 
.A1(n_4376),
.A2(n_4351),
.B(n_4369),
.C(n_4298),
.Y(n_4431)
);

NOR2x1_ASAP7_75t_L g4432 ( 
.A(n_4372),
.B(n_4322),
.Y(n_4432)
);

NOR3x1_ASAP7_75t_L g4433 ( 
.A(n_4374),
.B(n_4360),
.C(n_4327),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4402),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4402),
.Y(n_4435)
);

NAND4xp25_ASAP7_75t_L g4436 ( 
.A(n_4425),
.B(n_4345),
.C(n_4344),
.D(n_4362),
.Y(n_4436)
);

AOI21xp33_ASAP7_75t_L g4437 ( 
.A1(n_4397),
.A2(n_4398),
.B(n_4383),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4378),
.Y(n_4438)
);

AND2x2_ASAP7_75t_SL g4439 ( 
.A(n_4419),
.B(n_4358),
.Y(n_4439)
);

INVx2_ASAP7_75t_SL g4440 ( 
.A(n_4426),
.Y(n_4440)
);

AOI22xp5_ASAP7_75t_L g4441 ( 
.A1(n_4392),
.A2(n_4366),
.B1(n_4326),
.B2(n_661),
.Y(n_4441)
);

OR2x2_ASAP7_75t_L g4442 ( 
.A(n_4412),
.B(n_659),
.Y(n_4442)
);

HB1xp67_ASAP7_75t_L g4443 ( 
.A(n_4416),
.Y(n_4443)
);

XNOR2xp5_ASAP7_75t_L g4444 ( 
.A(n_4396),
.B(n_660),
.Y(n_4444)
);

BUFx2_ASAP7_75t_R g4445 ( 
.A(n_4373),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4410),
.B(n_660),
.Y(n_4446)
);

INVx1_ASAP7_75t_SL g4447 ( 
.A(n_4386),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4388),
.Y(n_4448)
);

AOI21xp5_ASAP7_75t_L g4449 ( 
.A1(n_4401),
.A2(n_4391),
.B(n_4389),
.Y(n_4449)
);

AOI31xp33_ASAP7_75t_L g4450 ( 
.A1(n_4406),
.A2(n_663),
.A3(n_661),
.B(n_662),
.Y(n_4450)
);

AOI22xp33_ASAP7_75t_L g4451 ( 
.A1(n_4407),
.A2(n_665),
.B1(n_662),
.B2(n_664),
.Y(n_4451)
);

AOI211xp5_ASAP7_75t_L g4452 ( 
.A1(n_4424),
.A2(n_666),
.B(n_664),
.C(n_665),
.Y(n_4452)
);

OAI21xp33_ASAP7_75t_L g4453 ( 
.A1(n_4380),
.A2(n_667),
.B(n_668),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4394),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4422),
.Y(n_4455)
);

NOR2x1_ASAP7_75t_L g4456 ( 
.A(n_4400),
.B(n_668),
.Y(n_4456)
);

AOI322xp5_ASAP7_75t_L g4457 ( 
.A1(n_4395),
.A2(n_676),
.A3(n_675),
.B1(n_673),
.B2(n_669),
.C1(n_672),
.C2(n_674),
.Y(n_4457)
);

AOI221xp5_ASAP7_75t_L g4458 ( 
.A1(n_4405),
.A2(n_673),
.B1(n_669),
.B2(n_672),
.C(n_675),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4411),
.Y(n_4459)
);

INVxp67_ASAP7_75t_L g4460 ( 
.A(n_4393),
.Y(n_4460)
);

NAND4xp75_ASAP7_75t_L g4461 ( 
.A(n_4432),
.B(n_4420),
.C(n_4408),
.D(n_4403),
.Y(n_4461)
);

NAND3xp33_ASAP7_75t_SL g4462 ( 
.A(n_4438),
.B(n_4417),
.C(n_4409),
.Y(n_4462)
);

NAND4xp25_ASAP7_75t_L g4463 ( 
.A(n_4437),
.B(n_4382),
.C(n_4413),
.D(n_4414),
.Y(n_4463)
);

NAND3x1_ASAP7_75t_L g4464 ( 
.A(n_4427),
.B(n_4387),
.C(n_4423),
.Y(n_4464)
);

NOR2x1_ASAP7_75t_L g4465 ( 
.A(n_4430),
.B(n_4399),
.Y(n_4465)
);

INVxp33_ASAP7_75t_SL g4466 ( 
.A(n_4444),
.Y(n_4466)
);

NAND5xp2_ASAP7_75t_L g4467 ( 
.A(n_4455),
.B(n_4384),
.C(n_4421),
.D(n_4418),
.E(n_4415),
.Y(n_4467)
);

NAND3xp33_ASAP7_75t_SL g4468 ( 
.A(n_4447),
.B(n_4385),
.C(n_4404),
.Y(n_4468)
);

NOR2x1_ASAP7_75t_L g4469 ( 
.A(n_4431),
.B(n_4390),
.Y(n_4469)
);

NAND3xp33_ASAP7_75t_SL g4470 ( 
.A(n_4434),
.B(n_676),
.C(n_678),
.Y(n_4470)
);

NOR3x2_ASAP7_75t_L g4471 ( 
.A(n_4442),
.B(n_689),
.C(n_679),
.Y(n_4471)
);

NAND3x1_ASAP7_75t_L g4472 ( 
.A(n_4428),
.B(n_680),
.C(n_681),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4440),
.B(n_680),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4443),
.Y(n_4474)
);

NOR3x1_ASAP7_75t_L g4475 ( 
.A(n_4436),
.B(n_683),
.C(n_684),
.Y(n_4475)
);

AND2x4_ASAP7_75t_L g4476 ( 
.A(n_4448),
.B(n_686),
.Y(n_4476)
);

AND2x2_ASAP7_75t_SL g4477 ( 
.A(n_4446),
.B(n_683),
.Y(n_4477)
);

OAI31xp33_ASAP7_75t_L g4478 ( 
.A1(n_4474),
.A2(n_4453),
.A3(n_4435),
.B(n_4454),
.Y(n_4478)
);

NOR2xp33_ASAP7_75t_L g4479 ( 
.A(n_4466),
.B(n_4445),
.Y(n_4479)
);

AOI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_4465),
.A2(n_4468),
.B(n_4473),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4477),
.Y(n_4481)
);

OAI311xp33_ASAP7_75t_L g4482 ( 
.A1(n_4463),
.A2(n_4441),
.A3(n_4459),
.B1(n_4460),
.C1(n_4429),
.Y(n_4482)
);

AOI22xp5_ASAP7_75t_L g4483 ( 
.A1(n_4462),
.A2(n_4439),
.B1(n_4456),
.B2(n_4449),
.Y(n_4483)
);

OAI211xp5_ASAP7_75t_L g4484 ( 
.A1(n_4469),
.A2(n_4452),
.B(n_4451),
.C(n_4458),
.Y(n_4484)
);

AOI221xp5_ASAP7_75t_L g4485 ( 
.A1(n_4467),
.A2(n_4450),
.B1(n_4433),
.B2(n_4457),
.C(n_689),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4471),
.Y(n_4486)
);

AOI211xp5_ASAP7_75t_L g4487 ( 
.A1(n_4470),
.A2(n_690),
.B(n_687),
.C(n_688),
.Y(n_4487)
);

AOI211xp5_ASAP7_75t_L g4488 ( 
.A1(n_4476),
.A2(n_690),
.B(n_687),
.C(n_688),
.Y(n_4488)
);

AOI221xp5_ASAP7_75t_L g4489 ( 
.A1(n_4479),
.A2(n_4461),
.B1(n_4475),
.B2(n_4464),
.C(n_4472),
.Y(n_4489)
);

OAI22xp33_ASAP7_75t_L g4490 ( 
.A1(n_4483),
.A2(n_693),
.B1(n_691),
.B2(n_692),
.Y(n_4490)
);

AOI21xp5_ASAP7_75t_L g4491 ( 
.A1(n_4480),
.A2(n_4478),
.B(n_4485),
.Y(n_4491)
);

OR2x2_ASAP7_75t_L g4492 ( 
.A(n_4481),
.B(n_693),
.Y(n_4492)
);

HB1xp67_ASAP7_75t_L g4493 ( 
.A(n_4486),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4487),
.B(n_4488),
.Y(n_4494)
);

NAND3xp33_ASAP7_75t_SL g4495 ( 
.A(n_4484),
.B(n_4482),
.C(n_694),
.Y(n_4495)
);

AOI211xp5_ASAP7_75t_L g4496 ( 
.A1(n_4495),
.A2(n_697),
.B(n_694),
.C(n_695),
.Y(n_4496)
);

OAI21xp33_ASAP7_75t_L g4497 ( 
.A1(n_4489),
.A2(n_4493),
.B(n_4491),
.Y(n_4497)
);

NOR2x1_ASAP7_75t_L g4498 ( 
.A(n_4492),
.B(n_695),
.Y(n_4498)
);

AND2x4_ASAP7_75t_L g4499 ( 
.A(n_4494),
.B(n_698),
.Y(n_4499)
);

OAI211xp5_ASAP7_75t_SL g4500 ( 
.A1(n_4490),
.A2(n_700),
.B(n_698),
.C(n_699),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4497),
.B(n_699),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4498),
.B(n_700),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4499),
.Y(n_4503)
);

NOR4xp25_ASAP7_75t_L g4504 ( 
.A(n_4500),
.B(n_4496),
.C(n_704),
.D(n_702),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_SL g4505 ( 
.A(n_4502),
.B(n_703),
.Y(n_4505)
);

XOR2xp5_ASAP7_75t_L g4506 ( 
.A(n_4503),
.B(n_4501),
.Y(n_4506)
);

OAI222xp33_ASAP7_75t_L g4507 ( 
.A1(n_4504),
.A2(n_706),
.B1(n_708),
.B2(n_703),
.C1(n_705),
.C2(n_707),
.Y(n_4507)
);

OAI221xp5_ASAP7_75t_R g4508 ( 
.A1(n_4501),
.A2(n_709),
.B1(n_705),
.B2(n_706),
.C(n_710),
.Y(n_4508)
);

XNOR2xp5_ASAP7_75t_L g4509 ( 
.A(n_4503),
.B(n_709),
.Y(n_4509)
);

AND2x4_ASAP7_75t_L g4510 ( 
.A(n_4503),
.B(n_710),
.Y(n_4510)
);

AOI22xp5_ASAP7_75t_L g4511 ( 
.A1(n_4501),
.A2(n_715),
.B1(n_713),
.B2(n_714),
.Y(n_4511)
);

XNOR2xp5_ASAP7_75t_L g4512 ( 
.A(n_4506),
.B(n_714),
.Y(n_4512)
);

OAI21xp5_ASAP7_75t_L g4513 ( 
.A1(n_4505),
.A2(n_715),
.B(n_716),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4510),
.Y(n_4514)
);

XNOR2x1_ASAP7_75t_L g4515 ( 
.A(n_4509),
.B(n_717),
.Y(n_4515)
);

XNOR2x1_ASAP7_75t_L g4516 ( 
.A(n_4511),
.B(n_717),
.Y(n_4516)
);

XNOR2xp5_ASAP7_75t_L g4517 ( 
.A(n_4508),
.B(n_718),
.Y(n_4517)
);

OAI22xp5_ASAP7_75t_L g4518 ( 
.A1(n_4507),
.A2(n_720),
.B1(n_718),
.B2(n_719),
.Y(n_4518)
);

BUFx2_ASAP7_75t_L g4519 ( 
.A(n_4514),
.Y(n_4519)
);

OR3x1_ASAP7_75t_L g4520 ( 
.A(n_4517),
.B(n_720),
.C(n_722),
.Y(n_4520)
);

OR2x2_ASAP7_75t_SL g4521 ( 
.A(n_4515),
.B(n_4512),
.Y(n_4521)
);

AOI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_4513),
.A2(n_723),
.B(n_724),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4516),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4518),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4514),
.Y(n_4525)
);

OAI22xp5_ASAP7_75t_L g4526 ( 
.A1(n_4512),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.Y(n_4526)
);

AND3x4_ASAP7_75t_L g4527 ( 
.A(n_4514),
.B(n_725),
.C(n_727),
.Y(n_4527)
);

AOI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_4512),
.A2(n_729),
.B1(n_727),
.B2(n_728),
.Y(n_4528)
);

OAI22xp5_ASAP7_75t_L g4529 ( 
.A1(n_4512),
.A2(n_731),
.B1(n_728),
.B2(n_730),
.Y(n_4529)
);

AOI22xp5_ASAP7_75t_L g4530 ( 
.A1(n_4512),
.A2(n_733),
.B1(n_731),
.B2(n_732),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4514),
.B(n_734),
.Y(n_4531)
);

AND2x4_ASAP7_75t_L g4532 ( 
.A(n_4514),
.B(n_734),
.Y(n_4532)
);

AOI21x1_ASAP7_75t_L g4533 ( 
.A1(n_4519),
.A2(n_736),
.B(n_737),
.Y(n_4533)
);

AOI22xp5_ASAP7_75t_L g4534 ( 
.A1(n_4520),
.A2(n_739),
.B1(n_736),
.B2(n_737),
.Y(n_4534)
);

OAI22x1_ASAP7_75t_SL g4535 ( 
.A1(n_4525),
.A2(n_743),
.B1(n_739),
.B2(n_740),
.Y(n_4535)
);

HB1xp67_ASAP7_75t_L g4536 ( 
.A(n_4521),
.Y(n_4536)
);

AOI22xp5_ASAP7_75t_L g4537 ( 
.A1(n_4527),
.A2(n_748),
.B1(n_744),
.B2(n_745),
.Y(n_4537)
);

INVx1_ASAP7_75t_SL g4538 ( 
.A(n_4523),
.Y(n_4538)
);

AOI222xp33_ASAP7_75t_L g4539 ( 
.A1(n_4524),
.A2(n_750),
.B1(n_752),
.B2(n_744),
.C1(n_749),
.C2(n_751),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4532),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4531),
.Y(n_4541)
);

XNOR2x1_ASAP7_75t_SL g4542 ( 
.A(n_4522),
.B(n_4526),
.Y(n_4542)
);

NOR2xp33_ASAP7_75t_L g4543 ( 
.A(n_4529),
.B(n_749),
.Y(n_4543)
);

AOI22x1_ASAP7_75t_L g4544 ( 
.A1(n_4528),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_4530),
.Y(n_4545)
);

XNOR2xp5_ASAP7_75t_L g4546 ( 
.A(n_4519),
.B(n_753),
.Y(n_4546)
);

AO22x2_ASAP7_75t_L g4547 ( 
.A1(n_4525),
.A2(n_755),
.B1(n_753),
.B2(n_754),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4536),
.B(n_754),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4538),
.Y(n_4549)
);

AOI22xp5_ASAP7_75t_SL g4550 ( 
.A1(n_4540),
.A2(n_757),
.B1(n_755),
.B2(n_756),
.Y(n_4550)
);

AO22x2_ASAP7_75t_L g4551 ( 
.A1(n_4541),
.A2(n_758),
.B1(n_756),
.B2(n_757),
.Y(n_4551)
);

OR2x6_ASAP7_75t_L g4552 ( 
.A(n_4545),
.B(n_758),
.Y(n_4552)
);

OAI22xp5_ASAP7_75t_SL g4553 ( 
.A1(n_4534),
.A2(n_761),
.B1(n_759),
.B2(n_760),
.Y(n_4553)
);

XNOR2xp5_ASAP7_75t_L g4554 ( 
.A(n_4542),
.B(n_762),
.Y(n_4554)
);

AND5x1_ASAP7_75t_L g4555 ( 
.A(n_4543),
.B(n_765),
.C(n_762),
.D(n_763),
.E(n_766),
.Y(n_4555)
);

OR2x2_ASAP7_75t_L g4556 ( 
.A(n_4537),
.B(n_763),
.Y(n_4556)
);

AOI22xp5_ASAP7_75t_SL g4557 ( 
.A1(n_4546),
.A2(n_772),
.B1(n_769),
.B2(n_770),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4533),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_4544),
.Y(n_4559)
);

AOI221xp5_ASAP7_75t_L g4560 ( 
.A1(n_4549),
.A2(n_4547),
.B1(n_4535),
.B2(n_4539),
.C(n_773),
.Y(n_4560)
);

AOI21xp5_ASAP7_75t_L g4561 ( 
.A1(n_4558),
.A2(n_769),
.B(n_770),
.Y(n_4561)
);

OAI22xp5_ASAP7_75t_L g4562 ( 
.A1(n_4552),
.A2(n_777),
.B1(n_774),
.B2(n_776),
.Y(n_4562)
);

OAI21xp5_ASAP7_75t_L g4563 ( 
.A1(n_4554),
.A2(n_774),
.B(n_776),
.Y(n_4563)
);

AO22x2_ASAP7_75t_L g4564 ( 
.A1(n_4559),
.A2(n_779),
.B1(n_777),
.B2(n_778),
.Y(n_4564)
);

AOI222xp33_ASAP7_75t_L g4565 ( 
.A1(n_4553),
.A2(n_784),
.B1(n_786),
.B2(n_778),
.C1(n_779),
.C2(n_785),
.Y(n_4565)
);

OAI22xp33_ASAP7_75t_L g4566 ( 
.A1(n_4556),
.A2(n_788),
.B1(n_785),
.B2(n_787),
.Y(n_4566)
);

AOI21xp5_ASAP7_75t_L g4567 ( 
.A1(n_4548),
.A2(n_787),
.B(n_788),
.Y(n_4567)
);

AOI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_4557),
.A2(n_789),
.B(n_791),
.Y(n_4568)
);

OR2x2_ASAP7_75t_L g4569 ( 
.A(n_4550),
.B(n_789),
.Y(n_4569)
);

AOI222xp33_ASAP7_75t_L g4570 ( 
.A1(n_4563),
.A2(n_4551),
.B1(n_4555),
.B2(n_793),
.C1(n_795),
.C2(n_791),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4569),
.Y(n_4571)
);

AOI222xp33_ASAP7_75t_L g4572 ( 
.A1(n_4560),
.A2(n_794),
.B1(n_796),
.B2(n_792),
.C1(n_793),
.C2(n_795),
.Y(n_4572)
);

NOR3xp33_ASAP7_75t_L g4573 ( 
.A(n_4568),
.B(n_794),
.C(n_797),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4567),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4566),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4561),
.Y(n_4576)
);

AOI222xp33_ASAP7_75t_L g4577 ( 
.A1(n_4571),
.A2(n_4576),
.B1(n_4574),
.B2(n_4575),
.C1(n_4562),
.C2(n_4570),
.Y(n_4577)
);

AOI21xp5_ASAP7_75t_L g4578 ( 
.A1(n_4573),
.A2(n_4565),
.B(n_4564),
.Y(n_4578)
);

AOI21xp33_ASAP7_75t_L g4579 ( 
.A1(n_4572),
.A2(n_4564),
.B(n_797),
.Y(n_4579)
);

AOI222xp33_ASAP7_75t_L g4580 ( 
.A1(n_4571),
.A2(n_800),
.B1(n_802),
.B2(n_798),
.C1(n_799),
.C2(n_801),
.Y(n_4580)
);

HB1xp67_ASAP7_75t_L g4581 ( 
.A(n_4578),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4577),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4582),
.B(n_4579),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_4583),
.A2(n_4581),
.B(n_4580),
.Y(n_4584)
);

AOI211xp5_ASAP7_75t_L g4585 ( 
.A1(n_4584),
.A2(n_803),
.B(n_798),
.C(n_800),
.Y(n_4585)
);


endmodule