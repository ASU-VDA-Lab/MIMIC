module fake_jpeg_26061_n_294 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_25),
.B1(n_30),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_26),
.B1(n_18),
.B2(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_33),
.A2(n_20),
.B(n_28),
.C(n_16),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_35),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_48),
.B(n_35),
.Y(n_90)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_73),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_36),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_35),
.C(n_38),
.Y(n_110)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_25),
.B1(n_34),
.B2(n_30),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_60),
.B1(n_51),
.B2(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx2_ASAP7_75t_SL g88 ( 
.A(n_74),
.Y(n_88)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_78),
.Y(n_98)
);

OAI22x1_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_72),
.B1(n_27),
.B2(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_30),
.B1(n_24),
.B2(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_60),
.B1(n_42),
.B2(n_17),
.Y(n_92)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_100),
.B1(n_104),
.B2(n_83),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_86),
.B(n_69),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_97),
.B1(n_111),
.B2(n_82),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_103),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_60),
.B1(n_24),
.B2(n_21),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_55),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_44),
.B1(n_50),
.B2(n_61),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_79),
.Y(n_107)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_53),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_120),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_112),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_118),
.B(n_119),
.Y(n_140)
);

XOR2x1_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_67),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_75),
.B1(n_71),
.B2(n_63),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_123),
.B1(n_106),
.B2(n_101),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_90),
.A2(n_65),
.B1(n_63),
.B2(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_127),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_37),
.C(n_38),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_131),
.B(n_136),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_38),
.C(n_64),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_69),
.B1(n_45),
.B2(n_41),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_106),
.B1(n_101),
.B2(n_108),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_41),
.C(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_41),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_0),
.B(n_2),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_95),
.B(n_16),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_136),
.B(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_147),
.B(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_156),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_102),
.B1(n_99),
.B2(n_94),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_102),
.B1(n_99),
.B2(n_94),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_19),
.Y(n_156)
);

AOI21x1_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_27),
.B(n_112),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_166),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_113),
.B(n_22),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_117),
.B(n_124),
.CI(n_134),
.CON(n_160),
.SN(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_114),
.A2(n_105),
.B1(n_109),
.B2(n_18),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_167),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_26),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_26),
.A3(n_18),
.B1(n_29),
.B2(n_41),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_109),
.B1(n_29),
.B2(n_27),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_177),
.B(n_167),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_181),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_131),
.B(n_133),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_126),
.C(n_133),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_183),
.C(n_185),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_117),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_185),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_120),
.C(n_127),
.Y(n_183)
);

AOI22x1_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_118),
.B1(n_115),
.B2(n_135),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_149),
.B1(n_31),
.B2(n_3),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_115),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_115),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_190),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_189),
.B(n_192),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_125),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_109),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_166),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_194),
.B(n_197),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_148),
.C(n_157),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_198),
.B(n_206),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_142),
.C(n_140),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_204),
.C(n_211),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_177),
.A2(n_160),
.B(n_143),
.C(n_152),
.D(n_142),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_155),
.B1(n_154),
.B2(n_145),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_143),
.C(n_147),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_168),
.B(n_164),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_141),
.B1(n_153),
.B2(n_151),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_149),
.C(n_135),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_171),
.B1(n_187),
.B2(n_170),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_31),
.B1(n_10),
.B2(n_11),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_15),
.C(n_9),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_182),
.C(n_174),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g217 ( 
.A(n_201),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_220),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_215),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_186),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_184),
.B(n_176),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_208),
.B(n_187),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_191),
.B1(n_190),
.B2(n_207),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_196),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_233),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_242),
.B1(n_231),
.B2(n_2),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_232),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_223),
.Y(n_251)
);

XOR2x1_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_174),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_239),
.A2(n_11),
.B(n_6),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_195),
.C(n_196),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_246),
.C(n_218),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_171),
.B1(n_204),
.B2(n_199),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_219),
.B1(n_226),
.B2(n_207),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_222),
.C(n_221),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_253),
.C(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_225),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_224),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_6),
.C(n_7),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_239),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_256),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_244),
.B1(n_240),
.B2(n_4),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_10),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_260),
.B(n_15),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_4),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_248),
.CI(n_243),
.CON(n_266),
.SN(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_270),
.B1(n_9),
.B2(n_12),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_247),
.B(n_246),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_268),
.A2(n_269),
.B(n_9),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_235),
.B(n_241),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_249),
.B(n_12),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_264),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_281),
.B(n_13),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_262),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_274),
.B1(n_271),
.B2(n_266),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_14),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_15),
.B(n_13),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_288),
.B(n_280),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_282),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_285),
.C(n_14),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_14),
.Y(n_294)
);


endmodule