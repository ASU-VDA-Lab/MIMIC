module fake_netlist_5_935_n_1177 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1177);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1177;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_1161;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_525;
wire n_493;
wire n_397;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_1157;
wire n_1099;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_173;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_212;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_568;
wire n_936;
wire n_947;
wire n_373;
wire n_820;
wire n_1090;
wire n_757;
wire n_509;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_929;
wire n_981;
wire n_941;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_1104;
wire n_792;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_1163;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1172;
wire n_976;
wire n_1095;
wire n_1096;
wire n_234;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_1009;
wire n_1148;
wire n_264;
wire n_742;
wire n_472;
wire n_669;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_1149;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1073;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_962;
wire n_436;
wire n_181;
wire n_930;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_974;
wire n_432;
wire n_553;
wire n_395;
wire n_727;
wire n_901;
wire n_839;
wire n_311;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_328;
wire n_214;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_928;
wire n_749;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_1164;
wire n_630;
wire n_420;
wire n_632;
wire n_699;
wire n_489;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_874;
wire n_1058;
wire n_838;
wire n_358;
wire n_465;
wire n_362;
wire n_876;
wire n_170;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_1106;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_1052;
wire n_174;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_210;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1131;
wire n_1059;
wire n_1084;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_513;
wire n_425;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_679;
wire n_832;
wire n_695;
wire n_857;
wire n_180;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_1027;
wire n_805;
wire n_490;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_187;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_53),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_24),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_103),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_70),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_35),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_56),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_85),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_139),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_134),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_31),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_86),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_34),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_38),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_5),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_29),
.Y(n_191)
);

BUFx8_ASAP7_75t_SL g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_115),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_84),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_104),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_19),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_51),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_15),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_67),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_94),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_37),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_102),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_33),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_32),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_120),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_24),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_39),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_105),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_41),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_48),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_0),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_170),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_190),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_180),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_182),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_184),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_183),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_187),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_204),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_205),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_171),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_177),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_232),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_233),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_234),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_253),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_231),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_225),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_227),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_235),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_228),
.B(n_178),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_248),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_229),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_238),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_237),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_232),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_232),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_232),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_232),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_250),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g304 ( 
.A(n_251),
.B(n_179),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_284),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_271),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_263),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_287),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_292),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_256),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_265),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_278),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_263),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_266),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_288),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_290),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_267),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_290),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_285),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_301),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_264),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_268),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_289),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_329),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_348),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_348),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_344),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_336),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_339),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_324),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_331),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_323),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_316),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_330),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_329),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_311),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_306),
.B(n_260),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_311),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_280),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_318),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_315),
.B(n_283),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_340),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_270),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_346),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_345),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_351),
.A2(n_320),
.B1(n_347),
.B2(n_334),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_347),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_385),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_372),
.B(n_175),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_275),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_387),
.A2(n_370),
.B1(n_373),
.B2(n_369),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_363),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_175),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_386),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_365),
.Y(n_409)
);

OAI22x1_ASAP7_75t_SL g410 ( 
.A1(n_355),
.A2(n_318),
.B1(n_335),
.B2(n_306),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_367),
.B(n_272),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_289),
.Y(n_413)
);

INVx5_ASAP7_75t_L g414 ( 
.A(n_360),
.Y(n_414)
);

CKINVDCx11_ASAP7_75t_R g415 ( 
.A(n_374),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

BUFx8_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_379),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

OAI22x1_ASAP7_75t_R g420 ( 
.A1(n_375),
.A2(n_273),
.B1(n_288),
.B2(n_258),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_359),
.B(n_257),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_335),
.B1(n_257),
.B2(n_258),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_362),
.A2(n_259),
.B1(n_262),
.B2(n_296),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_379),
.B(n_298),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_299),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_358),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_371),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_372),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_369),
.A2(n_259),
.B1(n_262),
.B2(n_296),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_371),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

BUFx8_ASAP7_75t_SL g446 ( 
.A(n_374),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_351),
.B(n_302),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_351),
.B(n_297),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_351),
.B(n_297),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_384),
.B(n_224),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_351),
.B(n_305),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_372),
.B(n_305),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_358),
.A2(n_314),
.B(n_313),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_355),
.Y(n_457)
);

BUFx8_ASAP7_75t_L g458 ( 
.A(n_372),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_351),
.B(n_308),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_372),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_358),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_371),
.B(n_308),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_358),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_379),
.A2(n_224),
.B1(n_172),
.B2(n_173),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_358),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_371),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_456),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_456),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_404),
.B(n_390),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_421),
.B(n_181),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_404),
.B(n_326),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

CKINVDCx8_ASAP7_75t_R g481 ( 
.A(n_457),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_391),
.B(n_218),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_404),
.B(n_332),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_401),
.B(n_453),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_438),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_390),
.B(n_338),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_421),
.B(n_321),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_442),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_439),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_400),
.B(n_207),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_442),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_448),
.B(n_218),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_392),
.A2(n_206),
.B1(n_222),
.B2(n_196),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_449),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_398),
.B(n_188),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_400),
.B(n_207),
.Y(n_501)
);

AND3x1_ASAP7_75t_L g502 ( 
.A(n_428),
.B(n_189),
.C(n_195),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_416),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_459),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_462),
.B(n_197),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_462),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_467),
.B(n_200),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_389),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_406),
.B(n_201),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_394),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_451),
.B(n_171),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_396),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_461),
.B(n_208),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_435),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_461),
.B(n_211),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_446),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_440),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_479),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_481),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_479),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_481),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_513),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_519),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_519),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_475),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_503),
.B(n_414),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_479),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_475),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_R g534 ( 
.A(n_475),
.B(n_457),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_475),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_511),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_480),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_422),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_477),
.B(n_414),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_515),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_517),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_473),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_R g544 ( 
.A(n_482),
.B(n_418),
.Y(n_544)
);

INVx8_ASAP7_75t_L g545 ( 
.A(n_479),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_474),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_474),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_474),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_478),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_520),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_488),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_SL g553 ( 
.A(n_487),
.B(n_419),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_478),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_493),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_514),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_512),
.B(n_452),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_516),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_483),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_499),
.Y(n_560)
);

INVx11_ASAP7_75t_L g561 ( 
.A(n_485),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_540),
.A2(n_500),
.B(n_471),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_525),
.B(n_418),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_425),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_534),
.Y(n_565)
);

INVxp33_ASAP7_75t_SL g566 ( 
.A(n_534),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_557),
.A2(n_424),
.B1(n_426),
.B2(n_429),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_539),
.B(n_425),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_538),
.B(n_427),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_524),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_553),
.B(n_443),
.C(n_450),
.Y(n_571)
);

BUFx6f_ASAP7_75t_SL g572 ( 
.A(n_558),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_530),
.B(n_419),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_547),
.B(n_546),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_548),
.B(n_411),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_543),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_545),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_549),
.B(n_413),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_527),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_553),
.A2(n_466),
.B1(n_405),
.B2(n_495),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_558),
.B(n_402),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_554),
.B(n_413),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_536),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_552),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_531),
.B(n_478),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_529),
.B(n_408),
.Y(n_588)
);

AND3x1_ASAP7_75t_L g589 ( 
.A(n_542),
.B(n_428),
.C(n_432),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_550),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_535),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_555),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_533),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_R g594 ( 
.A(n_522),
.B(n_415),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_544),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_560),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_545),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_521),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_544),
.B(n_402),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_545),
.Y(n_600)
);

AOI21x1_ASAP7_75t_L g601 ( 
.A1(n_561),
.A2(n_471),
.B(n_470),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_556),
.B(n_495),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_521),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_528),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_521),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_521),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_528),
.B(n_501),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_551),
.B(n_395),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_523),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_523),
.Y(n_610)
);

AOI21x1_ASAP7_75t_L g611 ( 
.A1(n_523),
.A2(n_472),
.B(n_470),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_523),
.B(n_419),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_532),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_551),
.B(n_395),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_532),
.B(n_446),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_532),
.B(n_501),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_532),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_559),
.A2(n_429),
.B1(n_423),
.B2(n_431),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_559),
.B(n_419),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_559),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_557),
.A2(n_414),
.B1(n_408),
.B2(n_397),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_557),
.A2(n_189),
.B1(n_409),
.B2(n_403),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_557),
.B(n_412),
.Y(n_624)
);

AND3x2_ASAP7_75t_L g625 ( 
.A(n_557),
.B(n_510),
.C(n_506),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_545),
.Y(n_627)
);

OAI21xp33_ASAP7_75t_SL g628 ( 
.A1(n_557),
.A2(n_484),
.B(n_476),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_534),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_557),
.A2(n_399),
.B1(n_433),
.B2(n_445),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_537),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_534),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_524),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_524),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_557),
.B(n_416),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_524),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_534),
.B(n_408),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_545),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_537),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_540),
.B(n_433),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_538),
.Y(n_643)
);

BUFx8_ASAP7_75t_SL g644 ( 
.A(n_522),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_571),
.B(n_408),
.Y(n_645)
);

BUFx6f_ASAP7_75t_SL g646 ( 
.A(n_565),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_597),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_624),
.B(n_414),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_564),
.B(n_476),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_569),
.B(n_445),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_591),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_564),
.B(n_518),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_644),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_630),
.B(n_469),
.Y(n_654)
);

INVx6_ASAP7_75t_L g655 ( 
.A(n_597),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_593),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_616),
.B(n_482),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_579),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_592),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_636),
.B(n_484),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_599),
.A2(n_430),
.B1(n_433),
.B2(n_432),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_586),
.B(n_505),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_596),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_434),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_596),
.Y(n_665)
);

NOR2x1p5_ASAP7_75t_L g666 ( 
.A(n_575),
.B(n_434),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_581),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_566),
.B(n_625),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_597),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_581),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_574),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_580),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_633),
.B(n_482),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_563),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_599),
.A2(n_430),
.B1(n_434),
.B2(n_407),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_585),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_568),
.B(n_502),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_582),
.A2(n_430),
.B1(n_434),
.B2(n_407),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_597),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_607),
.B(n_505),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_602),
.A2(n_430),
.B1(n_407),
.B2(n_415),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_585),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_590),
.Y(n_683)
);

BUFx4f_ASAP7_75t_L g684 ( 
.A(n_587),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_587),
.B(n_494),
.Y(n_685)
);

INVx8_ASAP7_75t_L g686 ( 
.A(n_572),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_632),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_570),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_569),
.B(n_441),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_598),
.B(n_507),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_643),
.B(n_444),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_568),
.B(n_595),
.Y(n_692)
);

AND2x2_ASAP7_75t_SL g693 ( 
.A(n_638),
.B(n_420),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_567),
.B(n_447),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_631),
.B(n_518),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_576),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_578),
.B(n_584),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_620),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_589),
.B(n_458),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_563),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_610),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_618),
.B(n_468),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_625),
.B(n_507),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_615),
.B(n_468),
.Y(n_704)
);

INVxp33_ASAP7_75t_SL g705 ( 
.A(n_594),
.Y(n_705)
);

CKINVDCx8_ASAP7_75t_R g706 ( 
.A(n_619),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_SL g707 ( 
.A1(n_623),
.A2(n_463),
.B1(n_393),
.B2(n_410),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_641),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_623),
.B(n_518),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_608),
.B(n_498),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_576),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_622),
.B(n_508),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_642),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_619),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_608),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_622),
.B(n_491),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_577),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_598),
.B(n_508),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_626),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_626),
.B(n_516),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_583),
.A2(n_407),
.B1(n_516),
.B2(n_486),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_629),
.Y(n_722)
);

BUFx4f_ASAP7_75t_L g723 ( 
.A(n_642),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_642),
.Y(n_724)
);

BUFx4f_ASAP7_75t_L g725 ( 
.A(n_619),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_614),
.B(n_417),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_682),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_692),
.B(n_606),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_703),
.B(n_606),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_713),
.B(n_603),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_723),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_648),
.B(n_583),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_664),
.B(n_612),
.C(n_614),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_672),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_683),
.Y(n_735)
);

AND2x6_ASAP7_75t_L g736 ( 
.A(n_703),
.B(n_609),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_724),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_653),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_698),
.B(n_609),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_715),
.B(n_659),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_687),
.B(n_629),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_694),
.B(n_628),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_723),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_645),
.B(n_562),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_686),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_708),
.B(n_605),
.Y(n_746)
);

CKINVDCx11_ASAP7_75t_R g747 ( 
.A(n_686),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_660),
.B(n_663),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_714),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_665),
.B(n_613),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_714),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_667),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_670),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_676),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_714),
.Y(n_755)
);

OR2x2_ASAP7_75t_SL g756 ( 
.A(n_695),
.B(n_594),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_711),
.B(n_613),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_719),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_671),
.B(n_617),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_722),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_688),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_704),
.Y(n_762)
);

BUFx12f_ASAP7_75t_L g763 ( 
.A(n_700),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_697),
.B(n_617),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_696),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_657),
.B(n_604),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_710),
.A2(n_707),
.B1(n_677),
.B2(n_678),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_662),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_R g769 ( 
.A(n_668),
.B(n_573),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_686),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_712),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_662),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_706),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_660),
.B(n_634),
.Y(n_774)
);

AND2x6_ASAP7_75t_L g775 ( 
.A(n_712),
.B(n_619),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_690),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_657),
.B(n_621),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_666),
.B(n_621),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_701),
.B(n_588),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_651),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_656),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_655),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_649),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_649),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_701),
.B(n_611),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_684),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_650),
.B(n_634),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_652),
.B(n_702),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_690),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_720),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_690),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_717),
.B(n_577),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_690),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_717),
.B(n_627),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_655),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_668),
.B(n_601),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_731),
.B(n_693),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_742),
.A2(n_707),
.B1(n_681),
.B2(n_709),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_767),
.A2(n_661),
.B1(n_675),
.B2(n_699),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_788),
.B(n_689),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_771),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_780),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_680),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_771),
.B(n_674),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_767),
.A2(n_732),
.B1(n_762),
.B2(n_737),
.Y(n_805)
);

O2A1O1Ixp5_ASAP7_75t_L g806 ( 
.A1(n_796),
.A2(n_716),
.B(n_726),
.C(n_684),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_734),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_731),
.B(n_705),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_734),
.B(n_691),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_759),
.B(n_658),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_790),
.B(n_680),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_783),
.B(n_680),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_735),
.Y(n_813)
);

INVx8_ASAP7_75t_L g814 ( 
.A(n_763),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_731),
.B(n_673),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_769),
.B(n_680),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_784),
.B(n_718),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_780),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_731),
.B(n_673),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_753),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_764),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_732),
.A2(n_646),
.B1(n_572),
.B2(n_721),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_780),
.Y(n_823)
);

AND3x1_ASAP7_75t_L g824 ( 
.A(n_773),
.B(n_669),
.C(n_647),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_756),
.A2(n_646),
.B1(n_654),
.B2(n_685),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_727),
.B(n_647),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_740),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_743),
.B(n_685),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_743),
.B(n_679),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_762),
.B(n_669),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_727),
.B(n_718),
.Y(n_831)
);

BUFx5_ASAP7_75t_L g832 ( 
.A(n_775),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_733),
.A2(n_679),
.B1(n_725),
.B2(n_637),
.Y(n_833)
);

BUFx8_ASAP7_75t_L g834 ( 
.A(n_763),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_753),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_748),
.B(n_718),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_758),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_787),
.B(n_718),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_781),
.B(n_417),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_744),
.A2(n_219),
.B(n_215),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_768),
.B(n_635),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_743),
.B(n_779),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_760),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_754),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_780),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_744),
.B(n_221),
.C(n_220),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_743),
.B(n_627),
.Y(n_847)
);

NAND3xp33_ASAP7_75t_L g848 ( 
.A(n_796),
.B(n_774),
.C(n_785),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_752),
.B(n_635),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_739),
.B(n_637),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_746),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_779),
.A2(n_407),
.B1(n_510),
.B2(n_506),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_776),
.B(n_640),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_746),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_785),
.A2(n_600),
.B1(n_640),
.B2(n_497),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_772),
.B(n_639),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_773),
.A2(n_639),
.B(n_454),
.C(n_460),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_778),
.A2(n_485),
.B1(n_497),
.B2(n_455),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_772),
.B(n_0),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_745),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_761),
.B(n_1),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_728),
.B(n_1),
.Y(n_862)
);

NAND2x1_ASAP7_75t_L g863 ( 
.A(n_729),
.B(n_485),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_769),
.B(n_725),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_765),
.B(n_2),
.Y(n_865)
);

NAND2x1_ASAP7_75t_L g866 ( 
.A(n_729),
.B(n_485),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_807),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_804),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_854),
.B(n_729),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_851),
.B(n_729),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_834),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_821),
.B(n_729),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_801),
.B(n_736),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_827),
.B(n_736),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_820),
.B(n_736),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_809),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_863),
.B(n_776),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_813),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_826),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_835),
.B(n_736),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_834),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_844),
.B(n_736),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_836),
.B(n_757),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_837),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_843),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_800),
.B(n_745),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_866),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_814),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_848),
.B(n_789),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_856),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_832),
.B(n_789),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_832),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_853),
.B(n_791),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_818),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_832),
.B(n_791),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_841),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_849),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_799),
.A2(n_775),
.B1(n_747),
.B2(n_766),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_832),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_850),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_803),
.B(n_812),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_817),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_818),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_832),
.B(n_793),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_865),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_853),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_831),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_811),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_842),
.B(n_775),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_810),
.B(n_775),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_838),
.B(n_757),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_818),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_802),
.B(n_823),
.Y(n_913)
);

BUFx4f_ASAP7_75t_L g914 ( 
.A(n_894),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_878),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_901),
.A2(n_840),
.B(n_846),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_L g917 ( 
.A(n_868),
.B(n_814),
.Y(n_917)
);

AOI21xp33_ASAP7_75t_L g918 ( 
.A1(n_905),
.A2(n_833),
.B(n_806),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_898),
.A2(n_816),
.B(n_825),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_898),
.A2(n_805),
.B1(n_798),
.B2(n_822),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_905),
.A2(n_797),
.B(n_857),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_871),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_905),
.B(n_845),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_888),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_888),
.B(n_824),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_880),
.A2(n_864),
.B(n_808),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_888),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_907),
.A2(n_830),
.B(n_861),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_R g929 ( 
.A(n_871),
.B(n_738),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_908),
.B(n_902),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_872),
.B(n_860),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_SL g932 ( 
.A(n_871),
.B(n_814),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_906),
.Y(n_933)
);

BUFx8_ASAP7_75t_L g934 ( 
.A(n_881),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_909),
.B(n_770),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_909),
.B(n_770),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_880),
.A2(n_829),
.B(n_828),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_881),
.B(n_747),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_908),
.B(n_900),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_879),
.A2(n_862),
.B(n_855),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_872),
.B(n_730),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_883),
.A2(n_819),
.B(n_815),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_877),
.A2(n_859),
.B(n_852),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_876),
.A2(n_858),
.B1(n_786),
.B2(n_847),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_909),
.B(n_738),
.Y(n_945)
);

OAI21xp33_ASAP7_75t_L g946 ( 
.A1(n_874),
.A2(n_730),
.B(n_778),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_909),
.A2(n_786),
.B1(n_795),
.B2(n_782),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_900),
.B(n_896),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_881),
.B(n_786),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_874),
.A2(n_911),
.B(n_889),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_889),
.B(n_750),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_877),
.A2(n_839),
.B(n_786),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_894),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_886),
.A2(n_795),
.B1(n_782),
.B2(n_794),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_889),
.A2(n_775),
.B1(n_794),
.B2(n_792),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_910),
.B(n_777),
.Y(n_956)
);

OAI21xp33_ASAP7_75t_L g957 ( 
.A1(n_889),
.A2(n_741),
.B(n_750),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_892),
.A2(n_755),
.B(n_751),
.C(n_749),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_887),
.B(n_749),
.Y(n_959)
);

AO21x1_ASAP7_75t_L g960 ( 
.A1(n_884),
.A2(n_3),
.B(n_4),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_897),
.B(n_4),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_890),
.B(n_5),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_904),
.A2(n_497),
.B(n_485),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_884),
.B(n_6),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_892),
.A2(n_899),
.B(n_873),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_885),
.B(n_7),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_910),
.B(n_869),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_916),
.A2(n_899),
.B(n_873),
.Y(n_968)
);

AO22x1_ASAP7_75t_L g969 ( 
.A1(n_934),
.A2(n_899),
.B1(n_869),
.B2(n_894),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_921),
.A2(n_895),
.B(n_891),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_920),
.A2(n_906),
.B1(n_887),
.B2(n_893),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_962),
.B(n_961),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_930),
.B(n_885),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_919),
.A2(n_895),
.B(n_891),
.C(n_870),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_918),
.A2(n_867),
.B(n_903),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_951),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_925),
.B(n_887),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_932),
.B(n_906),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_917),
.A2(n_870),
.B1(n_893),
.B2(n_882),
.Y(n_979)
);

NAND2xp33_ASAP7_75t_L g980 ( 
.A(n_929),
.B(n_887),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_967),
.B(n_951),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_932),
.A2(n_945),
.B(n_960),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_934),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_943),
.A2(n_867),
.B(n_875),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_915),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_981),
.B(n_924),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_982),
.B(n_972),
.Y(n_987)
);

BUFx4f_ASAP7_75t_L g988 ( 
.A(n_983),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_SL g989 ( 
.A(n_971),
.B(n_922),
.C(n_938),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_985),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_976),
.B(n_924),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_975),
.A2(n_940),
.B(n_952),
.C(n_928),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_980),
.A2(n_936),
.B1(n_935),
.B2(n_949),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_977),
.A2(n_955),
.B1(n_927),
.B2(n_914),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_975),
.B(n_977),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_968),
.B(n_927),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_984),
.A2(n_966),
.B(n_964),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_978),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_969),
.A2(n_974),
.B(n_970),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_979),
.B(n_933),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_973),
.B(n_950),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_981),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_982),
.A2(n_914),
.B1(n_947),
.B2(n_953),
.Y(n_1003)
);

OAI21xp33_ASAP7_75t_L g1004 ( 
.A1(n_975),
.A2(n_957),
.B(n_946),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_983),
.B(n_954),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_983),
.Y(n_1006)
);

AOI22x1_ASAP7_75t_L g1007 ( 
.A1(n_982),
.A2(n_926),
.B1(n_965),
.B2(n_937),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_982),
.A2(n_958),
.B(n_959),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_982),
.A2(n_944),
.B1(n_942),
.B2(n_963),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_983),
.B(n_939),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_990),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_996),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1006),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_1002),
.B(n_986),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_987),
.B(n_948),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_991),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_998),
.B(n_931),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_1013),
.A2(n_1003),
.B1(n_1009),
.B2(n_995),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1012),
.B(n_1016),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_1017),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_1018),
.A2(n_992),
.B(n_1008),
.C(n_999),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1020),
.B(n_1014),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1019),
.A2(n_989),
.B1(n_1014),
.B2(n_998),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_1021),
.A2(n_1007),
.B(n_988),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1022),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1025),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1024),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_1027),
.Y(n_1028)
);

OAI222xp33_ASAP7_75t_L g1029 ( 
.A1(n_1026),
.A2(n_1023),
.B1(n_1011),
.B2(n_1015),
.C1(n_993),
.C2(n_994),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1028),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1029),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_1030),
.B(n_1011),
.Y(n_1032)
);

OA21x2_ASAP7_75t_L g1033 ( 
.A1(n_1031),
.A2(n_1010),
.B(n_997),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_1032),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1033),
.A2(n_998),
.B1(n_1005),
.B2(n_1000),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_1034),
.B(n_1032),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_1035),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1034),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_1036),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1036),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1038),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_1039),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1040),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1042),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1043),
.B(n_1033),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1044),
.B(n_1033),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_1045),
.B(n_1037),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1046),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1047),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1049),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1048),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_1050),
.B(n_1041),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1051),
.B(n_1001),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1053),
.B(n_1052),
.Y(n_1054)
);

NAND4xp75_ASAP7_75t_L g1055 ( 
.A(n_1052),
.B(n_9),
.C(n_7),
.D(n_8),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1053),
.B(n_1000),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_1054),
.A2(n_1004),
.B(n_12),
.C(n_10),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1056),
.A2(n_173),
.B1(n_174),
.B2(n_172),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1055),
.B(n_10),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1059),
.B(n_11),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1058),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1060),
.B(n_1057),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1061),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1062),
.B(n_1063),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1062),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_L g1066 ( 
.A(n_1064),
.B(n_176),
.C(n_174),
.Y(n_1066)
);

OAI311xp33_ASAP7_75t_L g1067 ( 
.A1(n_1065),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.C1(n_15),
.Y(n_1067)
);

AOI32xp33_ASAP7_75t_L g1068 ( 
.A1(n_1067),
.A2(n_176),
.A3(n_214),
.B1(n_202),
.B2(n_209),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1066),
.B(n_923),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1069),
.Y(n_1070)
);

NAND3xp33_ASAP7_75t_SL g1071 ( 
.A(n_1068),
.B(n_214),
.C(n_210),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1070),
.B(n_13),
.Y(n_1072)
);

AOI221xp5_ASAP7_75t_L g1073 ( 
.A1(n_1071),
.A2(n_199),
.B1(n_212),
.B2(n_213),
.C(n_217),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_1070),
.A2(n_217),
.B(n_14),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1072),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1073),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_16),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1075),
.B(n_16),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1077),
.B(n_17),
.Y(n_1079)
);

AOI322xp5_ASAP7_75t_L g1080 ( 
.A1(n_1079),
.A2(n_1076),
.A3(n_217),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_22),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1078),
.A2(n_17),
.B(n_18),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1081),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1080),
.A2(n_18),
.B(n_20),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1082),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1083),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_1084),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1085),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_SL g1088 ( 
.A1(n_1087),
.A2(n_21),
.B(n_22),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_1086),
.B(n_23),
.Y(n_1089)
);

NAND4xp25_ASAP7_75t_SL g1090 ( 
.A(n_1088),
.B(n_23),
.C(n_25),
.D(n_26),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1089),
.Y(n_1091)
);

OAI211xp5_ASAP7_75t_L g1092 ( 
.A1(n_1088),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1091),
.Y(n_1093)
);

NAND4xp25_ASAP7_75t_SL g1094 ( 
.A(n_1092),
.B(n_27),
.C(n_28),
.D(n_29),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_1090),
.Y(n_1095)
);

AOI221xp5_ASAP7_75t_SL g1096 ( 
.A1(n_1093),
.A2(n_28),
.B1(n_30),
.B2(n_337),
.C(n_40),
.Y(n_1096)
);

NOR2x1_ASAP7_75t_L g1097 ( 
.A(n_1095),
.B(n_337),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1097),
.B(n_1094),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1096),
.B(n_30),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_1098),
.B(n_36),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1101),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_1100),
.B(n_894),
.Y(n_1103)
);

NOR2x1_ASAP7_75t_L g1104 ( 
.A(n_1102),
.B(n_337),
.Y(n_1104)
);

OA22x2_ASAP7_75t_L g1105 ( 
.A1(n_1103),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1104),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_1105),
.B(n_45),
.C(n_46),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1106),
.B(n_47),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1107),
.A2(n_337),
.B1(n_497),
.B2(n_455),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1106),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1110),
.B(n_49),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1109),
.B(n_50),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_1108),
.B(n_52),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1113),
.A2(n_337),
.B1(n_497),
.B2(n_894),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_SL g1116 ( 
.A1(n_1114),
.A2(n_1115),
.B1(n_1111),
.B2(n_57),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1114),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1117),
.A2(n_912),
.B1(n_894),
.B2(n_486),
.Y(n_1118)
);

XNOR2xp5_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_54),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1119),
.A2(n_912),
.B1(n_448),
.B2(n_486),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1118),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1121),
.A2(n_912),
.B1(n_903),
.B2(n_465),
.Y(n_1122)
);

NAND4xp75_ASAP7_75t_L g1123 ( 
.A(n_1120),
.B(n_55),
.C(n_58),
.D(n_59),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1122),
.B(n_60),
.Y(n_1124)
);

OAI22x1_ASAP7_75t_L g1125 ( 
.A1(n_1123),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1124),
.B(n_64),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_1125),
.B(n_912),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_SL g1128 ( 
.A1(n_1124),
.A2(n_912),
.B1(n_66),
.B2(n_68),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1124),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_912),
.B1(n_465),
.B2(n_489),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1127),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1126),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1128),
.A2(n_509),
.B1(n_504),
.B2(n_496),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1133),
.B(n_1130),
.Y(n_1134)
);

AOI221x1_ASAP7_75t_L g1135 ( 
.A1(n_1132),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.C(n_79),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1131),
.B(n_483),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_SL g1137 ( 
.A1(n_1134),
.A2(n_80),
.B(n_81),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1136),
.B(n_82),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1135),
.A2(n_83),
.B(n_88),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1134),
.A2(n_489),
.B1(n_504),
.B2(n_496),
.Y(n_1140)
);

OA21x2_ASAP7_75t_L g1141 ( 
.A1(n_1134),
.A2(n_89),
.B(n_90),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1134),
.B(n_91),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1134),
.B(n_92),
.Y(n_1143)
);

XNOR2xp5_ASAP7_75t_L g1144 ( 
.A(n_1134),
.B(n_93),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1134),
.Y(n_1145)
);

INVxp33_ASAP7_75t_L g1146 ( 
.A(n_1134),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1134),
.A2(n_95),
.B(n_96),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1134),
.B(n_97),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1145),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_SL g1150 ( 
.A1(n_1146),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1139),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1138),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1137),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1144),
.A2(n_489),
.B1(n_490),
.B2(n_483),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1143),
.A2(n_101),
.B1(n_106),
.B2(n_107),
.C(n_109),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1148),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1142),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1149),
.A2(n_1141),
.B1(n_1147),
.B2(n_1140),
.Y(n_1158)
);

AOI222xp33_ASAP7_75t_SL g1159 ( 
.A1(n_1157),
.A2(n_1141),
.B1(n_111),
.B2(n_113),
.C1(n_114),
.C2(n_116),
.Y(n_1159)
);

AOI222xp33_ASAP7_75t_L g1160 ( 
.A1(n_1153),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.C1(n_121),
.C2(n_122),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1151),
.A2(n_124),
.B(n_125),
.Y(n_1161)
);

AOI222xp33_ASAP7_75t_L g1162 ( 
.A1(n_1156),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.C1(n_130),
.C2(n_131),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1152),
.A2(n_483),
.B1(n_490),
.B2(n_492),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_R g1164 ( 
.A1(n_1154),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_R g1165 ( 
.A1(n_1158),
.A2(n_1150),
.B1(n_1155),
.B2(n_141),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1159),
.B(n_490),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1161),
.B(n_138),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1164),
.A2(n_1160),
.B(n_1162),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1168),
.A2(n_1163),
.B1(n_913),
.B2(n_144),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1166),
.A2(n_913),
.B1(n_142),
.B2(n_145),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1169),
.A2(n_1165),
.B1(n_1167),
.B2(n_147),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1171),
.A2(n_1170),
.B(n_146),
.Y(n_1172)
);

OAI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1172),
.A2(n_140),
.B1(n_149),
.B2(n_150),
.C(n_152),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1173),
.A2(n_153),
.B(n_154),
.C(n_155),
.Y(n_1174)
);

AOI21xp33_ASAP7_75t_L g1175 ( 
.A1(n_1174),
.A2(n_157),
.B(n_158),
.Y(n_1175)
);

AOI211xp5_ASAP7_75t_L g1176 ( 
.A1(n_1175),
.A2(n_956),
.B(n_160),
.C(n_161),
.Y(n_1176)
);

AOI211xp5_ASAP7_75t_L g1177 ( 
.A1(n_1176),
.A2(n_941),
.B(n_164),
.C(n_166),
.Y(n_1177)
);


endmodule