module fake_jpeg_24596_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_30),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_20),
.A2(n_32),
.B1(n_16),
.B2(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_36),
.B(n_37),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_66),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_14),
.C(n_10),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_79),
.B(n_29),
.Y(n_111)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_67),
.Y(n_114)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_36),
.CI(n_26),
.CON(n_79),
.SN(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_29),
.Y(n_80)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_80),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_43),
.B1(n_39),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_41),
.B1(n_38),
.B2(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_26),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_44),
.B1(n_20),
.B2(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_43),
.B1(n_44),
.B2(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_44),
.B1(n_38),
.B2(n_43),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_19),
.B1(n_27),
.B2(n_45),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_20),
.B1(n_16),
.B2(n_32),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_42),
.B(n_35),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_36),
.C(n_37),
.Y(n_98)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_60),
.B1(n_42),
.B2(n_35),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_96),
.B1(n_109),
.B2(n_123),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_97),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_45),
.B(n_31),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_99),
.A2(n_108),
.B1(n_113),
.B2(n_45),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_100),
.A2(n_31),
.B1(n_21),
.B2(n_45),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_36),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_120),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_20),
.B1(n_16),
.B2(n_32),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_42),
.B1(n_35),
.B2(n_26),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_26),
.B1(n_19),
.B2(n_36),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_36),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_90),
.B1(n_91),
.B2(n_77),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_140),
.B1(n_151),
.B2(n_152),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_25),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_129),
.B(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_78),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_64),
.B1(n_89),
.B2(n_83),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_137),
.B1(n_139),
.B2(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_141),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_92),
.B1(n_73),
.B2(n_70),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_72),
.B1(n_67),
.B2(n_69),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_28),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_21),
.B1(n_31),
.B2(n_27),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_140),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_150),
.B1(n_25),
.B2(n_23),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_25),
.B1(n_23),
.B2(n_28),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_24),
.B1(n_17),
.B2(n_33),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_110),
.CI(n_100),
.CON(n_157),
.SN(n_157)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_157),
.B(n_159),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_169),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_117),
.B1(n_107),
.B2(n_102),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_163),
.B1(n_34),
.B2(n_33),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_170),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_100),
.B1(n_117),
.B2(n_107),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_102),
.B(n_118),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_172),
.B(n_143),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_28),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_17),
.B(n_24),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_185),
.B(n_33),
.Y(n_218)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_177),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_116),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_179),
.Y(n_207)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_182),
.B1(n_164),
.B2(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_112),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_18),
.Y(n_182)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_34),
.C(n_33),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_34),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_128),
.B(n_18),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_215),
.B1(n_216),
.B2(n_165),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_190),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_135),
.B(n_137),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_192),
.A2(n_194),
.B(n_204),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_181),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_193),
.B(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_132),
.C(n_149),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_201),
.C(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_103),
.B1(n_115),
.B2(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_197),
.A2(n_199),
.B1(n_208),
.B2(n_212),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_161),
.B1(n_172),
.B2(n_153),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_202),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_103),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_33),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_0),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_23),
.B(n_129),
.C(n_17),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_205),
.B(n_9),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_115),
.B1(n_74),
.B2(n_24),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_0),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_177),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_157),
.A2(n_127),
.B1(n_148),
.B2(n_34),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_148),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_127),
.C(n_34),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_159),
.C(n_180),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_1),
.B(n_2),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_156),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_22),
.B(n_2),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_222),
.B1(n_199),
.B2(n_208),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_168),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_217),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_229),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_239),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_165),
.B1(n_171),
.B2(n_169),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_232),
.A2(n_212),
.B1(n_209),
.B2(n_194),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_197),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_238),
.C(n_243),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_22),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_22),
.C(n_2),
.Y(n_238)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_215),
.B(n_200),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_22),
.C(n_3),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_22),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_214),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_204),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_249),
.B(n_260),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_206),
.B(n_192),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_203),
.B(n_233),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_228),
.B1(n_243),
.B2(n_222),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_223),
.B(n_218),
.C(n_210),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_221),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_188),
.B1(n_192),
.B2(n_205),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_210),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_262),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_240),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_238),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_241),
.B1(n_234),
.B2(n_226),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_273),
.B1(n_266),
.B2(n_267),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_219),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_272),
.C(n_276),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_219),
.C(n_235),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_232),
.B1(n_230),
.B2(n_244),
.Y(n_274)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_253),
.C(n_252),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_242),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_277),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_279),
.A2(n_280),
.B(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_225),
.C(n_236),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_281),
.A2(n_255),
.B1(n_252),
.B2(n_245),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_247),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_286),
.B(n_272),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_255),
.B1(n_254),
.B2(n_249),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_293),
.B1(n_281),
.B2(n_276),
.Y(n_298)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_1),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_10),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_271),
.A2(n_254),
.B1(n_259),
.B2(n_251),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_258),
.B1(n_248),
.B2(n_257),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_263),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_257),
.B1(n_204),
.B2(n_5),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_268),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_299),
.B(n_308),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_280),
.B1(n_282),
.B2(n_270),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_300),
.A2(n_287),
.B1(n_284),
.B2(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_304),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_305),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_289),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_15),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_294),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_307),
.A2(n_285),
.B(n_295),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_300),
.C(n_298),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_284),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_304),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_321),
.B(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_317),
.B(n_295),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_314),
.B1(n_311),
.B2(n_318),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_327),
.B(n_319),
.Y(n_328)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

A2O1A1O1Ixp25_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_325),
.B(n_11),
.C(n_12),
.D(n_7),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_12),
.B(n_5),
.C(n_6),
.Y(n_330)
);

A2O1A1O1Ixp25_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_4),
.B(n_6),
.C(n_7),
.D(n_313),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_4),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_4),
.B(n_6),
.Y(n_333)
);


endmodule