module real_jpeg_26654_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_60),
.Y(n_104)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_1),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_27),
.B1(n_92),
.B2(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_2),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_2),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_68),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_24),
.B(n_76),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_94),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_5),
.A2(n_51),
.B(n_66),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_5),
.A2(n_86),
.B1(n_161),
.B2(n_162),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_7),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_153)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_71),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_12),
.Y(n_88)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_15),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_115),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_113),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_19),
.B(n_81),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.C(n_73),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_20),
.A2(n_21),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_22),
.B(n_41),
.C(n_47),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_33),
.B2(n_38),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_23),
.A2(n_28),
.B1(n_33),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_44),
.Y(n_90)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_25),
.A2(n_35),
.A3(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_25),
.A2(n_90),
.B1(n_91),
.B2(n_95),
.Y(n_89)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_28),
.A2(n_33),
.B1(n_38),
.B2(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_30),
.B(n_36),
.Y(n_77)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_33),
.Y(n_143)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_36),
.A2(n_64),
.B(n_94),
.C(n_138),
.Y(n_137)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_43),
.A2(n_91),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_43),
.A2(n_44),
.B(n_92),
.C(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_92),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B(n_55),
.Y(n_47)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_49),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_57),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_51),
.B1(n_64),
.B2(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_50),
.B(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_56),
.A2(n_57),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_57),
.B(n_79),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_61),
.B(n_73),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B(n_69),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_65),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_62),
.A2(n_65),
.B1(n_125),
.B2(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_65),
.B(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_78),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_98),
.B1(n_99),
.B2(n_112),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_96),
.B2(n_97),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_86),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_86),
.A2(n_153),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

HAxp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.CON(n_91),
.SN(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_94),
.B(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_101),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_129),
.B(n_176),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_117),
.B(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_123),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_118),
.A2(n_119),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_170),
.B(n_175),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_149),
.B(n_169),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_132),
.B(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_145),
.C(n_146),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_157),
.B(n_168),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_155),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_163),
.B(n_167),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_172),
.Y(n_175)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);


endmodule