module fake_ariane_1067_n_2154 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_478, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_496, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2154);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_478;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2154;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_552;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_1467;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_519;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_504;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_523;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_162),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_433),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_349),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_406),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_157),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_45),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_57),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_465),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_67),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_41),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_140),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_340),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_255),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_473),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_487),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_145),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_188),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_362),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_86),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_482),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_499),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_436),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_422),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_483),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_402),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_208),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_480),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_485),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_156),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_491),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_157),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_430),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_249),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_42),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_51),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_77),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_179),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_345),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_63),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_5),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_212),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_88),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_301),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_171),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_213),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_136),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_67),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_474),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_459),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_496),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_371),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_404),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_41),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_262),
.Y(n_558)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_250),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_118),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_469),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_51),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_445),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_369),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_373),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_64),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_111),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_381),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_438),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_222),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_128),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_394),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_114),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_77),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_376),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_463),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_87),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_46),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_27),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_429),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_98),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_233),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_165),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_83),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_440),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_479),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_234),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_336),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_494),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_154),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_320),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_167),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_448),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_28),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_458),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_300),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_197),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_481),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_107),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_195),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_261),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_352),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_71),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_248),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_237),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_121),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_285),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_235),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_162),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_401),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_175),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_384),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_72),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_23),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_61),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_447),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_15),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_1),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_39),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_461),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_42),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_15),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_410),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_492),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_414),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_164),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_420),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_450),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_309),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_444),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_168),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_190),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_271),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_12),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_318),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_392),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_27),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_428),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_382),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_191),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_454),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_146),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_403),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_385),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_89),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_71),
.Y(n_646)
);

CKINVDCx14_ASAP7_75t_R g647 ( 
.A(n_417),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_342),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_434),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_238),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_423),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_311),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_327),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_216),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_399),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_302),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_61),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_103),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_493),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_446),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_231),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_164),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_9),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_475),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_471),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_432),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_466),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_435),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_144),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_395),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_33),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_419),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_326),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_180),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_37),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_253),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_105),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_40),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_143),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_337),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_135),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_462),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_284),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_477),
.Y(n_684)
);

CKINVDCx16_ASAP7_75t_R g685 ( 
.A(n_425),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_363),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_490),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_36),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_441),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_113),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_43),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_443),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_484),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_437),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_380),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_196),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_415),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_14),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_431),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_17),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_78),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_274),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_53),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_193),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_409),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_28),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_101),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_476),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_372),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_66),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_79),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_411),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_89),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_453),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_56),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_177),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_81),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_85),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_30),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_87),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_128),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_449),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_100),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_292),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_106),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_20),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_442),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_460),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_272),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_0),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_468),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_91),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_159),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_424),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_102),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_228),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_353),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_102),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_146),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_148),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_260),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_185),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_151),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_364),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_452),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_456),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_478),
.Y(n_747)
);

CKINVDCx14_ASAP7_75t_R g748 ( 
.A(n_464),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_105),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_472),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_343),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_451),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_298),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_488),
.Y(n_754)
);

BUFx2_ASAP7_75t_SL g755 ( 
.A(n_69),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_467),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_457),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_94),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_280),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_426),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_270),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_316),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_348),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_68),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_40),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_470),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_427),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_215),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_149),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_93),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_158),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_205),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_542),
.Y(n_773)
);

CKINVDCx16_ASAP7_75t_R g774 ( 
.A(n_540),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_542),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_597),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_615),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_615),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_534),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_543),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_701),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_669),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_545),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_574),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_616),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_577),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_666),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_579),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_556),
.Y(n_789)
);

INVxp33_ASAP7_75t_SL g790 ( 
.A(n_755),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_583),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_696),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_594),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_737),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_599),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_619),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_556),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_642),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_663),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_677),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_678),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_691),
.Y(n_802)
);

INVx4_ASAP7_75t_R g803 ( 
.A(n_591),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_621),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_700),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_717),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_720),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_723),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_732),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_594),
.Y(n_810)
);

INVxp67_ASAP7_75t_SL g811 ( 
.A(n_621),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_735),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_738),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_645),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_740),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_556),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_594),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_594),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_657),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_645),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_764),
.Y(n_821)
);

INVxp67_ASAP7_75t_SL g822 ( 
.A(n_671),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_771),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_671),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_749),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_749),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_532),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_761),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_562),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_657),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_768),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_657),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_657),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_538),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_504),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_707),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_707),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_500),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_707),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_707),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_610),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_715),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_505),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_743),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_726),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_708),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_517),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_517),
.Y(n_848)
);

INVxp67_ASAP7_75t_SL g849 ( 
.A(n_614),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_506),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_509),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_656),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_656),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_692),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_516),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_692),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_716),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_508),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_716),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_510),
.Y(n_860)
);

CKINVDCx14_ASAP7_75t_R g861 ( 
.A(n_559),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_591),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_847),
.B(n_561),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_776),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_781),
.A2(n_662),
.B1(n_613),
.B2(n_685),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_861),
.B(n_501),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_862),
.B(n_766),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_789),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_787),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_789),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_848),
.B(n_766),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_789),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_777),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_838),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_774),
.B(n_647),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_852),
.B(n_521),
.Y(n_877)
);

CKINVDCx11_ASAP7_75t_R g878 ( 
.A(n_835),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_793),
.Y(n_879)
);

CKINVDCx6p67_ASAP7_75t_R g880 ( 
.A(n_785),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_779),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_827),
.B(n_748),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_797),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_810),
.A2(n_515),
.B(n_511),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_817),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_797),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_797),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_780),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_782),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_850),
.Y(n_890)
);

OA21x2_ASAP7_75t_L g891 ( 
.A1(n_832),
.A2(n_523),
.B(n_522),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_816),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_816),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_853),
.B(n_611),
.Y(n_895)
);

OAI22x1_ASAP7_75t_L g896 ( 
.A1(n_845),
.A2(n_646),
.B1(n_679),
.B2(n_622),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_783),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_782),
.A2(n_719),
.B1(n_578),
.B2(n_675),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_816),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_820),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_819),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_830),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_784),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_833),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_836),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_837),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_786),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_839),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_794),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_840),
.Y(n_910)
);

OA21x2_ASAP7_75t_L g911 ( 
.A1(n_824),
.A2(n_530),
.B(n_526),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_845),
.A2(n_551),
.B1(n_560),
.B2(n_539),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_788),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_791),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_820),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_773),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_795),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_854),
.B(n_856),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_825),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_775),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_796),
.Y(n_921)
);

AND2x6_ASAP7_75t_L g922 ( 
.A(n_857),
.B(n_611),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_778),
.Y(n_923)
);

BUFx12f_ASAP7_75t_L g924 ( 
.A(n_831),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_829),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_881),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_878),
.Y(n_927)
);

INVxp33_ASAP7_75t_L g928 ( 
.A(n_871),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_919),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_868),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_888),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_R g932 ( 
.A(n_890),
.B(n_790),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_897),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_864),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_869),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_868),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_909),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_878),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_903),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_924),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_875),
.B(n_851),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_880),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_919),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_919),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_907),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_913),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_914),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_871),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_889),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_889),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_917),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_900),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_919),
.Y(n_953)
);

CKINVDCx6p67_ASAP7_75t_R g954 ( 
.A(n_876),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_904),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_904),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_916),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_916),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_900),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_915),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_921),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_905),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_882),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_915),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_905),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_920),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_R g967 ( 
.A(n_920),
.B(n_855),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_875),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_865),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_863),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_863),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_912),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_918),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_923),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_925),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_923),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_877),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_877),
.B(n_546),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_925),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_866),
.B(n_792),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_898),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_906),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_874),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_872),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_872),
.B(n_859),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_911),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_901),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_895),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_895),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_896),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_922),
.B(n_843),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_867),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_911),
.Y(n_993)
);

AO21x2_ASAP7_75t_L g994 ( 
.A1(n_884),
.A2(n_549),
.B(n_547),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_922),
.B(n_828),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_911),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_906),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_906),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_867),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_901),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_867),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_867),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_867),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_906),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_922),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_908),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_908),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_908),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_908),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_SL g1010 ( 
.A(n_934),
.B(n_858),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_987),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_929),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_964),
.B(n_827),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_963),
.A2(n_922),
.B1(n_841),
.B2(n_846),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_937),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_1004),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_973),
.B(n_922),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_970),
.B(n_860),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_963),
.B(n_804),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_985),
.B(n_804),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_926),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_929),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_975),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_1006),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_949),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_985),
.B(n_811),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_935),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_931),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_933),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_979),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_941),
.B(n_520),
.Y(n_1031)
);

INVx4_ASAP7_75t_SL g1032 ( 
.A(n_974),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_SL g1033 ( 
.A(n_940),
.B(n_968),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_955),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_929),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_977),
.B(n_849),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_952),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_939),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_950),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_956),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1000),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_957),
.B(n_849),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_993),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_962),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_993),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_959),
.B(n_928),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_959),
.B(n_834),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_1007),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_942),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_929),
.Y(n_1050)
);

BUFx10_ASAP7_75t_L g1051 ( 
.A(n_971),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_957),
.B(n_879),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_981),
.A2(n_891),
.B1(n_910),
.B2(n_668),
.Y(n_1053)
);

CKINVDCx8_ASAP7_75t_R g1054 ( 
.A(n_948),
.Y(n_1054)
);

OR2x2_ASAP7_75t_SL g1055 ( 
.A(n_932),
.B(n_798),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_986),
.A2(n_891),
.B1(n_910),
.B2(n_668),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_943),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_945),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_960),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_972),
.B(n_537),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_965),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_L g1062 ( 
.A(n_932),
.B(n_842),
.C(n_834),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_984),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_1009),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_946),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_991),
.A2(n_891),
.B(n_887),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_930),
.Y(n_1067)
);

INVx6_ASAP7_75t_L g1068 ( 
.A(n_998),
.Y(n_1068)
);

NAND2xp33_ASAP7_75t_R g1069 ( 
.A(n_995),
.B(n_844),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_988),
.B(n_842),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_947),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_930),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_936),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_951),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_961),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_969),
.B(n_811),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_958),
.B(n_879),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_976),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_936),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_989),
.B(n_814),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_967),
.B(n_814),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_927),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_958),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_967),
.B(n_550),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_1008),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_1008),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_978),
.A2(n_566),
.B(n_557),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_966),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_995),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_966),
.B(n_885),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_998),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_998),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_944),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_953),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_954),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_978),
.B(n_567),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_998),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_982),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_938),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_997),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_999),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1005),
.B(n_885),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_983),
.B(n_571),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_992),
.Y(n_1104)
);

BUFx10_ASAP7_75t_L g1105 ( 
.A(n_1001),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_992),
.B(n_799),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1002),
.B(n_893),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1003),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_994),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_994),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_980),
.B(n_573),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_996),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_980),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_990),
.Y(n_1114)
);

AND2x4_ASAP7_75t_SL g1115 ( 
.A(n_954),
.B(n_726),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_964),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_935),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_975),
.Y(n_1118)
);

AND2x6_ASAP7_75t_L g1119 ( 
.A(n_991),
.B(n_512),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_941),
.B(n_581),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_987),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_973),
.B(n_893),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_975),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_935),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_964),
.B(n_822),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_929),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_987),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1004),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_929),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_949),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_987),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_970),
.B(n_584),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_970),
.B(n_590),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_964),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_935),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_987),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_975),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_968),
.Y(n_1138)
);

OA22x2_ASAP7_75t_L g1139 ( 
.A1(n_964),
.A2(n_801),
.B1(n_802),
.B2(n_800),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_964),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_964),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_973),
.B(n_902),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_1141),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1060),
.A2(n_826),
.B1(n_822),
.B2(n_603),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1027),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1021),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1034),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1081),
.B(n_826),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1036),
.B(n_902),
.Y(n_1149)
);

AO22x2_ASAP7_75t_L g1150 ( 
.A1(n_1112),
.A2(n_805),
.B1(n_807),
.B2(n_806),
.Y(n_1150)
);

OAI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1132),
.A2(n_609),
.B1(n_617),
.B2(n_606),
.C(n_592),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1116),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1117),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1028),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1134),
.B(n_618),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1040),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1133),
.A2(n_552),
.B1(n_572),
.B2(n_570),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1013),
.B(n_808),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1029),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_SL g1160 ( 
.A(n_1015),
.B(n_513),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1125),
.B(n_809),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1019),
.B(n_626),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1019),
.B(n_1042),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1032),
.B(n_812),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_1140),
.Y(n_1165)
);

AO22x2_ASAP7_75t_L g1166 ( 
.A1(n_1076),
.A2(n_815),
.B1(n_821),
.B2(n_813),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1044),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1020),
.B(n_634),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1038),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1058),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1065),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_1138),
.B(n_823),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1022),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1061),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1018),
.B(n_637),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1096),
.A2(n_681),
.B1(n_688),
.B2(n_658),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1037),
.B(n_690),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_1032),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1039),
.B(n_698),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1054),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_1095),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1020),
.B(n_703),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_1124),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1071),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1074),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1026),
.B(n_706),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1135),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1023),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1059),
.B(n_710),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1030),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1046),
.B(n_711),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1106),
.B(n_575),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1010),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1139),
.A2(n_718),
.B1(n_721),
.B2(n_713),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1118),
.Y(n_1195)
);

INVxp33_ASAP7_75t_SL g1196 ( 
.A(n_1033),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1123),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1075),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_L g1199 ( 
.A(n_1017),
.B(n_725),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1137),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1011),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1106),
.A2(n_596),
.B1(n_604),
.B2(n_582),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1049),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1082),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1016),
.B(n_730),
.Y(n_1205)
);

AND2x6_ASAP7_75t_L g1206 ( 
.A(n_1043),
.B(n_512),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1103),
.B(n_733),
.Y(n_1207)
);

BUFx8_ASAP7_75t_L g1208 ( 
.A(n_1025),
.Y(n_1208)
);

NAND2x1p5_ASAP7_75t_L g1209 ( 
.A(n_1095),
.B(n_873),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1011),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1041),
.Y(n_1211)
);

AND2x2_ASAP7_75t_SL g1212 ( 
.A(n_1089),
.B(n_529),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1041),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1016),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1121),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1121),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1127),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1127),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1026),
.B(n_739),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1131),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1131),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1022),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1024),
.A2(n_620),
.B1(n_629),
.B2(n_607),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_1130),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1080),
.B(n_758),
.Y(n_1225)
);

AO22x2_ASAP7_75t_L g1226 ( 
.A1(n_1114),
.A2(n_555),
.B1(n_563),
.B2(n_529),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1136),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1136),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1047),
.B(n_765),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1070),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1057),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1063),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1024),
.B(n_769),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1078),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1052),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1048),
.B(n_873),
.Y(n_1236)
);

CKINVDCx11_ASAP7_75t_R g1237 ( 
.A(n_1051),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1077),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1057),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1090),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1048),
.B(n_887),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1093),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1094),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1100),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1083),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1064),
.B(n_1128),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1088),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1099),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1067),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1055),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1072),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1073),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1051),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1079),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1064),
.B(n_770),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1128),
.B(n_502),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1098),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1087),
.A2(n_633),
.B(n_636),
.C(n_632),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1043),
.B(n_531),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1085),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1122),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1085),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1142),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1105),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1086),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_L g1266 ( 
.A(n_1062),
.B(n_639),
.C(n_638),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1113),
.B(n_585),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1108),
.B(n_1115),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1108),
.B(n_894),
.Y(n_1269)
);

NAND3xp33_ASAP7_75t_L g1270 ( 
.A(n_1014),
.B(n_643),
.C(n_641),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1084),
.B(n_625),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1086),
.Y(n_1272)
);

AO22x2_ASAP7_75t_L g1273 ( 
.A1(n_1045),
.A2(n_555),
.B1(n_744),
.B2(n_563),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1097),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1045),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1012),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1069),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1012),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1105),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1108),
.B(n_644),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1104),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1102),
.Y(n_1282)
);

OR2x4_ASAP7_75t_L g1283 ( 
.A(n_1031),
.B(n_651),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1120),
.B(n_654),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1107),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1126),
.Y(n_1286)
);

NAND2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1101),
.B(n_894),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1126),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1101),
.B(n_1119),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1022),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1111),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1035),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1068),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1068),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1035),
.B(n_655),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1035),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1053),
.B(n_1056),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1050),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_SL g1299 ( 
.A(n_1119),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1050),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1119),
.B(n_757),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1050),
.B(n_503),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1091),
.B(n_659),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1091),
.B(n_507),
.Y(n_1304)
);

NAND2x1p5_ASAP7_75t_L g1305 ( 
.A(n_1091),
.B(n_661),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1092),
.B(n_673),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1092),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1119),
.B(n_683),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1129),
.B(n_686),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1092),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1129),
.A2(n_689),
.B1(n_697),
.B2(n_687),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1109),
.Y(n_1312)
);

NAND2x1p5_ASAP7_75t_L g1313 ( 
.A(n_1129),
.B(n_705),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1066),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1110),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1021),
.Y(n_1316)
);

AO22x2_ASAP7_75t_L g1317 ( 
.A1(n_1112),
.A2(n_762),
.B1(n_744),
.B2(n_714),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1034),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1021),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1081),
.A2(n_742),
.B1(n_753),
.B2(n_709),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1021),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1095),
.B(n_760),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1021),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1081),
.B(n_763),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1016),
.B(n_514),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1021),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1032),
.B(n_533),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1021),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1022),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1034),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1116),
.B(n_518),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1021),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1013),
.B(n_0),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1178),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1207),
.B(n_519),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1314),
.A2(n_762),
.B(n_631),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1199),
.A2(n_525),
.B(n_524),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1148),
.B(n_1),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1235),
.A2(n_528),
.B(n_527),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1163),
.B(n_1161),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1196),
.B(n_535),
.Y(n_1342)
);

OAI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1175),
.A2(n_1177),
.B(n_1176),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1238),
.A2(n_541),
.B(n_536),
.Y(n_1344)
);

AOI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1289),
.A2(n_883),
.B(n_870),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1301),
.A2(n_1308),
.B(n_1309),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1158),
.B(n_2),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1240),
.A2(n_548),
.B(n_544),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1157),
.A2(n_554),
.B(n_558),
.C(n_553),
.Y(n_1349)
);

AO22x1_ASAP7_75t_L g1350 ( 
.A1(n_1208),
.A2(n_564),
.B1(n_568),
.B2(n_565),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1211),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1201),
.A2(n_1215),
.B(n_1210),
.Y(n_1352)
);

CKINVDCx16_ASAP7_75t_R g1353 ( 
.A(n_1248),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_L g1354 ( 
.A(n_1160),
.B(n_1284),
.C(n_1151),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1183),
.B(n_569),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1152),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1216),
.A2(n_883),
.B(n_870),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_SL g1358 ( 
.A(n_1180),
.B(n_576),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1218),
.A2(n_586),
.B(n_580),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1275),
.A2(n_588),
.B(n_587),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1285),
.A2(n_589),
.B(n_595),
.C(n_593),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1281),
.A2(n_600),
.B(n_598),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1261),
.B(n_2),
.Y(n_1363)
);

O2A1O1Ixp5_ASAP7_75t_L g1364 ( 
.A1(n_1302),
.A2(n_803),
.B(n_5),
.C(n_3),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1271),
.A2(n_601),
.B(n_605),
.C(n_602),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1146),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1221),
.A2(n_883),
.B(n_870),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1178),
.Y(n_1368)
);

AOI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1227),
.A2(n_883),
.B(n_870),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1263),
.B(n_1333),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1230),
.B(n_3),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1324),
.B(n_4),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1143),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_SL g1374 ( 
.A(n_1208),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1212),
.B(n_608),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1228),
.A2(n_612),
.B(n_624),
.C(n_623),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1155),
.B(n_627),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1246),
.B(n_4),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1231),
.A2(n_892),
.B(n_886),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1260),
.A2(n_630),
.B(n_628),
.Y(n_1380)
);

NOR2xp67_ASAP7_75t_L g1381 ( 
.A(n_1165),
.B(n_635),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1154),
.A2(n_640),
.B1(n_649),
.B2(n_648),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1181),
.B(n_650),
.Y(n_1383)
);

AND2x6_ASAP7_75t_L g1384 ( 
.A(n_1297),
.B(n_556),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1262),
.A2(n_653),
.B(n_652),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1277),
.B(n_6),
.Y(n_1386)
);

AOI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1239),
.A2(n_1288),
.B(n_1286),
.Y(n_1387)
);

OAI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1179),
.A2(n_664),
.B(n_660),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1265),
.A2(n_670),
.B(n_665),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1272),
.A2(n_674),
.B(n_672),
.Y(n_1390)
);

AOI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1213),
.A2(n_892),
.B(n_886),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1232),
.B(n_676),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1246),
.B(n_6),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1145),
.B(n_886),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1282),
.B(n_7),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1229),
.B(n_7),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1189),
.A2(n_680),
.B1(n_684),
.B2(n_682),
.Y(n_1397)
);

AOI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1217),
.A2(n_892),
.B(n_886),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1153),
.B(n_693),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1220),
.A2(n_695),
.B(n_694),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1276),
.A2(n_702),
.B(n_699),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1225),
.B(n_8),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1188),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1258),
.A2(n_704),
.B(n_722),
.C(n_712),
.Y(n_1404)
);

NOR2x1_ASAP7_75t_L g1405 ( 
.A(n_1181),
.B(n_892),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1332),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1204),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1166),
.B(n_8),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1278),
.A2(n_727),
.B(n_724),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1259),
.A2(n_729),
.B(n_728),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1245),
.A2(n_734),
.B(n_731),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1247),
.A2(n_741),
.B(n_736),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1233),
.A2(n_746),
.B(n_745),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1331),
.B(n_747),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1224),
.B(n_667),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1298),
.A2(n_899),
.B(n_772),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1255),
.A2(n_751),
.B(n_750),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1149),
.A2(n_754),
.B(n_752),
.Y(n_1418)
);

OAI21xp33_ASAP7_75t_L g1419 ( 
.A1(n_1144),
.A2(n_759),
.B(n_756),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1268),
.B(n_9),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1251),
.A2(n_767),
.B(n_10),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1267),
.B(n_10),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1159),
.B(n_11),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1169),
.B(n_11),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1252),
.A2(n_12),
.B(n_13),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1268),
.B(n_13),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1187),
.B(n_899),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1304),
.A2(n_772),
.B(n_667),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1256),
.A2(n_772),
.B(n_667),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1325),
.A2(n_1307),
.B(n_1171),
.Y(n_1430)
);

AO21x1_ASAP7_75t_L g1431 ( 
.A1(n_1303),
.A2(n_772),
.B(n_667),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_1250),
.Y(n_1432)
);

AO21x1_ASAP7_75t_L g1433 ( 
.A1(n_1295),
.A2(n_170),
.B(n_169),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1170),
.A2(n_899),
.B(n_173),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1184),
.A2(n_899),
.B(n_174),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1185),
.A2(n_176),
.B(n_172),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1190),
.Y(n_1437)
);

AO32x1_ASAP7_75t_L g1438 ( 
.A1(n_1311),
.A2(n_17),
.A3(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1254),
.A2(n_16),
.B(n_18),
.Y(n_1439)
);

OAI21xp33_ASAP7_75t_L g1440 ( 
.A1(n_1191),
.A2(n_19),
.B(n_20),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1166),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1198),
.A2(n_181),
.B(n_178),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1249),
.A2(n_21),
.B(n_22),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1223),
.A2(n_23),
.B(n_24),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1316),
.A2(n_183),
.B(n_182),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1250),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1172),
.B(n_24),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1319),
.B(n_1321),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1164),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1193),
.B(n_25),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1323),
.A2(n_186),
.B(n_184),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1291),
.B(n_25),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1326),
.B(n_1328),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1237),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1290),
.A2(n_189),
.B(n_187),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1164),
.B(n_26),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1150),
.B(n_26),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1320),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_1458)
);

NOR2xp67_ASAP7_75t_L g1459 ( 
.A(n_1264),
.B(n_1214),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1292),
.A2(n_194),
.B(n_192),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1234),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1173),
.Y(n_1462)
);

INVx4_ASAP7_75t_L g1463 ( 
.A(n_1253),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1209),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1295),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1296),
.A2(n_199),
.B(n_198),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1206),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1269),
.A2(n_201),
.B(n_200),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1310),
.A2(n_203),
.B(n_202),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1242),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1243),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1205),
.A2(n_206),
.B(n_204),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1274),
.A2(n_1300),
.B(n_1222),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1300),
.A2(n_209),
.B(n_207),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1173),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1192),
.B(n_32),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1202),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1266),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1244),
.A2(n_37),
.B(n_38),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1194),
.B(n_38),
.C(n_39),
.Y(n_1480)
);

AOI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1273),
.A2(n_211),
.B(n_210),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1173),
.A2(n_217),
.B(n_214),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1222),
.A2(n_219),
.B(n_218),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1222),
.A2(n_221),
.B(n_220),
.Y(n_1484)
);

BUFx8_ASAP7_75t_L g1485 ( 
.A(n_1299),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_L g1486 ( 
.A(n_1279),
.B(n_43),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_SL g1487 ( 
.A(n_1322),
.B(n_44),
.C(n_45),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1195),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1197),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1329),
.A2(n_224),
.B(n_223),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1192),
.B(n_44),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1280),
.B(n_46),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1280),
.B(n_47),
.Y(n_1493)
);

BUFx8_ASAP7_75t_L g1494 ( 
.A(n_1327),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1206),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1329),
.A2(n_226),
.B(n_225),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1329),
.Y(n_1497)
);

NAND2x1p5_ASAP7_75t_L g1498 ( 
.A(n_1294),
.B(n_227),
.Y(n_1498)
);

O2A1O1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1162),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1168),
.B(n_50),
.Y(n_1500)
);

NOR2xp67_ASAP7_75t_L g1501 ( 
.A(n_1182),
.B(n_229),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1150),
.B(n_52),
.Y(n_1502)
);

AOI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1273),
.A2(n_1306),
.B(n_1257),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1293),
.A2(n_1312),
.B(n_1287),
.Y(n_1504)
);

AO21x1_ASAP7_75t_L g1505 ( 
.A1(n_1306),
.A2(n_232),
.B(n_230),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1327),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1200),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1186),
.A2(n_239),
.B(n_236),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1270),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1509)
);

NOR2x1p5_ASAP7_75t_SL g1510 ( 
.A(n_1147),
.B(n_240),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1305),
.A2(n_242),
.B(n_241),
.Y(n_1511)
);

AOI21xp33_ASAP7_75t_L g1512 ( 
.A1(n_1219),
.A2(n_54),
.B(n_55),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1156),
.A2(n_55),
.B(n_56),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1283),
.B(n_57),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1315),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1167),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1174),
.A2(n_58),
.B(n_59),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1318),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1330),
.A2(n_244),
.B(n_243),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1206),
.B(n_58),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1315),
.A2(n_246),
.B(n_245),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1236),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1408),
.B(n_1317),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1356),
.B(n_1313),
.Y(n_1524)
);

AOI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1345),
.A2(n_1226),
.B(n_1317),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1351),
.Y(n_1526)
);

O2A1O1Ixp5_ASAP7_75t_L g1527 ( 
.A1(n_1335),
.A2(n_1241),
.B(n_1226),
.C(n_1315),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_SL g1528 ( 
.A(n_1343),
.B(n_59),
.C(n_60),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1403),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1354),
.B(n_60),
.Y(n_1530)
);

O2A1O1Ixp5_ASAP7_75t_L g1531 ( 
.A1(n_1414),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1377),
.A2(n_62),
.B(n_65),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1366),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1500),
.A2(n_68),
.B(n_65),
.C(n_66),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1406),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1422),
.A2(n_72),
.B(n_69),
.C(n_70),
.Y(n_1536)
);

INVx6_ASAP7_75t_L g1537 ( 
.A(n_1494),
.Y(n_1537)
);

INVx4_ASAP7_75t_L g1538 ( 
.A(n_1353),
.Y(n_1538)
);

O2A1O1Ixp5_ASAP7_75t_L g1539 ( 
.A1(n_1421),
.A2(n_74),
.B(n_70),
.C(n_73),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1357),
.A2(n_251),
.B(n_247),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1461),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1334),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1373),
.B(n_73),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1352),
.A2(n_254),
.B(n_252),
.Y(n_1544)
);

OR2x6_ASAP7_75t_SL g1545 ( 
.A(n_1454),
.B(n_74),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1370),
.B(n_75),
.Y(n_1546)
);

INVx4_ASAP7_75t_L g1547 ( 
.A(n_1334),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1448),
.A2(n_257),
.B(n_256),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1334),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1437),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1449),
.B(n_498),
.Y(n_1551)
);

AND2x2_ASAP7_75t_SL g1552 ( 
.A(n_1441),
.B(n_75),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1340),
.B(n_76),
.Y(n_1553)
);

BUFx2_ASAP7_75t_SL g1554 ( 
.A(n_1341),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1378),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_1555)
);

A2O1A1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1440),
.A2(n_1444),
.B(n_1372),
.C(n_1480),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1432),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1358),
.B(n_80),
.Y(n_1558)
);

AO21x1_ASAP7_75t_L g1559 ( 
.A1(n_1513),
.A2(n_1517),
.B(n_1443),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1453),
.A2(n_259),
.B(n_258),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1378),
.B(n_1393),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1488),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1489),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1507),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1486),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1393),
.B(n_82),
.Y(n_1566)
);

A2O1A1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1375),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_SL g1568 ( 
.A(n_1463),
.B(n_84),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1436),
.A2(n_264),
.B(n_263),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1470),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1506),
.B(n_86),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1420),
.B(n_88),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1458),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1407),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1442),
.A2(n_266),
.B(n_265),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1518),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1445),
.A2(n_268),
.B(n_267),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1388),
.A2(n_93),
.B(n_90),
.C(n_92),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1471),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1396),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1402),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1450),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1368),
.B(n_1497),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1497),
.B(n_99),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1451),
.A2(n_273),
.B(n_269),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_SL g1586 ( 
.A(n_1487),
.B(n_1477),
.C(n_1399),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1423),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1465),
.B(n_100),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1420),
.B(n_101),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1452),
.A2(n_106),
.B1(n_103),
.B2(n_104),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1347),
.B(n_104),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1516),
.B(n_107),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1446),
.B(n_108),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1387),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1497),
.B(n_108),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1479),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1426),
.B(n_109),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1426),
.B(n_110),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1485),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1424),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1462),
.B(n_112),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_R g1602 ( 
.A(n_1374),
.B(n_275),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1494),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1515),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1395),
.B(n_112),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1492),
.B(n_113),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1338),
.B(n_114),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1493),
.B(n_115),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1430),
.A2(n_277),
.B(n_276),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1368),
.B(n_278),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1508),
.A2(n_281),
.B(n_279),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1450),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1434),
.A2(n_283),
.B(n_282),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1368),
.B(n_116),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1386),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1522),
.B(n_497),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1342),
.B(n_117),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1435),
.A2(n_287),
.B(n_286),
.Y(n_1618)
);

AOI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1474),
.A2(n_289),
.B(n_288),
.Y(n_1619)
);

XNOR2xp5_ASAP7_75t_L g1620 ( 
.A(n_1350),
.B(n_118),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1457),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1502),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_SL g1623 ( 
.A(n_1485),
.B(n_290),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1363),
.B(n_119),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1462),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1476),
.B(n_119),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1467),
.B(n_120),
.C(n_121),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1478),
.A2(n_123),
.B(n_120),
.C(n_122),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1464),
.B(n_291),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_SL g1630 ( 
.A1(n_1361),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1425),
.A2(n_294),
.B(n_293),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1371),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1491),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1515),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1397),
.B(n_124),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1439),
.A2(n_296),
.B(n_295),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1462),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1475),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1360),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1429),
.A2(n_299),
.B(n_297),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1362),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1475),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1519),
.A2(n_304),
.B(n_303),
.Y(n_1643)
);

AOI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1472),
.A2(n_306),
.B(n_305),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1456),
.B(n_129),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1520),
.Y(n_1646)
);

INVxp67_ASAP7_75t_SL g1647 ( 
.A(n_1515),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1459),
.B(n_495),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1365),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_1649)
);

O2A1O1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1512),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_1650)
);

AO221x2_ASAP7_75t_L g1651 ( 
.A1(n_1438),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.C(n_135),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1475),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1499),
.A2(n_136),
.B(n_133),
.C(n_134),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1447),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1504),
.B(n_137),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1427),
.A2(n_308),
.B(n_307),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_SL g1657 ( 
.A1(n_1433),
.A2(n_1505),
.B(n_1481),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1415),
.B(n_137),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1455),
.A2(n_312),
.B(n_310),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1509),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1349),
.A2(n_141),
.B(n_138),
.C(n_139),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1415),
.B(n_141),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1514),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1392),
.Y(n_1664)
);

O2A1O1Ixp33_ASAP7_75t_SL g1665 ( 
.A1(n_1376),
.A2(n_142),
.B(n_145),
.C(n_147),
.Y(n_1665)
);

AND2x6_ASAP7_75t_L g1666 ( 
.A(n_1495),
.B(n_313),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1460),
.A2(n_315),
.B(n_314),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1382),
.B(n_147),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1466),
.A2(n_1469),
.B(n_1418),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1501),
.B(n_148),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1404),
.A2(n_149),
.B(n_150),
.C(n_151),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1381),
.B(n_150),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1473),
.A2(n_319),
.B(n_317),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1394),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1428),
.A2(n_322),
.B(n_321),
.Y(n_1675)
);

AO21x2_ASAP7_75t_L g1676 ( 
.A1(n_1336),
.A2(n_324),
.B(n_323),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1355),
.B(n_152),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1346),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1503),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1542),
.Y(n_1680)
);

INVx6_ASAP7_75t_L g1681 ( 
.A(n_1537),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1583),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1533),
.Y(n_1683)
);

INVx4_ASAP7_75t_L g1684 ( 
.A(n_1537),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1603),
.Y(n_1685)
);

INVx5_ASAP7_75t_L g1686 ( 
.A(n_1542),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1599),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1574),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1561),
.B(n_152),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1633),
.B(n_1384),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1538),
.B(n_1583),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1597),
.B(n_1383),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1557),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1554),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1572),
.B(n_153),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1549),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1549),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1679),
.Y(n_1698)
);

BUFx4f_ASAP7_75t_L g1699 ( 
.A(n_1614),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1652),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1523),
.B(n_1384),
.Y(n_1701)
);

NAND2x1p5_ASAP7_75t_L g1702 ( 
.A(n_1547),
.B(n_1405),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1587),
.B(n_1384),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1535),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1625),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1589),
.B(n_153),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1526),
.Y(n_1707)
);

BUFx4f_ASAP7_75t_SL g1708 ( 
.A(n_1652),
.Y(n_1708)
);

INVx8_ASAP7_75t_L g1709 ( 
.A(n_1614),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1541),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1566),
.B(n_1419),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1678),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1524),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1570),
.Y(n_1714)
);

BUFx2_ASAP7_75t_SL g1715 ( 
.A(n_1666),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1579),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1638),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1621),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1564),
.Y(n_1719)
);

INVxp67_ASAP7_75t_SL g1720 ( 
.A(n_1646),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1622),
.Y(n_1721)
);

INVx3_ASAP7_75t_SL g1722 ( 
.A(n_1662),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1552),
.A2(n_1384),
.B1(n_1400),
.B2(n_1339),
.Y(n_1723)
);

CKINVDCx20_ASAP7_75t_R g1724 ( 
.A(n_1602),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1616),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1642),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1616),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1604),
.Y(n_1728)
);

INVx5_ASAP7_75t_L g1729 ( 
.A(n_1662),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1576),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1529),
.Y(n_1731)
);

INVx6_ASAP7_75t_L g1732 ( 
.A(n_1637),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1546),
.Y(n_1733)
);

NAND2x1p5_ASAP7_75t_L g1734 ( 
.A(n_1551),
.B(n_1511),
.Y(n_1734)
);

BUFx4_ASAP7_75t_SL g1735 ( 
.A(n_1632),
.Y(n_1735)
);

CKINVDCx14_ASAP7_75t_R g1736 ( 
.A(n_1545),
.Y(n_1736)
);

OR2x6_ASAP7_75t_L g1737 ( 
.A(n_1629),
.B(n_1498),
.Y(n_1737)
);

INVx5_ASAP7_75t_L g1738 ( 
.A(n_1666),
.Y(n_1738)
);

INVx1_ASAP7_75t_SL g1739 ( 
.A(n_1598),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1664),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1648),
.Y(n_1741)
);

INVx6_ASAP7_75t_SL g1742 ( 
.A(n_1648),
.Y(n_1742)
);

CKINVDCx20_ASAP7_75t_R g1743 ( 
.A(n_1620),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1550),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1543),
.B(n_154),
.Y(n_1745)
);

INVx3_ASAP7_75t_SL g1746 ( 
.A(n_1610),
.Y(n_1746)
);

BUFx2_ASAP7_75t_SL g1747 ( 
.A(n_1610),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1593),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1562),
.Y(n_1749)
);

BUFx12f_ASAP7_75t_L g1750 ( 
.A(n_1551),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1634),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1674),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1674),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1563),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1674),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1592),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1588),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1600),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1654),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1658),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1571),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1635),
.A2(n_1344),
.B1(n_1348),
.B2(n_1359),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1668),
.Y(n_1763)
);

BUFx2_ASAP7_75t_SL g1764 ( 
.A(n_1666),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1672),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1615),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1594),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1553),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1607),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1626),
.Y(n_1770)
);

BUFx4f_ASAP7_75t_L g1771 ( 
.A(n_1623),
.Y(n_1771)
);

INVx4_ASAP7_75t_L g1772 ( 
.A(n_1676),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1647),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1606),
.B(n_1411),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1584),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1558),
.B(n_155),
.Y(n_1776)
);

INVx3_ASAP7_75t_SL g1777 ( 
.A(n_1595),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1591),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1525),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1530),
.Y(n_1780)
);

BUFx8_ASAP7_75t_L g1781 ( 
.A(n_1582),
.Y(n_1781)
);

BUFx12f_ASAP7_75t_L g1782 ( 
.A(n_1612),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1605),
.Y(n_1783)
);

NAND2x1p5_ASAP7_75t_L g1784 ( 
.A(n_1655),
.B(n_1468),
.Y(n_1784)
);

INVx6_ASAP7_75t_L g1785 ( 
.A(n_1617),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1540),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1677),
.B(n_1413),
.Y(n_1787)
);

AO21x1_ASAP7_75t_L g1788 ( 
.A1(n_1532),
.A2(n_1521),
.B(n_1483),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1624),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1608),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1528),
.A2(n_1412),
.B1(n_1409),
.B2(n_1401),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1531),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1527),
.Y(n_1793)
);

BUFx5_ASAP7_75t_L g1794 ( 
.A(n_1673),
.Y(n_1794)
);

INVx4_ASAP7_75t_L g1795 ( 
.A(n_1568),
.Y(n_1795)
);

BUFx2_ASAP7_75t_SL g1796 ( 
.A(n_1601),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1738),
.A2(n_1590),
.B1(n_1567),
.B2(n_1534),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1787),
.A2(n_1565),
.B(n_1596),
.C(n_1556),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1683),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1689),
.B(n_1645),
.Y(n_1800)
);

AO21x2_ASAP7_75t_L g1801 ( 
.A1(n_1793),
.A2(n_1657),
.B(n_1431),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1738),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1681),
.Y(n_1803)
);

OAI21x1_ASAP7_75t_L g1804 ( 
.A1(n_1779),
.A2(n_1369),
.B(n_1367),
.Y(n_1804)
);

OR2x6_ASAP7_75t_L g1805 ( 
.A(n_1715),
.B(n_1631),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1719),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1715),
.A2(n_1651),
.B1(n_1663),
.B2(n_1627),
.Y(n_1807)
);

NAND2x1p5_ASAP7_75t_L g1808 ( 
.A(n_1771),
.B(n_1670),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1711),
.A2(n_1636),
.B(n_1539),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1704),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1693),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1774),
.A2(n_1578),
.B(n_1641),
.Y(n_1812)
);

NAND2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1699),
.B(n_1482),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1784),
.A2(n_1416),
.B(n_1398),
.Y(n_1814)
);

OR3x4_ASAP7_75t_SL g1815 ( 
.A(n_1736),
.B(n_1651),
.C(n_155),
.Y(n_1815)
);

NAND3xp33_ASAP7_75t_L g1816 ( 
.A(n_1738),
.B(n_1536),
.C(n_1639),
.Y(n_1816)
);

NOR2xp67_ASAP7_75t_R g1817 ( 
.A(n_1795),
.B(n_1559),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1730),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1710),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1714),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1716),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1707),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1761),
.B(n_1555),
.Y(n_1823)
);

OAI21x1_ASAP7_75t_L g1824 ( 
.A1(n_1734),
.A2(n_1391),
.B(n_1379),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1764),
.A2(n_1573),
.B(n_1586),
.C(n_1661),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1720),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1766),
.B(n_1580),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1782),
.A2(n_1581),
.B1(n_1649),
.B2(n_1653),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1792),
.A2(n_1669),
.B(n_1611),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1726),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1758),
.B(n_1718),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1694),
.B(n_156),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1723),
.A2(n_1660),
.B(n_1628),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1718),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1740),
.B(n_158),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1788),
.A2(n_1544),
.B(n_1619),
.Y(n_1836)
);

AO21x2_ASAP7_75t_L g1837 ( 
.A1(n_1703),
.A2(n_1609),
.B(n_1643),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1773),
.B(n_1510),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1778),
.A2(n_1671),
.B(n_1650),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1686),
.B(n_1484),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1731),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1721),
.Y(n_1842)
);

NOR2xp67_ASAP7_75t_L g1843 ( 
.A(n_1772),
.B(n_1548),
.Y(n_1843)
);

AOI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1786),
.A2(n_1560),
.B(n_1644),
.Y(n_1844)
);

OAI21x1_ASAP7_75t_L g1845 ( 
.A1(n_1690),
.A2(n_1618),
.B(n_1613),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1786),
.A2(n_1575),
.B(n_1569),
.Y(n_1846)
);

OAI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1759),
.A2(n_1585),
.B(n_1577),
.Y(n_1847)
);

OAI21x1_ASAP7_75t_L g1848 ( 
.A1(n_1767),
.A2(n_1667),
.B(n_1659),
.Y(n_1848)
);

OAI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1702),
.A2(n_1640),
.B(n_1675),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1721),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1763),
.B(n_1665),
.Y(n_1851)
);

AO32x2_ASAP7_75t_L g1852 ( 
.A1(n_1725),
.A2(n_1438),
.A3(n_1630),
.B1(n_1364),
.B2(n_163),
.Y(n_1852)
);

OAI21x1_ASAP7_75t_L g1853 ( 
.A1(n_1769),
.A2(n_1656),
.B(n_1496),
.Y(n_1853)
);

AO21x2_ASAP7_75t_L g1854 ( 
.A1(n_1701),
.A2(n_1417),
.B(n_1410),
.Y(n_1854)
);

INVx3_ASAP7_75t_L g1855 ( 
.A(n_1741),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1681),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1698),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1791),
.A2(n_1490),
.B(n_1385),
.Y(n_1858)
);

OA21x2_ASAP7_75t_L g1859 ( 
.A1(n_1712),
.A2(n_1389),
.B(n_1380),
.Y(n_1859)
);

OAI21x1_ASAP7_75t_L g1860 ( 
.A1(n_1768),
.A2(n_1749),
.B(n_1744),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1698),
.Y(n_1861)
);

OAI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1754),
.A2(n_1390),
.B(n_1337),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1733),
.B(n_159),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1712),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1783),
.A2(n_328),
.B(n_325),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1685),
.B(n_160),
.Y(n_1866)
);

OAI21x1_ASAP7_75t_L g1867 ( 
.A1(n_1836),
.A2(n_1682),
.B(n_1789),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1830),
.Y(n_1868)
);

CKINVDCx8_ASAP7_75t_R g1869 ( 
.A(n_1815),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1831),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1806),
.Y(n_1871)
);

OA21x2_ASAP7_75t_L g1872 ( 
.A1(n_1829),
.A2(n_1762),
.B(n_1770),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1807),
.A2(n_1764),
.B1(n_1785),
.B2(n_1790),
.Y(n_1873)
);

BUFx4f_ASAP7_75t_SL g1874 ( 
.A(n_1803),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1797),
.A2(n_1729),
.B1(n_1747),
.B2(n_1785),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1818),
.Y(n_1876)
);

BUFx3_ASAP7_75t_L g1877 ( 
.A(n_1856),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1860),
.Y(n_1878)
);

INVx2_ASAP7_75t_SL g1879 ( 
.A(n_1857),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1811),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1834),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1799),
.Y(n_1882)
);

CKINVDCx11_ASAP7_75t_R g1883 ( 
.A(n_1805),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1850),
.B(n_1826),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1810),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1819),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1820),
.Y(n_1887)
);

OA21x2_ASAP7_75t_L g1888 ( 
.A1(n_1846),
.A2(n_1748),
.B(n_1776),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1821),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1864),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1822),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1805),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1842),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1841),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1861),
.B(n_1757),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1838),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1838),
.Y(n_1897)
);

AOI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1809),
.A2(n_1780),
.B(n_1739),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1828),
.A2(n_1777),
.B1(n_1796),
.B2(n_1729),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1797),
.A2(n_1816),
.B1(n_1828),
.B2(n_1833),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1801),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1801),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1827),
.Y(n_1903)
);

AO21x2_ASAP7_75t_L g1904 ( 
.A1(n_1809),
.A2(n_1692),
.B(n_1745),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1804),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1903),
.B(n_1800),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1900),
.A2(n_1798),
.B(n_1805),
.Y(n_1907)
);

NOR3xp33_ASAP7_75t_SL g1908 ( 
.A(n_1880),
.B(n_1835),
.C(n_1825),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1868),
.B(n_1823),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1877),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1869),
.A2(n_1816),
.B1(n_1833),
.B2(n_1839),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1893),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1903),
.B(n_1817),
.Y(n_1913)
);

CKINVDCx16_ASAP7_75t_R g1914 ( 
.A(n_1877),
.Y(n_1914)
);

CKINVDCx16_ASAP7_75t_R g1915 ( 
.A(n_1868),
.Y(n_1915)
);

OR2x6_ASAP7_75t_L g1916 ( 
.A(n_1888),
.B(n_1802),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1886),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1870),
.B(n_1817),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1879),
.B(n_1688),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1874),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_R g1921 ( 
.A(n_1880),
.B(n_1724),
.Y(n_1921)
);

NOR2x1_ASAP7_75t_R g1922 ( 
.A(n_1883),
.B(n_1684),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1871),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1871),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1886),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1879),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1881),
.B(n_1802),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1890),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1890),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1896),
.B(n_1855),
.Y(n_1930)
);

NOR2x1_ASAP7_75t_L g1931 ( 
.A(n_1913),
.B(n_1904),
.Y(n_1931)
);

INVxp67_ASAP7_75t_L g1932 ( 
.A(n_1918),
.Y(n_1932)
);

INVx3_ASAP7_75t_L g1933 ( 
.A(n_1910),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1915),
.B(n_1892),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1910),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1926),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1926),
.B(n_1892),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1917),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1909),
.B(n_1892),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1925),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1916),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_SL g1942 ( 
.A1(n_1911),
.A2(n_1888),
.B(n_1904),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1916),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1928),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1906),
.B(n_1884),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1911),
.A2(n_1904),
.B1(n_1812),
.B2(n_1765),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1929),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1938),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1946),
.A2(n_1888),
.B1(n_1907),
.B2(n_1899),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1940),
.Y(n_1950)
);

NOR2xp67_ASAP7_75t_L g1951 ( 
.A(n_1936),
.B(n_1920),
.Y(n_1951)
);

OA21x2_ASAP7_75t_L g1952 ( 
.A1(n_1941),
.A2(n_1912),
.B(n_1902),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1932),
.A2(n_1869),
.B1(n_1908),
.B2(n_1914),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1944),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1934),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1949),
.B(n_1942),
.C(n_1931),
.Y(n_1956)
);

INVx4_ASAP7_75t_L g1957 ( 
.A(n_1955),
.Y(n_1957)
);

AOI221xp5_ASAP7_75t_L g1958 ( 
.A1(n_1953),
.A2(n_1942),
.B1(n_1873),
.B2(n_1839),
.C(n_1812),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1954),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1948),
.B(n_1945),
.Y(n_1960)
);

AOI221xp5_ASAP7_75t_L g1961 ( 
.A1(n_1956),
.A2(n_1832),
.B1(n_1898),
.B2(n_1950),
.C(n_1943),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1959),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1957),
.B(n_1951),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1960),
.B(n_1933),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1958),
.B(n_1945),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1960),
.B(n_1947),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1963),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1962),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1964),
.B(n_1934),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1968),
.B(n_1965),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1967),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1971),
.Y(n_1972)
);

O2A1O1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1970),
.B(n_1967),
.C(n_1866),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1973),
.B(n_1969),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1973),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1975),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1974),
.Y(n_1977)
);

NAND3xp33_ASAP7_75t_L g1978 ( 
.A(n_1977),
.B(n_1781),
.C(n_1961),
.Y(n_1978)
);

NOR3xp33_ASAP7_75t_L g1979 ( 
.A(n_1976),
.B(n_1687),
.C(n_1863),
.Y(n_1979)
);

NOR2xp67_ASAP7_75t_L g1980 ( 
.A(n_1977),
.B(n_1969),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1980),
.A2(n_1969),
.B(n_1966),
.Y(n_1981)
);

NAND2xp33_ASAP7_75t_SL g1982 ( 
.A(n_1979),
.B(n_1921),
.Y(n_1982)
);

NAND2x1_ASAP7_75t_L g1983 ( 
.A(n_1978),
.B(n_1910),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1981),
.A2(n_1729),
.B(n_1709),
.C(n_1706),
.Y(n_1984)
);

AOI211xp5_ASAP7_75t_L g1985 ( 
.A1(n_1982),
.A2(n_1722),
.B(n_1922),
.C(n_1695),
.Y(n_1985)
);

NAND3xp33_ASAP7_75t_SL g1986 ( 
.A(n_1983),
.B(n_1743),
.C(n_1808),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1981),
.Y(n_1987)
);

OAI211xp5_ASAP7_75t_L g1988 ( 
.A1(n_1981),
.A2(n_1709),
.B(n_1935),
.C(n_1933),
.Y(n_1988)
);

AOI221xp5_ASAP7_75t_L g1989 ( 
.A1(n_1981),
.A2(n_1756),
.B1(n_1765),
.B2(n_1760),
.C(n_1919),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1983),
.A2(n_1708),
.B1(n_1943),
.B2(n_1941),
.Y(n_1990)
);

AO22x1_ASAP7_75t_L g1991 ( 
.A1(n_1987),
.A2(n_1933),
.B1(n_1935),
.B2(n_1691),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1985),
.B(n_1935),
.Y(n_1992)
);

AOI211xp5_ASAP7_75t_L g1993 ( 
.A1(n_1988),
.A2(n_1756),
.B(n_1760),
.C(n_1746),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1986),
.A2(n_1952),
.B1(n_1854),
.B2(n_1937),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1984),
.Y(n_1995)
);

INVxp67_ASAP7_75t_SL g1996 ( 
.A(n_1990),
.Y(n_1996)
);

AOI22xp33_ASAP7_75t_L g1997 ( 
.A1(n_1989),
.A2(n_1952),
.B1(n_1854),
.B2(n_1916),
.Y(n_1997)
);

INVxp67_ASAP7_75t_SL g1998 ( 
.A(n_1987),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_SL g1999 ( 
.A1(n_1987),
.A2(n_1735),
.B1(n_1750),
.B2(n_1732),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1987),
.B(n_160),
.Y(n_2000)
);

NOR3xp33_ASAP7_75t_L g2001 ( 
.A(n_1998),
.B(n_1700),
.C(n_1865),
.Y(n_2001)
);

NAND4xp75_ASAP7_75t_L g2002 ( 
.A(n_2000),
.B(n_1994),
.C(n_1996),
.D(n_1995),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1991),
.B(n_1895),
.Y(n_2003)
);

CKINVDCx6p67_ASAP7_75t_R g2004 ( 
.A(n_1992),
.Y(n_2004)
);

AND4x2_ASAP7_75t_L g2005 ( 
.A(n_1992),
.B(n_165),
.C(n_161),
.D(n_163),
.Y(n_2005)
);

NOR3xp33_ASAP7_75t_SL g2006 ( 
.A(n_1999),
.B(n_161),
.C(n_166),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1993),
.A2(n_166),
.B(n_167),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1997),
.B(n_1937),
.Y(n_2008)
);

NOR4xp75_ASAP7_75t_L g2009 ( 
.A(n_1998),
.B(n_1851),
.C(n_1855),
.D(n_1939),
.Y(n_2009)
);

NAND3xp33_ASAP7_75t_L g2010 ( 
.A(n_2000),
.B(n_1705),
.C(n_1680),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_2000),
.B(n_1737),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_2000),
.Y(n_2012)
);

NAND4xp75_ASAP7_75t_L g2013 ( 
.A(n_2000),
.B(n_1697),
.C(n_1696),
.D(n_1939),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_2000),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1998),
.B(n_1713),
.Y(n_2015)
);

NAND3xp33_ASAP7_75t_L g2016 ( 
.A(n_2000),
.B(n_1680),
.C(n_1727),
.Y(n_2016)
);

A2O1A1Ixp33_ASAP7_75t_SL g2017 ( 
.A1(n_1998),
.A2(n_1905),
.B(n_331),
.C(n_329),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1998),
.A2(n_1813),
.B1(n_1737),
.B2(n_1775),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_2000),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_2000),
.Y(n_2020)
);

XOR2xp5_ASAP7_75t_L g2021 ( 
.A(n_1999),
.B(n_1727),
.Y(n_2021)
);

NAND2x1p5_ASAP7_75t_L g2022 ( 
.A(n_2000),
.B(n_1686),
.Y(n_2022)
);

NOR3xp33_ASAP7_75t_L g2023 ( 
.A(n_1998),
.B(n_1875),
.C(n_1742),
.Y(n_2023)
);

BUFx2_ASAP7_75t_L g2024 ( 
.A(n_2000),
.Y(n_2024)
);

NAND2x1p5_ASAP7_75t_L g2025 ( 
.A(n_2000),
.B(n_1686),
.Y(n_2025)
);

OAI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1998),
.A2(n_1732),
.B1(n_1775),
.B2(n_1796),
.C(n_1859),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_2024),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_2014),
.Y(n_2028)
);

CKINVDCx16_ASAP7_75t_R g2029 ( 
.A(n_2019),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_2020),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_2022),
.Y(n_2031)
);

NAND2xp33_ASAP7_75t_L g2032 ( 
.A(n_2006),
.B(n_1780),
.Y(n_2032)
);

AO22x2_ASAP7_75t_L g2033 ( 
.A1(n_2012),
.A2(n_1717),
.B1(n_1885),
.B2(n_1882),
.Y(n_2033)
);

XNOR2xp5_ASAP7_75t_L g2034 ( 
.A(n_2011),
.B(n_1742),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_2015),
.A2(n_1887),
.B1(n_1889),
.B2(n_1896),
.C(n_1897),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_2004),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2025),
.B(n_1927),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_2021),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_2007),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_2010),
.Y(n_2040)
);

CKINVDCx20_ASAP7_75t_R g2041 ( 
.A(n_2005),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2002),
.Y(n_2042)
);

BUFx4f_ASAP7_75t_L g2043 ( 
.A(n_2003),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2013),
.Y(n_2044)
);

NAND3xp33_ASAP7_75t_SL g2045 ( 
.A(n_2017),
.B(n_2023),
.C(n_2016),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_2018),
.B(n_1752),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_2008),
.Y(n_2047)
);

CKINVDCx16_ASAP7_75t_R g2048 ( 
.A(n_2009),
.Y(n_2048)
);

BUFx2_ASAP7_75t_L g2049 ( 
.A(n_2001),
.Y(n_2049)
);

CKINVDCx20_ASAP7_75t_R g2050 ( 
.A(n_2026),
.Y(n_2050)
);

CKINVDCx20_ASAP7_75t_R g2051 ( 
.A(n_2004),
.Y(n_2051)
);

NAND2x1_ASAP7_75t_SL g2052 ( 
.A(n_2014),
.B(n_1930),
.Y(n_2052)
);

AOI211x1_ASAP7_75t_SL g2053 ( 
.A1(n_2007),
.A2(n_1843),
.B(n_1901),
.C(n_1902),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_2024),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2028),
.Y(n_2055)
);

OAI22xp5_ASAP7_75t_SL g2056 ( 
.A1(n_2051),
.A2(n_1752),
.B1(n_1859),
.B2(n_1840),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2041),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2029),
.B(n_2030),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2048),
.A2(n_1883),
.B1(n_1843),
.B2(n_1872),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_2027),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2027),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_2036),
.A2(n_2042),
.B(n_2054),
.Y(n_2062)
);

AO21x2_ASAP7_75t_L g2063 ( 
.A1(n_2045),
.A2(n_1930),
.B(n_1844),
.Y(n_2063)
);

XNOR2x1_ASAP7_75t_SL g2064 ( 
.A(n_2047),
.B(n_1753),
.Y(n_2064)
);

OA22x2_ASAP7_75t_L g2065 ( 
.A1(n_2031),
.A2(n_1897),
.B1(n_1867),
.B2(n_1905),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_2054),
.A2(n_1862),
.B(n_1872),
.Y(n_2066)
);

AO21x2_ASAP7_75t_L g2067 ( 
.A1(n_2044),
.A2(n_330),
.B(n_332),
.Y(n_2067)
);

OAI22x1_ASAP7_75t_L g2068 ( 
.A1(n_2039),
.A2(n_1755),
.B1(n_1872),
.B2(n_1901),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2043),
.A2(n_1858),
.B(n_1853),
.Y(n_2069)
);

AO21x2_ASAP7_75t_L g2070 ( 
.A1(n_2032),
.A2(n_333),
.B(n_334),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2052),
.Y(n_2071)
);

AO22x2_ASAP7_75t_L g2072 ( 
.A1(n_2038),
.A2(n_1878),
.B1(n_338),
.B2(n_339),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2040),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_2049),
.Y(n_2074)
);

AO21x2_ASAP7_75t_L g2075 ( 
.A1(n_2037),
.A2(n_335),
.B(n_341),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_2034),
.B(n_1867),
.Y(n_2076)
);

XOR2x2_ASAP7_75t_L g2077 ( 
.A(n_2046),
.B(n_344),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2050),
.Y(n_2078)
);

AOI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_2033),
.A2(n_1837),
.B1(n_1881),
.B2(n_1751),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2033),
.Y(n_2080)
);

XOR2xp5_ASAP7_75t_L g2081 ( 
.A(n_2053),
.B(n_346),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2035),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_2029),
.B(n_1751),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2029),
.B(n_347),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2028),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2028),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2029),
.A2(n_1837),
.B1(n_1728),
.B2(n_1794),
.Y(n_2087)
);

OAI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2029),
.A2(n_1876),
.B1(n_1878),
.B2(n_1924),
.Y(n_2088)
);

HB1xp67_ASAP7_75t_L g2089 ( 
.A(n_2058),
.Y(n_2089)
);

AO22x2_ASAP7_75t_L g2090 ( 
.A1(n_2055),
.A2(n_2086),
.B1(n_2085),
.B2(n_2071),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2064),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2060),
.A2(n_2057),
.B1(n_2061),
.B2(n_2062),
.Y(n_2092)
);

AOI21xp33_ASAP7_75t_L g2093 ( 
.A1(n_2074),
.A2(n_350),
.B(n_351),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2075),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2073),
.A2(n_1794),
.B1(n_1845),
.B2(n_1847),
.Y(n_2095)
);

OAI22x1_ASAP7_75t_L g2096 ( 
.A1(n_2081),
.A2(n_1876),
.B1(n_1923),
.B2(n_356),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_2067),
.Y(n_2097)
);

XNOR2xp5_ASAP7_75t_L g2098 ( 
.A(n_2078),
.B(n_354),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2084),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2070),
.Y(n_2100)
);

XNOR2xp5_ASAP7_75t_L g2101 ( 
.A(n_2077),
.B(n_355),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2083),
.A2(n_1794),
.B1(n_1891),
.B2(n_1894),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2080),
.B(n_1852),
.Y(n_2103)
);

NAND2x1_ASAP7_75t_SL g2104 ( 
.A(n_2082),
.B(n_2079),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2072),
.Y(n_2105)
);

AOI31xp33_ASAP7_75t_L g2106 ( 
.A1(n_2076),
.A2(n_357),
.A3(n_358),
.B(n_359),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_2072),
.Y(n_2107)
);

NAND3xp33_ASAP7_75t_L g2108 ( 
.A(n_2087),
.B(n_2088),
.C(n_2066),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_2063),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2097),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2089),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2107),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2090),
.Y(n_2113)
);

CKINVDCx20_ASAP7_75t_R g2114 ( 
.A(n_2092),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2100),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2090),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2094),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2105),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2098),
.Y(n_2119)
);

CKINVDCx20_ASAP7_75t_R g2120 ( 
.A(n_2101),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2096),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2099),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2109),
.Y(n_2123)
);

XNOR2xp5_ASAP7_75t_L g2124 ( 
.A(n_2091),
.B(n_2068),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2113),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2116),
.A2(n_2093),
.B(n_2106),
.Y(n_2126)
);

AOI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_2111),
.A2(n_2103),
.B1(n_2108),
.B2(n_2065),
.Y(n_2127)
);

CKINVDCx20_ASAP7_75t_R g2128 ( 
.A(n_2114),
.Y(n_2128)
);

OAI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2110),
.A2(n_2102),
.B1(n_2104),
.B2(n_2059),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2123),
.Y(n_2130)
);

BUFx4f_ASAP7_75t_SL g2131 ( 
.A(n_2120),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_2112),
.A2(n_2069),
.B(n_2095),
.Y(n_2132)
);

AOI22x1_ASAP7_75t_L g2133 ( 
.A1(n_2124),
.A2(n_2056),
.B1(n_361),
.B2(n_365),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_2131),
.A2(n_2115),
.B1(n_2117),
.B2(n_2118),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2128),
.A2(n_2122),
.B1(n_2121),
.B2(n_2119),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2125),
.B(n_360),
.Y(n_2136)
);

XNOR2xp5_ASAP7_75t_L g2137 ( 
.A(n_2130),
.B(n_366),
.Y(n_2137)
);

OAI21x1_ASAP7_75t_L g2138 ( 
.A1(n_2126),
.A2(n_1849),
.B(n_1814),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2133),
.A2(n_1794),
.B1(n_1848),
.B2(n_1824),
.Y(n_2139)
);

BUFx2_ASAP7_75t_L g2140 ( 
.A(n_2127),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2134),
.B(n_2129),
.Y(n_2141)
);

OAI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_2140),
.A2(n_2132),
.B1(n_1852),
.B2(n_370),
.Y(n_2142)
);

OAI221xp5_ASAP7_75t_L g2143 ( 
.A1(n_2135),
.A2(n_367),
.B1(n_368),
.B2(n_374),
.C(n_375),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2136),
.B(n_377),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2141),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_2144),
.A2(n_2137),
.B1(n_2139),
.B2(n_2138),
.Y(n_2146)
);

AOI22xp33_ASAP7_75t_SL g2147 ( 
.A1(n_2143),
.A2(n_378),
.B1(n_379),
.B2(n_383),
.Y(n_2147)
);

AOI222xp33_ASAP7_75t_L g2148 ( 
.A1(n_2142),
.A2(n_386),
.B1(n_387),
.B2(n_388),
.C1(n_389),
.C2(n_390),
.Y(n_2148)
);

NOR4xp25_ASAP7_75t_L g2149 ( 
.A(n_2145),
.B(n_391),
.C(n_393),
.D(n_396),
.Y(n_2149)
);

AOI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_2146),
.A2(n_397),
.B1(n_398),
.B2(n_400),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2150),
.A2(n_2148),
.B1(n_2147),
.B2(n_408),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_SL g2152 ( 
.A1(n_2149),
.A2(n_405),
.B(n_407),
.Y(n_2152)
);

AOI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_2152),
.A2(n_2151),
.B(n_413),
.Y(n_2153)
);

AOI211xp5_ASAP7_75t_L g2154 ( 
.A1(n_2153),
.A2(n_412),
.B(n_416),
.C(n_418),
.Y(n_2154)
);


endmodule