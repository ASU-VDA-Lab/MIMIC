module fake_jpeg_32104_n_527 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_57),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_58),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_64),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_70),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_67),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_68),
.Y(n_127)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_1),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_71),
.B(n_84),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_16),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_99),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_33),
.B(n_2),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_85),
.B(n_97),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_33),
.B(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_101),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_41),
.B(n_3),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_48),
.B(n_3),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_4),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_105),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

BUFx12f_ASAP7_75t_SL g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_105),
.B(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_110),
.B(n_117),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_29),
.B1(n_50),
.B2(n_49),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_122),
.A2(n_88),
.B1(n_86),
.B2(n_74),
.Y(n_182)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_79),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_144),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_19),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_148),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_17),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_19),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_156),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_82),
.Y(n_156)
);

INVx2_ASAP7_75t_R g163 ( 
.A(n_85),
.Y(n_163)
);

CKINVDCx9p33_ASAP7_75t_R g194 ( 
.A(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_67),
.B(n_28),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_167),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_72),
.B(n_53),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_132),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_113),
.A2(n_106),
.B1(n_96),
.B2(n_54),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_174),
.A2(n_183),
.B1(n_206),
.B2(n_122),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_176),
.Y(n_236)
);

AOI22x1_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_68),
.B1(n_57),
.B2(n_56),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_177),
.B(n_191),
.Y(n_248)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_196),
.Y(n_244)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_127),
.A2(n_75),
.B1(n_61),
.B2(n_69),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_181),
.A2(n_208),
.B1(n_214),
.B2(n_216),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_182),
.A2(n_193),
.B1(n_209),
.B2(n_34),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_120),
.A2(n_62),
.B1(n_50),
.B2(n_49),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_115),
.B(n_28),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_221),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_192),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_123),
.A2(n_92),
.B1(n_37),
.B2(n_50),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_160),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_195),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_125),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_36),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_212),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_199),
.Y(n_245)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_132),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_138),
.A2(n_49),
.B1(n_37),
.B2(n_100),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_127),
.A2(n_100),
.B1(n_30),
.B2(n_60),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_138),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_209)
);

BUFx24_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_121),
.B(n_44),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_140),
.Y(n_213)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_146),
.B(n_45),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_114),
.Y(n_228)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_137),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_220),
.B1(n_126),
.B2(n_166),
.Y(n_249)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_218),
.B(n_118),
.Y(n_262)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_124),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_228),
.B(n_17),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_144),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_242),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_152),
.B1(n_141),
.B2(n_168),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_230),
.A2(n_239),
.B1(n_240),
.B2(n_243),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_194),
.A2(n_152),
.B1(n_149),
.B2(n_168),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_177),
.A2(n_141),
.B1(n_161),
.B2(n_149),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_241),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_172),
.B(n_212),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_201),
.A2(n_194),
.B(n_212),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_208),
.B(n_195),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_174),
.A2(n_171),
.B1(n_150),
.B2(n_142),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_260),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_173),
.A2(n_161),
.B1(n_169),
.B2(n_133),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_173),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_202),
.A2(n_164),
.B(n_158),
.C(n_43),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_210),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_268),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_204),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_269),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_219),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_181),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_284),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_271),
.B(n_280),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_222),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_277),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_232),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_275),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_223),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_200),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_190),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_184),
.Y(n_279)
);

INVx6_ASAP7_75t_SL g280 ( 
.A(n_232),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_226),
.B(n_178),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_281),
.B(n_282),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_176),
.Y(n_282)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_228),
.A2(n_36),
.B(n_43),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_287),
.B(n_31),
.Y(n_308)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_225),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_217),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_292),
.B(n_293),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_214),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_260),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_319),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_249),
.B(n_258),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_300),
.A2(n_267),
.B(n_263),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_240),
.B1(n_230),
.B2(n_243),
.Y(n_301)
);

OA22x2_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_276),
.B1(n_265),
.B2(n_266),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_308),
.B(n_310),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_241),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_321),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_273),
.B(n_245),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_277),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_268),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_294),
.A2(n_253),
.A3(n_254),
.B1(n_235),
.B2(n_238),
.Y(n_315)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_317),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_254),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_271),
.A2(n_220),
.B1(n_216),
.B2(n_186),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_320),
.A2(n_324),
.B1(n_285),
.B2(n_312),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_272),
.B(n_235),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_272),
.A2(n_175),
.B1(n_224),
.B2(n_231),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_313),
.B(n_279),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_325),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_281),
.C(n_269),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_337),
.C(n_338),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_264),
.Y(n_328)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_306),
.A2(n_270),
.B(n_269),
.Y(n_331)
);

AO21x1_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_342),
.B(n_284),
.Y(n_374)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_270),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_280),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_335),
.A2(n_343),
.B1(n_326),
.B2(n_301),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_336),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_303),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_265),
.C(n_266),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_296),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_340),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_296),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_308),
.B(n_287),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_341),
.B(n_344),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_274),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_299),
.B(n_275),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_347),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_305),
.B(n_275),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_274),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_311),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_321),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_350),
.B(n_351),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_324),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_352),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_307),
.A2(n_292),
.B(n_293),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_353),
.A2(n_323),
.B(n_309),
.Y(n_359)
);

AO22x1_ASAP7_75t_L g355 ( 
.A1(n_333),
.A2(n_318),
.B1(n_300),
.B2(n_315),
.Y(n_355)
);

AO22x1_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_335),
.B1(n_342),
.B2(n_354),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_297),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_329),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_361),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_359),
.B(n_360),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_333),
.A2(n_312),
.B(n_320),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_326),
.A2(n_351),
.B1(n_353),
.B2(n_346),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_311),
.C(n_322),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_357),
.C(n_362),
.Y(n_392)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_372),
.A2(n_335),
.B1(n_331),
.B2(n_354),
.Y(n_388)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_334),
.Y(n_373)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

XOR2x1_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_343),
.Y(n_405)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_376),
.Y(n_401)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_377),
.Y(n_403)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_379),
.B(n_383),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_380),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_347),
.A2(n_336),
.B1(n_350),
.B2(n_340),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_385),
.Y(n_393)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_330),
.B(n_317),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_376),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_339),
.A2(n_276),
.B1(n_304),
.B2(n_298),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_399),
.B1(n_410),
.B2(n_411),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_390),
.B(n_394),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_364),
.B(n_341),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_391),
.B(n_412),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_392),
.B(n_395),
.C(n_397),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_338),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_329),
.C(n_335),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_396),
.A2(n_236),
.B(n_348),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_335),
.C(n_330),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_261),
.Y(n_398)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_355),
.B1(n_371),
.B2(n_358),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_402),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_298),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_380),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_405),
.A2(n_380),
.B1(n_374),
.B2(n_382),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_261),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_359),
.B(n_286),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_385),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_355),
.A2(n_304),
.B1(n_316),
.B2(n_283),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_366),
.A2(n_316),
.B1(n_283),
.B2(n_289),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_289),
.C(n_234),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_413),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_386),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_415),
.B(n_436),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_431),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_417),
.B(n_428),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_387),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_429),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_404),
.A2(n_366),
.B1(n_383),
.B2(n_379),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_419),
.A2(n_410),
.B1(n_397),
.B2(n_412),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_360),
.B(n_370),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_421),
.A2(n_432),
.B(n_438),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_393),
.Y(n_427)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_427),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_375),
.B1(n_377),
.B2(n_373),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_378),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_369),
.B(n_368),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_396),
.A2(n_368),
.B(n_367),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_434),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_408),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_411),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_393),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_437),
.B(n_231),
.Y(n_458)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_401),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_414),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_405),
.B1(n_387),
.B2(n_388),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_447),
.B1(n_423),
.B2(n_259),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_419),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_420),
.A2(n_400),
.B1(n_407),
.B2(n_403),
.Y(n_443)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_456),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_413),
.B1(n_394),
.B2(n_390),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_433),
.B(n_395),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_449),
.B(n_424),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_430),
.A2(n_352),
.B(n_285),
.Y(n_450)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_450),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_250),
.C(n_234),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_454),
.C(n_426),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_250),
.C(n_237),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_252),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_218),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_460),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_453),
.A2(n_416),
.B1(n_434),
.B2(n_435),
.Y(n_460)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_461),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_469),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_455),
.A2(n_421),
.B(n_432),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_463),
.B(n_467),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_446),
.A2(n_424),
.B(n_417),
.Y(n_466)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_454),
.B(n_423),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_237),
.C(n_236),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_474),
.C(n_456),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_439),
.A2(n_259),
.B1(n_286),
.B2(n_238),
.Y(n_472)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_189),
.C(n_166),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_476),
.B(n_452),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_477),
.B(n_479),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_481),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_444),
.C(n_448),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_465),
.A2(n_468),
.B1(n_460),
.B2(n_471),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_457),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_487),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_462),
.A2(n_441),
.B1(n_445),
.B2(n_444),
.Y(n_486)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_486),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_463),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_448),
.C(n_441),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_488),
.B(n_474),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_464),
.A2(n_207),
.B1(n_192),
.B2(n_203),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_489),
.B(n_162),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_198),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_491),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

OAI321xp33_ASAP7_75t_L g496 ( 
.A1(n_483),
.A2(n_473),
.A3(n_198),
.B1(n_211),
.B2(n_162),
.C(n_145),
.Y(n_496)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

NOR3xp33_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_473),
.C(n_60),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_499),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_480),
.B(n_31),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_503),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_484),
.B(n_145),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_492),
.B(n_44),
.Y(n_504)
);

AOI322xp5_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_505),
.A3(n_498),
.B1(n_129),
.B2(n_111),
.C1(n_157),
.C2(n_497),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g505 ( 
.A1(n_492),
.A2(n_211),
.B(n_109),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_500),
.C(n_479),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_510),
.C(n_513),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_502),
.A2(n_490),
.B1(n_486),
.B2(n_491),
.Y(n_510)
);

OAI31xp33_ASAP7_75t_L g515 ( 
.A1(n_511),
.A2(n_58),
.A3(n_159),
.B(n_129),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_494),
.A2(n_488),
.B1(n_477),
.B2(n_34),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_512),
.A2(n_159),
.B(n_58),
.Y(n_514)
);

AOI322xp5_ASAP7_75t_L g521 ( 
.A1(n_514),
.A2(n_518),
.A3(n_6),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_515),
.A2(n_508),
.B1(n_39),
.B2(n_10),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_512),
.A2(n_4),
.B(n_5),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_516),
.B(n_506),
.Y(n_519)
);

AOI21xp33_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_6),
.B(n_7),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_519),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_520),
.A2(n_521),
.B(n_517),
.Y(n_523)
);

AOI322xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_522),
.A3(n_509),
.B1(n_12),
.B2(n_15),
.C1(n_9),
.C2(n_6),
.Y(n_524)
);

INVx11_ASAP7_75t_L g525 ( 
.A(n_524),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_525),
.A2(n_9),
.B1(n_12),
.B2(n_15),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_525),
.B1(n_12),
.B2(n_15),
.Y(n_527)
);


endmodule