module fake_netlist_5_2071_n_30 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_30);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_30;

wire n_29;
wire n_16;
wire n_12;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_10;
wire n_24;
wire n_28;
wire n_21;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_26;
wire n_20;
wire n_14;
wire n_23;
wire n_13;

INVx6_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

NAND3xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_4),
.C(n_8),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_3),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_9),
.B(n_2),
.Y(n_16)
);

AND2x4_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

AO31x2_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_0),
.A3(n_1),
.B(n_3),
.Y(n_18)
);

OAI22x1_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_12),
.B(n_14),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_11),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_21),
.B(n_17),
.Y(n_25)
);

AOI221xp5_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_10),
.B1(n_18),
.B2(n_19),
.C(n_23),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

AOI211x1_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_26),
.B(n_18),
.C(n_10),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_27),
.B(n_25),
.Y(n_30)
);


endmodule