module fake_aes_8241_n_653 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_653);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_653;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_504;
wire n_170;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_67), .Y(n_77) );
INVxp33_ASAP7_75t_SL g78 ( .A(n_45), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_69), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_17), .Y(n_80) );
INVx1_ASAP7_75t_SL g81 ( .A(n_6), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_8), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_33), .Y(n_83) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_64), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_47), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_13), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_72), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_22), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_71), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_65), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_14), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_55), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_73), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_1), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_63), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_27), .Y(n_99) );
BUFx2_ASAP7_75t_L g100 ( .A(n_21), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_14), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_66), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_36), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_35), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_1), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_9), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_32), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_62), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_50), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_28), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_76), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_11), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_52), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_25), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_57), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_54), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_48), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_51), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_8), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_44), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_23), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_100), .B(n_0), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_100), .B(n_0), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_101), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_89), .B(n_80), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_101), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_77), .A2(n_34), .B(n_74), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_124), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
NOR2xp33_ASAP7_75t_R g137 ( .A(n_124), .B(n_31), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_101), .Y(n_138) );
INVxp67_ASAP7_75t_SL g139 ( .A(n_80), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_108), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_82), .B(n_2), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_112), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_78), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_77), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_122), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_79), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_86), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_93), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_83), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_110), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_79), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_121), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_85), .Y(n_157) );
BUFx8_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_94), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_81), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_87), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_81), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_107), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_107), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_121), .B(n_3), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_87), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_163), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_127), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_127), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_133), .A2(n_96), .B1(n_97), .B2(n_103), .Y(n_171) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_165), .B(n_123), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_127), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_158), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_158), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_137), .Y(n_177) );
AND2x6_ASAP7_75t_L g178 ( .A(n_165), .B(n_123), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_165), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_165), .B(n_97), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_139), .B(n_96), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_125), .B(n_120), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_127), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_127), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_129), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_130), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_139), .B(n_103), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_132), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_142), .B(n_106), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_130), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_133), .B(n_106), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_140), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_131), .B(n_104), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_158), .Y(n_197) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_125), .B(n_120), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_125), .B(n_105), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_157), .B(n_104), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_128), .B(n_115), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_132), .Y(n_206) );
NAND3x1_ASAP7_75t_L g207 ( .A(n_128), .B(n_115), .C(n_92), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
NAND3xp33_ASAP7_75t_L g209 ( .A(n_142), .B(n_105), .C(n_90), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_145), .B(n_113), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_156), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_131), .B(n_113), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_132), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_159), .B(n_92), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_156), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_126), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_134), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_132), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g220 ( .A1(n_160), .A2(n_95), .B1(n_109), .B2(n_117), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_151), .A2(n_111), .B1(n_98), .B2(n_117), .Y(n_221) );
OR2x2_ASAP7_75t_SL g222 ( .A(n_145), .B(n_95), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_126), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_126), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_146), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_153), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_134), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_126), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_167), .B(n_128), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_213), .A2(n_152), .B(n_146), .C(n_148), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_167), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_210), .B(n_152), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_187), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_200), .A2(n_144), .B1(n_143), .B2(n_135), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_190), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_196), .B(n_154), .Y(n_236) );
OR2x2_ASAP7_75t_SL g237 ( .A(n_177), .B(n_147), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_210), .B(n_166), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_200), .A2(n_141), .B1(n_164), .B2(n_162), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_195), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_191), .B(n_141), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_226), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_210), .B(n_166), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_190), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_215), .B(n_161), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_194), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_187), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_192), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_200), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_200), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_192), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_199), .Y(n_254) );
OR2x6_ASAP7_75t_L g255 ( .A(n_183), .B(n_198), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_175), .B(n_161), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_191), .B(n_141), .Y(n_257) );
NAND3xp33_ASAP7_75t_L g258 ( .A(n_203), .B(n_155), .C(n_148), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_199), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_176), .Y(n_260) );
BUFx4f_ASAP7_75t_L g261 ( .A(n_200), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_179), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_200), .A2(n_155), .B1(n_114), .B2(n_118), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_200), .A2(n_111), .B1(n_109), .B2(n_98), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_208), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_226), .B(n_134), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_207), .A2(n_116), .B1(n_99), .B2(n_102), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_208), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_179), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_177), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_212), .Y(n_271) );
INVx4_ASAP7_75t_L g272 ( .A(n_176), .Y(n_272) );
NAND2xp33_ASAP7_75t_L g273 ( .A(n_178), .B(n_84), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_191), .B(n_90), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_204), .B(n_88), .Y(n_275) );
NOR3xp33_ASAP7_75t_SL g276 ( .A(n_220), .B(n_3), .C(n_4), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_221), .Y(n_277) );
NOR3xp33_ASAP7_75t_SL g278 ( .A(n_209), .B(n_4), .C(n_5), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_201), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_201), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_178), .Y(n_281) );
NAND2xp33_ASAP7_75t_SL g282 ( .A(n_179), .B(n_119), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_183), .Y(n_283) );
NOR3xp33_ASAP7_75t_SL g284 ( .A(n_206), .B(n_5), .C(n_6), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_183), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_212), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_205), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_198), .Y(n_288) );
INVx3_ASAP7_75t_SL g289 ( .A(n_204), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_198), .B(n_119), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_182), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_175), .A2(n_134), .B(n_119), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_204), .B(n_181), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_206), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_255), .A2(n_172), .B1(n_222), .B2(n_180), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_240), .B(n_222), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_255), .B(n_181), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_235), .Y(n_298) );
HAxp5_ASAP7_75t_L g299 ( .A(n_277), .B(n_207), .CON(n_299), .SN(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_256), .A2(n_172), .B(n_182), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_293), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_262), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_257), .B(n_204), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_255), .Y(n_304) );
OR2x6_ASAP7_75t_L g305 ( .A(n_283), .B(n_172), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_241), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_233), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_248), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_289), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_256), .A2(n_197), .B(n_180), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_257), .B(n_181), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_231), .Y(n_313) );
INVx5_ASAP7_75t_L g314 ( .A(n_291), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_257), .B(n_181), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_235), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_288), .A2(n_180), .B1(n_188), .B2(n_197), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_291), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_291), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_262), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_250), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
NOR2xp33_ASAP7_75t_SL g325 ( .A(n_250), .B(n_178), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_230), .A2(n_193), .B(n_188), .C(n_225), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_292), .A2(n_180), .B(n_227), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_242), .B(n_229), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_232), .B(n_238), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_232), .A2(n_178), .B1(n_188), .B2(n_193), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_249), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_252), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_251), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_261), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_262), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_243), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_238), .A2(n_178), .B1(n_188), .B2(n_225), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_244), .B(n_178), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_282), .A2(n_227), .B(n_218), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_282), .A2(n_227), .B(n_218), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_261), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_281), .B(n_205), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_260), .Y(n_343) );
OR2x6_ASAP7_75t_L g344 ( .A(n_260), .B(n_205), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_281), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_328), .A2(n_277), .B1(n_246), .B2(n_244), .C(n_171), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_297), .B(n_246), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_297), .A2(n_239), .B1(n_178), .B2(n_236), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_313), .Y(n_349) );
NAND3xp33_ASAP7_75t_L g350 ( .A(n_327), .B(n_276), .C(n_284), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_305), .A2(n_290), .B1(n_274), .B2(n_264), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_298), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_308), .B(n_243), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_339), .A2(n_266), .B(n_218), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_297), .B(n_281), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_326), .A2(n_258), .B(n_275), .C(n_279), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_329), .B(n_263), .Y(n_360) );
INVx4_ASAP7_75t_SL g361 ( .A(n_305), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_312), .B(n_254), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_309), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_305), .A2(n_259), .B1(n_280), .B2(n_275), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_317), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_260), .B(n_272), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_328), .A2(n_267), .B1(n_269), .B2(n_270), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_332), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_314), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_316), .Y(n_371) );
NAND2xp33_ASAP7_75t_L g372 ( .A(n_324), .B(n_287), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_317), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_301), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_302), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_334), .B(n_272), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_303), .A2(n_270), .B1(n_234), .B2(n_214), .C(n_219), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_374), .B(n_306), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_361), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_348), .A2(n_305), .B1(n_295), .B2(n_330), .Y(n_380) );
INVx4_ASAP7_75t_SL g381 ( .A(n_370), .Y(n_381) );
OAI22xp33_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_336), .B1(n_296), .B2(n_325), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_346), .A2(n_312), .B1(n_296), .B2(n_315), .C(n_304), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_365), .A2(n_336), .B1(n_308), .B2(n_299), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_347), .A2(n_318), .B1(n_338), .B2(n_337), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_373), .A2(n_299), .B1(n_333), .B2(n_310), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_347), .B(n_189), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_350), .A2(n_344), .B(n_310), .Y(n_388) );
AOI222xp33_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_237), .B1(n_273), .B2(n_214), .C1(n_219), .C2(n_189), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_361), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_368), .A2(n_278), .B1(n_311), .B2(n_300), .C(n_189), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_371), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_377), .A2(n_302), .B1(n_322), .B2(n_335), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_361), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_374), .B(n_322), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_362), .B(n_173), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_359), .A2(n_335), .B1(n_273), .B2(n_343), .C(n_266), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_364), .A2(n_335), .B1(n_343), .B2(n_294), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_362), .A2(n_272), .B1(n_344), .B2(n_341), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_354), .A2(n_186), .B1(n_173), .B2(n_168), .C(n_269), .Y(n_400) );
AOI222xp33_ASAP7_75t_L g401 ( .A1(n_354), .A2(n_186), .B1(n_341), .B2(n_334), .C1(n_168), .C2(n_323), .Y(n_401) );
AOI211xp5_ASAP7_75t_L g402 ( .A1(n_353), .A2(n_84), .B(n_342), .C(n_323), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_361), .Y(n_403) );
OAI211xp5_ASAP7_75t_SL g404 ( .A1(n_363), .A2(n_269), .B(n_286), .C(n_265), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_379), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_390), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_392), .B(n_371), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_392), .Y(n_408) );
AND2x4_ASAP7_75t_SL g409 ( .A(n_394), .B(n_352), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_395), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g411 ( .A1(n_391), .A2(n_351), .B(n_357), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_396), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_396), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_378), .B(n_363), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_378), .B(n_367), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_387), .B(n_352), .Y(n_417) );
NOR4xp25_ASAP7_75t_SL g418 ( .A(n_390), .B(n_367), .C(n_369), .D(n_361), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_403), .Y(n_420) );
NAND4xp25_ASAP7_75t_SL g421 ( .A(n_384), .B(n_369), .C(n_355), .D(n_356), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_403), .B(n_352), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_381), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_380), .A2(n_355), .B1(n_356), .B2(n_375), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_397), .A2(n_357), .B(n_366), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_383), .A2(n_375), .B1(n_370), .B2(n_355), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_387), .B(n_356), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_389), .A2(n_370), .B1(n_344), .B2(n_372), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_381), .B(n_386), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_404), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_402), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g434 ( .A(n_385), .B(n_202), .C(n_211), .D(n_216), .Y(n_434) );
NOR4xp25_ASAP7_75t_SL g435 ( .A(n_402), .B(n_342), .C(n_134), .D(n_10), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_398), .A2(n_321), .B(n_314), .C(n_319), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_401), .B(n_245), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g439 ( .A1(n_393), .A2(n_319), .B(n_314), .C(n_271), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_414), .B(n_382), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_407), .B(n_7), .Y(n_442) );
AOI221x1_ASAP7_75t_L g443 ( .A1(n_433), .A2(n_126), .B1(n_127), .B2(n_136), .C(n_149), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_438), .A2(n_399), .B1(n_400), .B2(n_376), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_430), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_432), .B(n_126), .C(n_127), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_407), .B(n_7), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_414), .B(n_9), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_415), .A2(n_217), .B(n_223), .C(n_224), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_415), .B(n_10), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_408), .B(n_11), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_421), .A2(n_321), .B1(n_314), .B2(n_319), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_410), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_417), .B(n_13), .Y(n_455) );
INVx4_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_406), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_417), .B(n_15), .Y(n_458) );
OAI31xp33_ASAP7_75t_L g459 ( .A1(n_433), .A2(n_358), .A3(n_376), .B(n_211), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_439), .A2(n_320), .B(n_314), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_405), .B(n_15), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_427), .B(n_16), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_409), .Y(n_465) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_434), .A2(n_358), .B1(n_319), .B2(n_320), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_416), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_432), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_430), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_432), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_427), .B(n_16), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_420), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_420), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_412), .B(n_18), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_412), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_405), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_425), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_425), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_422), .Y(n_483) );
AOI221xp5_ASAP7_75t_SL g484 ( .A1(n_426), .A2(n_136), .B1(n_149), .B2(n_265), .C(n_268), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_431), .B(n_136), .C(n_149), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_440), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_442), .B(n_429), .Y(n_487) );
NAND2xp33_ASAP7_75t_SL g488 ( .A(n_456), .B(n_419), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_477), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_474), .B(n_411), .Y(n_490) );
INVx1_ASAP7_75t_SL g491 ( .A(n_457), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_477), .Y(n_492) );
AOI31xp33_ASAP7_75t_L g493 ( .A1(n_462), .A2(n_423), .A3(n_428), .B(n_437), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_442), .B(n_424), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_447), .B(n_424), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_478), .Y(n_496) );
NAND2x2_ASAP7_75t_L g497 ( .A(n_450), .B(n_418), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_474), .B(n_411), .Y(n_498) );
NAND2xp33_ASAP7_75t_SL g499 ( .A(n_456), .B(n_418), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_447), .B(n_423), .Y(n_500) );
INVx1_ASAP7_75t_SL g501 ( .A(n_465), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_478), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_474), .B(n_425), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_465), .Y(n_504) );
OR2x6_ASAP7_75t_L g505 ( .A(n_456), .B(n_439), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_480), .B(n_431), .Y(n_506) );
NAND2xp33_ASAP7_75t_SL g507 ( .A(n_456), .B(n_435), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_480), .B(n_425), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_454), .Y(n_510) );
OAI33xp33_ASAP7_75t_L g511 ( .A1(n_451), .A2(n_19), .A3(n_20), .B1(n_228), .B2(n_223), .B3(n_217), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_483), .B(n_436), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_471), .B(n_149), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_471), .B(n_149), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_467), .Y(n_515) );
NAND2xp33_ASAP7_75t_R g516 ( .A(n_462), .B(n_451), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_460), .B(n_149), .Y(n_517) );
NAND2xp33_ASAP7_75t_R g518 ( .A(n_445), .B(n_24), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_460), .B(n_136), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_455), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_450), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_479), .B(n_136), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_463), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_463), .B(n_136), .Y(n_525) );
NAND2xp33_ASAP7_75t_L g526 ( .A(n_453), .B(n_345), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_473), .Y(n_527) );
NOR3xp33_ASAP7_75t_SL g528 ( .A(n_448), .B(n_26), .C(n_29), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_467), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_455), .B(n_253), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_468), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_473), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_458), .B(n_253), .Y(n_533) );
AOI22x1_ASAP7_75t_L g534 ( .A1(n_452), .A2(n_341), .B1(n_345), .B2(n_324), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_475), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_458), .B(n_247), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_452), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_493), .A2(n_450), .B1(n_441), .B2(n_444), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_528), .A2(n_459), .B(n_464), .Y(n_539) );
AO22x1_ASAP7_75t_L g540 ( .A1(n_522), .A2(n_521), .B1(n_491), .B2(n_501), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_537), .B(n_464), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_515), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_504), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_529), .Y(n_544) );
AOI311xp33_ASAP7_75t_L g545 ( .A1(n_487), .A2(n_466), .A3(n_461), .B(n_472), .C(n_476), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_488), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_489), .B(n_472), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_516), .A2(n_476), .B1(n_469), .B2(n_445), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_488), .B(n_484), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_486), .Y(n_550) );
NAND4xp25_ASAP7_75t_L g551 ( .A(n_516), .B(n_484), .C(n_468), .D(n_470), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_492), .B(n_468), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_511), .B(n_469), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_520), .B(n_470), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g555 ( .A(n_500), .B(n_470), .C(n_482), .D(n_481), .Y(n_555) );
NOR3xp33_ASAP7_75t_SL g556 ( .A(n_518), .B(n_485), .C(n_446), .Y(n_556) );
OAI222xp33_ASAP7_75t_L g557 ( .A1(n_505), .A2(n_469), .B1(n_445), .B2(n_481), .C1(n_482), .C2(n_446), .Y(n_557) );
AOI21xp33_ASAP7_75t_L g558 ( .A1(n_518), .A2(n_482), .B(n_481), .Y(n_558) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_505), .B(n_485), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_508), .A2(n_445), .B(n_449), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
OAI211xp5_ASAP7_75t_SL g562 ( .A1(n_512), .A2(n_228), .B(n_224), .C(n_245), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_502), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_527), .B(n_443), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_532), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_506), .A2(n_169), .B1(n_170), .B2(n_174), .C(n_184), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_535), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_505), .A2(n_443), .B1(n_345), .B2(n_324), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_509), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_509), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g571 ( .A1(n_494), .A2(n_345), .B(n_247), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_490), .B(n_37), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_505), .A2(n_216), .B1(n_287), .B2(n_40), .Y(n_573) );
OAI221xp5_ASAP7_75t_L g574 ( .A1(n_507), .A2(n_185), .B1(n_184), .B2(n_174), .C(n_170), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_510), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_510), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_507), .B(n_38), .C(n_39), .Y(n_577) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_523), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_530), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_495), .B(n_533), .Y(n_581) );
AOI211x1_ASAP7_75t_L g582 ( .A1(n_536), .A2(n_41), .B(n_42), .C(n_43), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_565), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_549), .A2(n_499), .B(n_526), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_570), .Y(n_585) );
OAI21xp5_ASAP7_75t_SL g586 ( .A1(n_546), .A2(n_490), .B(n_498), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_559), .B(n_499), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_543), .Y(n_588) );
AOI211xp5_ASAP7_75t_L g589 ( .A1(n_540), .A2(n_526), .B(n_498), .C(n_503), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_542), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_581), .B(n_503), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_580), .B(n_531), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_555), .B(n_513), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_579), .Y(n_594) );
INVx3_ASAP7_75t_SL g595 ( .A(n_549), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_581), .B(n_514), .Y(n_596) );
XNOR2x2_ASAP7_75t_SL g597 ( .A(n_548), .B(n_497), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_544), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_547), .B(n_514), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_538), .A2(n_534), .B1(n_513), .B2(n_519), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_554), .Y(n_601) );
AO21x1_ASAP7_75t_L g602 ( .A1(n_553), .A2(n_525), .B(n_519), .Y(n_602) );
NOR2xp67_ASAP7_75t_SL g603 ( .A(n_574), .B(n_525), .Y(n_603) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_545), .B(n_517), .C(n_49), .D(n_53), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_539), .A2(n_517), .B1(n_185), .B2(n_184), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_579), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_550), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_561), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_578), .B(n_46), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_571), .A2(n_56), .B(n_58), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_584), .A2(n_577), .B(n_557), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_595), .A2(n_553), .B1(n_577), .B2(n_541), .Y(n_613) );
BUFx3_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_602), .A2(n_567), .B1(n_551), .B2(n_558), .C(n_582), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_604), .B(n_573), .C(n_562), .Y(n_616) );
OAI32xp33_ASAP7_75t_L g617 ( .A1(n_587), .A2(n_564), .A3(n_568), .B1(n_572), .B2(n_569), .Y(n_617) );
AOI322xp5_ASAP7_75t_L g618 ( .A1(n_587), .A2(n_556), .A3(n_576), .B1(n_575), .B2(n_560), .C1(n_552), .C2(n_566), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_611), .A2(n_556), .B(n_60), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_601), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_600), .A2(n_169), .B1(n_184), .B2(n_174), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_605), .B(n_610), .C(n_586), .Y(n_622) );
OAI22xp5_ASAP7_75t_SL g623 ( .A1(n_600), .A2(n_59), .B1(n_61), .B2(n_68), .Y(n_623) );
OAI31xp33_ASAP7_75t_L g624 ( .A1(n_593), .A2(n_70), .A3(n_75), .B(n_169), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_594), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_602), .B(n_170), .Y(n_626) );
NOR2xp33_ASAP7_75t_R g627 ( .A(n_614), .B(n_596), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g628 ( .A(n_613), .B(n_619), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_620), .Y(n_629) );
OAI322xp33_ASAP7_75t_L g630 ( .A1(n_612), .A2(n_591), .A3(n_583), .B1(n_593), .B2(n_592), .C1(n_590), .C2(n_608), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_615), .B(n_592), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_626), .A2(n_597), .B(n_599), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_625), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_625), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_619), .A2(n_594), .B(n_606), .Y(n_635) );
AND4x1_ASAP7_75t_L g636 ( .A(n_624), .B(n_603), .C(n_598), .D(n_607), .Y(n_636) );
OAI22xp5_ASAP7_75t_SL g637 ( .A1(n_623), .A2(n_606), .B1(n_609), .B2(n_585), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_618), .B(n_185), .C(n_585), .D(n_616), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_617), .A2(n_185), .B(n_621), .C(n_622), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_626), .A2(n_595), .B(n_587), .C(n_604), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_612), .A2(n_595), .B1(n_620), .B2(n_589), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_638), .B(n_639), .C(n_641), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_627), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_628), .A2(n_631), .B1(n_636), .B2(n_632), .C(n_637), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_640), .B(n_633), .Y(n_645) );
AO22x2_ASAP7_75t_L g646 ( .A1(n_645), .A2(n_628), .B1(n_633), .B2(n_635), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_643), .B(n_629), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_644), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_647), .Y(n_649) );
XNOR2x1_ASAP7_75t_L g650 ( .A(n_647), .B(n_642), .Y(n_650) );
NOR2x1p5_ASAP7_75t_L g651 ( .A(n_649), .B(n_648), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_651), .A2(n_646), .B1(n_650), .B2(n_634), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_646), .B(n_630), .Y(n_653) );
endmodule