module fake_aes_3526_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
OAI22x1_ASAP7_75t_R g13 ( .A1(n_2), .A2(n_7), .B1(n_8), .B2(n_1), .Y(n_13) );
CKINVDCx11_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
CKINVDCx11_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_12), .B(n_0), .Y(n_16) );
INVx3_ASAP7_75t_SL g17 ( .A(n_11), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
OA21x2_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_12), .B(n_13), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_17), .B(n_15), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_16), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_18), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_19), .B1(n_18), .B2(n_14), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_21), .Y(n_25) );
INVx2_ASAP7_75t_SL g26 ( .A(n_24), .Y(n_26) );
OAI211xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_0), .B(n_3), .C(n_4), .Y(n_27) );
OAI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_3), .B1(n_5), .B2(n_9), .C(n_10), .Y(n_28) );
BUFx8_ASAP7_75t_SL g29 ( .A(n_27), .Y(n_29) );
O2A1O1Ixp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_25), .B(n_26), .C(n_5), .Y(n_30) );
INVxp67_ASAP7_75t_SL g31 ( .A(n_29), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
OAI22xp33_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_25), .B1(n_30), .B2(n_32), .Y(n_33) );
NOR2xp33_ASAP7_75t_L g34 ( .A(n_33), .B(n_32), .Y(n_34) );
endmodule