module fake_jpeg_9025_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_21),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_28),
.B1(n_32),
.B2(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_26),
.B1(n_19),
.B2(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_17),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_73),
.B(n_83),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_34),
.C(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_68),
.Y(n_96)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_89),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_22),
.B(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_75),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_84),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_28),
.B1(n_32),
.B2(n_17),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_44),
.A2(n_28),
.B1(n_32),
.B2(n_17),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_79),
.B1(n_31),
.B2(n_30),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_25),
.B(n_19),
.C(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_61),
.B1(n_51),
.B2(n_54),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_22),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_18),
.B1(n_26),
.B2(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_100),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_18),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_71),
.C(n_92),
.Y(n_138)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_27),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_64),
.B1(n_82),
.B2(n_67),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_59),
.B1(n_33),
.B2(n_31),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_30),
.B1(n_27),
.B2(n_16),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

OAI22x1_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_31),
.B1(n_23),
.B2(n_16),
.Y(n_134)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_80),
.B1(n_31),
.B2(n_23),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_1),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_23),
.B(n_30),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_83),
.B(n_69),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_126),
.B(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_123),
.B(n_127),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_64),
.B(n_69),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_68),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_134),
.B1(n_141),
.B2(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_132),
.B(n_133),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_144),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_1),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_129),
.B(n_144),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_95),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_23),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_149),
.C(n_110),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_82),
.B(n_67),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_93),
.B1(n_88),
.B2(n_86),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_30),
.B1(n_27),
.B2(n_16),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_16),
.Y(n_147)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_80),
.C(n_27),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_152),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_1),
.B(n_2),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_99),
.B(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_121),
.B1(n_118),
.B2(n_101),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_156),
.B(n_159),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_114),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_160),
.C(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_165),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_167),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_172),
.B(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_95),
.Y(n_168)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_179),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_116),
.B1(n_109),
.B2(n_98),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_96),
.C(n_119),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_123),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_121),
.B1(n_96),
.B2(n_118),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_124),
.A2(n_105),
.B1(n_100),
.B2(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_139),
.C(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_177),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_180),
.B(n_167),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_183),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_125),
.B1(n_124),
.B2(n_150),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_210),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_137),
.B(n_130),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_194),
.A2(n_206),
.B(n_207),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_135),
.B1(n_125),
.B2(n_130),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_197),
.B1(n_154),
.B2(n_156),
.Y(n_215)
);

OAI22x1_ASAP7_75t_SL g196 ( 
.A1(n_161),
.A2(n_137),
.B1(n_136),
.B2(n_142),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_180),
.B1(n_183),
.B2(n_163),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_179),
.B1(n_166),
.B2(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_5),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_158),
.B(n_177),
.C(n_176),
.D(n_171),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_174),
.Y(n_221)
);

AO32x1_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_142),
.A3(n_9),
.B1(n_11),
.B2(n_15),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_160),
.C(n_182),
.Y(n_216)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_197),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_226),
.B1(n_210),
.B2(n_190),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_218),
.C(n_219),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_154),
.C(n_172),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_157),
.C(n_174),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_222),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_8),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_224),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_236),
.B(n_194),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_195),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_4),
.C(n_5),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_233),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_211),
.C(n_199),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_196),
.B(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_209),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_239),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_200),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_198),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_215),
.A2(n_192),
.B1(n_190),
.B2(n_201),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_225),
.B1(n_212),
.B2(n_203),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_251),
.B(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_226),
.Y(n_268)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_218),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_270),
.C(n_271),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_217),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_221),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_266),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_192),
.B(n_219),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_248),
.B1(n_253),
.B2(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_243),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_216),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_239),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_233),
.C(n_222),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_229),
.C(n_203),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_247),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_278),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_251),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_240),
.B1(n_250),
.B2(n_230),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_284),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_256),
.C(n_230),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_266),
.C(n_260),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_205),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_290),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_269),
.C(n_258),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_267),
.B(n_259),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_14),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_259),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_287),
.A2(n_283),
.B1(n_281),
.B2(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_274),
.C(n_263),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_286),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_292),
.A2(n_274),
.B1(n_11),
.B2(n_13),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_303),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_11),
.B(n_13),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_285),
.C(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_307),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_289),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_293),
.B(n_302),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_305),
.B(n_302),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_310),
.B(n_306),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_14),
.C(n_15),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_5),
.C(n_7),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_7),
.C(n_102),
.Y(n_315)
);


endmodule