module fake_jpeg_19575_n_356 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_38),
.B(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_50),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_55),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_44),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_24),
.B(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_44),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_34),
.B1(n_17),
.B2(n_22),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_76),
.B(n_74),
.C(n_85),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_35),
.B1(n_32),
.B2(n_26),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_83),
.B1(n_87),
.B2(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_68),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_44),
.Y(n_104)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_17),
.B1(n_35),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_55),
.B1(n_43),
.B2(n_53),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_31),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_44),
.C(n_48),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_35),
.B1(n_32),
.B2(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_44),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_32),
.B1(n_26),
.B2(n_17),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_89),
.B(n_112),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_94),
.B1(n_113),
.B2(n_117),
.Y(n_133)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_36),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_60),
.C(n_44),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_54),
.B1(n_45),
.B2(n_16),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_95),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_22),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_20),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_20),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_82),
.B(n_19),
.Y(n_146)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_60),
.B(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_45),
.Y(n_134)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx9p33_ASAP7_75t_R g109 ( 
.A(n_59),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_42),
.B1(n_43),
.B2(n_41),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_71),
.B1(n_57),
.B2(n_45),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_41),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_114),
.Y(n_148)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_125),
.Y(n_141)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_18),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_119),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_67),
.B(n_18),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_29),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_67),
.Y(n_125)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_127),
.A2(n_90),
.B1(n_107),
.B2(n_56),
.Y(n_145)
);

AOI22x1_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_65),
.B1(n_58),
.B2(n_57),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_128),
.A2(n_56),
.B1(n_62),
.B2(n_51),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_89),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_116),
.C(n_112),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_75),
.B1(n_117),
.B2(n_127),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_131),
.A2(n_145),
.B1(n_146),
.B2(n_56),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_70),
.B(n_82),
.C(n_51),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_152),
.B1(n_89),
.B2(n_93),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_58),
.B1(n_81),
.B2(n_75),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_48),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_99),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_154),
.B(n_155),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_48),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_95),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_119),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_160),
.B(n_165),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_177),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_189),
.B(n_132),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_123),
.B1(n_93),
.B2(n_125),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_168),
.B1(n_171),
.B2(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_115),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_182),
.C(n_134),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_123),
.B1(n_124),
.B2(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_29),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_183),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_92),
.B1(n_126),
.B2(n_120),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_158),
.A2(n_24),
.B(n_33),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_172),
.A2(n_191),
.B(n_143),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_132),
.B(n_143),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_135),
.B1(n_158),
.B2(n_156),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_126),
.B1(n_114),
.B2(n_108),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_192),
.B1(n_193),
.B2(n_149),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_121),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_97),
.C(n_96),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_97),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_0),
.B(n_1),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_96),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_30),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_128),
.A2(n_90),
.B1(n_62),
.B2(n_31),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_31),
.B1(n_30),
.B2(n_8),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_129),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_195),
.B(n_208),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_141),
.B1(n_133),
.B2(n_130),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_197),
.B(n_206),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_201),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_209),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_151),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_147),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_216),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_220),
.B1(n_191),
.B2(n_180),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_181),
.A2(n_145),
.B1(n_142),
.B2(n_150),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_222),
.B1(n_211),
.B2(n_220),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_140),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_9),
.C(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_140),
.Y(n_218)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_142),
.B1(n_144),
.B2(n_8),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_170),
.Y(n_223)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_144),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_13),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_163),
.B(n_1),
.Y(n_228)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_233),
.B1(n_235),
.B2(n_238),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_240),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_191),
.B1(n_179),
.B2(n_183),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_188),
.B1(n_163),
.B2(n_187),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_213),
.A2(n_161),
.B1(n_175),
.B2(n_164),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_171),
.B1(n_173),
.B2(n_186),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_248),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_173),
.B1(n_185),
.B2(n_189),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_241),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_203),
.A2(n_193),
.B1(n_178),
.B2(n_10),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_204),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_195),
.B(n_210),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_206),
.C(n_212),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_261),
.C(n_275),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_203),
.B1(n_208),
.B2(n_197),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_260),
.A2(n_248),
.B1(n_250),
.B2(n_237),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_209),
.C(n_198),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_278),
.B1(n_263),
.B2(n_277),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_255),
.B(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_201),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_227),
.C(n_226),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_277),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_228),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_296),
.B1(n_273),
.B2(n_272),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_234),
.B1(n_244),
.B2(n_255),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_287),
.B1(n_276),
.B2(n_264),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_289),
.B(n_262),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_265),
.Y(n_285)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_236),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_298),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_255),
.B1(n_239),
.B2(n_237),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_257),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_294),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_238),
.B(n_231),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_245),
.Y(n_294)
);

A2O1A1O1Ixp25_ASAP7_75t_L g297 ( 
.A1(n_263),
.A2(n_252),
.B(n_243),
.C(n_242),
.D(n_10),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_274),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_266),
.A2(n_10),
.B(n_9),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_309),
.B1(n_313),
.B2(n_3),
.Y(n_323)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_305),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_275),
.C(n_259),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_315),
.C(n_299),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_312),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_264),
.B1(n_262),
.B2(n_9),
.Y(n_309)
);

OAI321xp33_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_298),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_2),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_280),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_5),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_293),
.C(n_287),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_317),
.C(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_292),
.C(n_282),
.Y(n_317)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_320),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_289),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_321),
.B(n_306),
.Y(n_331)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_323),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_3),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_4),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_303),
.C(n_308),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_322),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_331),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_319),
.A2(n_301),
.B1(n_302),
.B2(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_325),
.B(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_328),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_341),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_338),
.B1(n_336),
.B2(n_335),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_317),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_342),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_316),
.B(n_324),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_7),
.Y(n_348)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_339),
.A2(n_326),
.B(n_5),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_348),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_349),
.B(n_344),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_342),
.B(n_346),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_350),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_345),
.B(n_7),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_7),
.Y(n_356)
);


endmodule