module real_aes_8162_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g124 ( .A(n_0), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_1), .A2(n_153), .B(n_156), .C(n_159), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_2), .A2(n_179), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g539 ( .A(n_3), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_4), .B(n_202), .Y(n_225) );
AOI21xp33_ASAP7_75t_L g466 ( .A1(n_5), .A2(n_179), .B(n_467), .Y(n_466) );
AND2x6_ASAP7_75t_L g153 ( .A(n_6), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g186 ( .A(n_7), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_8), .B(n_107), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_8), .B(n_41), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_9), .A2(n_233), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_10), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g471 ( .A(n_11), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_12), .B(n_208), .Y(n_510) );
INVx1_ASAP7_75t_L g145 ( .A(n_13), .Y(n_145) );
INVx1_ASAP7_75t_L g522 ( .A(n_14), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_15), .A2(n_187), .B(n_197), .C(n_200), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_16), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_17), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_18), .B(n_478), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_19), .B(n_179), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_20), .B(n_243), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_21), .A2(n_208), .B(n_209), .C(n_211), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_22), .B(n_202), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_23), .B(n_165), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_24), .A2(n_199), .B(n_200), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_25), .B(n_165), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_26), .Y(n_261) );
INVx1_ASAP7_75t_L g251 ( .A(n_27), .Y(n_251) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_29), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_30), .B(n_165), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_31), .A2(n_65), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_31), .Y(n_130) );
INVx1_ASAP7_75t_L g238 ( .A(n_32), .Y(n_238) );
INVx1_ASAP7_75t_L g460 ( .A(n_33), .Y(n_460) );
INVx2_ASAP7_75t_L g151 ( .A(n_34), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_35), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_36), .A2(n_208), .B(n_221), .C(n_223), .Y(n_220) );
INVxp67_ASAP7_75t_L g240 ( .A(n_37), .Y(n_240) );
CKINVDCx14_ASAP7_75t_R g219 ( .A(n_38), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_39), .A2(n_156), .B(n_250), .C(n_254), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_40), .A2(n_153), .B(n_156), .C(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g107 ( .A(n_41), .Y(n_107) );
INVx1_ASAP7_75t_L g459 ( .A(n_42), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_43), .A2(n_167), .B(n_184), .C(n_185), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_44), .B(n_165), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_45), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_46), .Y(n_235) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_47), .A2(n_448), .B1(n_723), .B2(n_726), .C1(n_727), .C2(n_729), .Y(n_447) );
INVx1_ASAP7_75t_L g206 ( .A(n_48), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_49), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_50), .B(n_179), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_51), .A2(n_156), .B1(n_211), .B2(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_52), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_53), .Y(n_536) );
CKINVDCx14_ASAP7_75t_R g181 ( .A(n_54), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_55), .A2(n_184), .B(n_223), .C(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_56), .Y(n_502) );
INVx1_ASAP7_75t_L g468 ( .A(n_57), .Y(n_468) );
INVx1_ASAP7_75t_L g154 ( .A(n_58), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_59), .A2(n_78), .B1(n_724), .B2(n_725), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_59), .Y(n_725) );
INVx1_ASAP7_75t_L g144 ( .A(n_60), .Y(n_144) );
INVx1_ASAP7_75t_SL g222 ( .A(n_61), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_62), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_63), .A2(n_102), .B1(n_113), .B2(n_733), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_64), .B(n_202), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_65), .Y(n_129) );
INVx1_ASAP7_75t_L g264 ( .A(n_66), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_SL g477 ( .A1(n_67), .A2(n_223), .B(n_478), .C(n_479), .Y(n_477) );
INVxp67_ASAP7_75t_L g480 ( .A(n_68), .Y(n_480) );
INVx1_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_70), .A2(n_179), .B(n_180), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_71), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_72), .A2(n_179), .B(n_194), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_73), .Y(n_463) );
INVx1_ASAP7_75t_L g496 ( .A(n_74), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_75), .A2(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g195 ( .A(n_76), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_77), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_78), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_79), .A2(n_153), .B(n_156), .C(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_80), .A2(n_179), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g198 ( .A(n_81), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_82), .B(n_239), .Y(n_490) );
INVx2_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g160 ( .A(n_84), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_85), .B(n_478), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_86), .A2(n_153), .B(n_156), .C(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g121 ( .A(n_87), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g722 ( .A(n_87), .B(n_123), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_88), .A2(n_156), .B(n_263), .C(n_266), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_89), .B(n_141), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_90), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_91), .A2(n_153), .B(n_156), .C(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_92), .Y(n_514) );
INVx1_ASAP7_75t_L g476 ( .A(n_93), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_94), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_95), .B(n_239), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_96), .B(n_172), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_97), .B(n_172), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g210 ( .A(n_99), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_100), .A2(n_179), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g734 ( .A(n_105), .Y(n_734) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
OR2x2_ASAP7_75t_L g719 ( .A(n_109), .B(n_123), .Y(n_719) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_109), .B(n_122), .Y(n_731) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_446), .Y(n_113) );
BUFx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g732 ( .A(n_118), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_126), .B(n_443), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_121), .Y(n_445) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_131), .B2(n_132), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g448 ( .A1(n_131), .A2(n_449), .B1(n_717), .B2(n_720), .Y(n_448) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_132), .A2(n_717), .B1(n_722), .B2(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_398), .Y(n_132) );
NAND5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_310), .C(n_348), .D(n_369), .E(n_386), .Y(n_133) );
NOR3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_282), .C(n_303), .Y(n_134) );
OAI221xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_214), .B1(n_245), .B2(n_269), .C(n_273), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_174), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_138), .B(n_271), .Y(n_290) );
OR2x2_ASAP7_75t_L g317 ( .A(n_138), .B(n_191), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_138), .B(n_191), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_138), .B(n_177), .Y(n_345) );
AND2x2_ASAP7_75t_L g383 ( .A(n_138), .B(n_347), .Y(n_383) );
AND2x2_ASAP7_75t_L g412 ( .A(n_138), .B(n_322), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_138), .B(n_294), .Y(n_429) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g309 ( .A(n_139), .B(n_190), .Y(n_309) );
BUFx3_ASAP7_75t_L g334 ( .A(n_139), .Y(n_334) );
AND2x2_ASAP7_75t_L g363 ( .A(n_139), .B(n_191), .Y(n_363) );
AND3x2_ASAP7_75t_L g376 ( .A(n_139), .B(n_377), .C(n_378), .Y(n_376) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_146), .B(n_169), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_140), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_140), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_140), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_141), .A2(n_178), .B(n_189), .Y(n_177) );
INVx2_ASAP7_75t_L g244 ( .A(n_141), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_141), .A2(n_148), .B(n_248), .C(n_249), .Y(n_247) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_141), .A2(n_517), .B(n_523), .Y(n_516) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g173 ( .A(n_142), .B(n_143), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_155), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_148), .A2(n_261), .B(n_262), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_148), .A2(n_188), .B1(n_457), .B2(n_461), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_148), .A2(n_496), .B(n_497), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_148), .A2(n_536), .B(n_537), .Y(n_535) );
NAND2x1p5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
AND2x4_ASAP7_75t_L g179 ( .A(n_149), .B(n_153), .Y(n_179) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g241 ( .A(n_150), .Y(n_241) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx1_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
INVx3_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
INVx1_ASAP7_75t_L g478 ( .A(n_152), .Y(n_478) );
INVx4_ASAP7_75t_SL g188 ( .A(n_153), .Y(n_188) );
BUFx3_ASAP7_75t_L g254 ( .A(n_153), .Y(n_254) );
INVx5_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx3_ASAP7_75t_L g168 ( .A(n_157), .Y(n_168) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
O2A1O1Ixp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_164), .C(n_166), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_161), .A2(n_166), .B(n_264), .C(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_162), .A2(n_163), .B1(n_459), .B2(n_460), .Y(n_458) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx4_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
INVx2_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
INVx4_ASAP7_75t_L g208 ( .A(n_165), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_166), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_166), .A2(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx3_ASAP7_75t_L g202 ( .A(n_171), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_171), .B(n_256), .Y(n_255) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_171), .A2(n_260), .B(n_267), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g492 ( .A(n_171), .B(n_493), .Y(n_492) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_172), .Y(n_192) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_172), .A2(n_474), .B(n_481), .Y(n_473) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g231 ( .A(n_173), .Y(n_231) );
INVx1_ASAP7_75t_L g299 ( .A(n_174), .Y(n_299) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_190), .Y(n_174) );
AOI32xp33_ASAP7_75t_L g354 ( .A1(n_175), .A2(n_306), .A3(n_355), .B1(n_358), .B2(n_359), .Y(n_354) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g281 ( .A(n_176), .B(n_190), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_176), .B(n_309), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_176), .B(n_331), .Y(n_359) );
OR2x2_ASAP7_75t_L g365 ( .A(n_176), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_176), .B(n_320), .Y(n_390) );
OR2x2_ASAP7_75t_L g408 ( .A(n_176), .B(n_227), .Y(n_408) );
BUFx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g272 ( .A(n_177), .B(n_203), .Y(n_272) );
INVx2_ASAP7_75t_L g294 ( .A(n_177), .Y(n_294) );
OR2x2_ASAP7_75t_L g316 ( .A(n_177), .B(n_203), .Y(n_316) );
AND2x2_ASAP7_75t_L g321 ( .A(n_177), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_177), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g377 ( .A(n_177), .B(n_271), .Y(n_377) );
BUFx2_ASAP7_75t_L g233 ( .A(n_179), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_SL g180 ( .A1(n_181), .A2(n_182), .B(n_183), .C(n_188), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_SL g194 ( .A1(n_182), .A2(n_188), .B(n_195), .C(n_196), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_SL g205 ( .A1(n_182), .A2(n_188), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_182), .A2(n_188), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_SL g234 ( .A1(n_182), .A2(n_188), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_182), .A2(n_188), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_182), .A2(n_188), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_182), .A2(n_188), .B(n_519), .C(n_520), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx5_ASAP7_75t_L g239 ( .A(n_187), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_187), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_187), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g266 ( .A(n_188), .Y(n_266) );
INVx1_ASAP7_75t_SL g428 ( .A(n_190), .Y(n_428) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_203), .Y(n_190) );
INVx1_ASAP7_75t_SL g271 ( .A(n_191), .Y(n_271) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_191), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_191), .B(n_357), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_191), .B(n_294), .C(n_412), .Y(n_423) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_201), .Y(n_191) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_192), .A2(n_204), .B(n_213), .Y(n_203) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_192), .A2(n_217), .B(n_225), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_199), .B(n_210), .Y(n_209) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_199), .A2(n_238), .B1(n_239), .B2(n_240), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_199), .B(n_522), .Y(n_521) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_202), .A2(n_466), .B(n_472), .Y(n_465) );
INVx2_ASAP7_75t_L g322 ( .A(n_203), .Y(n_322) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_203), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_208), .B(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g541 ( .A(n_211), .Y(n_541) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_226), .Y(n_214) );
INVx1_ASAP7_75t_L g358 ( .A(n_215), .Y(n_358) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g276 ( .A(n_216), .B(n_258), .Y(n_276) );
INVx2_ASAP7_75t_L g293 ( .A(n_216), .Y(n_293) );
AND2x2_ASAP7_75t_L g298 ( .A(n_216), .B(n_259), .Y(n_298) );
AND2x2_ASAP7_75t_L g313 ( .A(n_216), .B(n_246), .Y(n_313) );
AND2x2_ASAP7_75t_L g325 ( .A(n_216), .B(n_297), .Y(n_325) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_224), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_226), .B(n_341), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_226), .B(n_298), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_226), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_226), .B(n_292), .Y(n_420) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g257 ( .A(n_227), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_227), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g302 ( .A(n_227), .B(n_246), .Y(n_302) );
AND2x2_ASAP7_75t_L g328 ( .A(n_227), .B(n_258), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_227), .B(n_368), .Y(n_367) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_232), .B(n_242), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_229), .A2(n_287), .B(n_288), .Y(n_286) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_229), .A2(n_495), .B(n_501), .Y(n_494) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AOI21xp5_ASAP7_75t_SL g486 ( .A1(n_230), .A2(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_231), .A2(n_456), .B(n_462), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_231), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_231), .A2(n_535), .B(n_542), .Y(n_534) );
INVx1_ASAP7_75t_L g287 ( .A(n_232), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_237), .B(n_241), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_239), .A2(n_251), .B(n_252), .C(n_253), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_239), .A2(n_539), .B(n_540), .C(n_541), .Y(n_538) );
INVx2_ASAP7_75t_L g253 ( .A(n_241), .Y(n_253) );
INVx1_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_244), .B(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_244), .A2(n_506), .B(n_513), .Y(n_505) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_257), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_246), .B(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g292 ( .A(n_246), .B(n_293), .Y(n_292) );
INVx3_ASAP7_75t_SL g297 ( .A(n_246), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_246), .B(n_284), .Y(n_350) );
OR2x2_ASAP7_75t_L g360 ( .A(n_246), .B(n_286), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_246), .B(n_328), .Y(n_388) );
OR2x2_ASAP7_75t_L g418 ( .A(n_246), .B(n_258), .Y(n_418) );
AND2x2_ASAP7_75t_L g422 ( .A(n_246), .B(n_259), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_246), .B(n_298), .Y(n_435) );
AND2x2_ASAP7_75t_L g442 ( .A(n_246), .B(n_324), .Y(n_442) );
OR2x6_ASAP7_75t_L g246 ( .A(n_247), .B(n_255), .Y(n_246) );
INVx1_ASAP7_75t_SL g385 ( .A(n_257), .Y(n_385) );
AND2x2_ASAP7_75t_L g324 ( .A(n_258), .B(n_286), .Y(n_324) );
AND2x2_ASAP7_75t_L g338 ( .A(n_258), .B(n_293), .Y(n_338) );
AND2x2_ASAP7_75t_L g341 ( .A(n_258), .B(n_297), .Y(n_341) );
INVx1_ASAP7_75t_L g368 ( .A(n_258), .Y(n_368) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_L g280 ( .A(n_259), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_270), .A2(n_316), .B(n_440), .C(n_441), .Y(n_439) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g346 ( .A(n_271), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_272), .B(n_289), .Y(n_304) );
AND2x2_ASAP7_75t_L g330 ( .A(n_272), .B(n_331), .Y(n_330) );
OAI21xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_277), .B(n_281), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_275), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g301 ( .A(n_276), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_276), .B(n_297), .Y(n_342) );
AND2x2_ASAP7_75t_L g433 ( .A(n_276), .B(n_284), .Y(n_433) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g306 ( .A(n_280), .B(n_293), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_280), .B(n_291), .Y(n_307) );
OAI322xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_290), .A3(n_291), .B1(n_294), .B2(n_295), .C1(n_299), .C2(n_300), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_289), .Y(n_283) );
AND2x2_ASAP7_75t_L g394 ( .A(n_284), .B(n_306), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_284), .B(n_358), .Y(n_440) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g337 ( .A(n_286), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g403 ( .A(n_290), .B(n_316), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_291), .B(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_292), .B(n_324), .Y(n_381) );
AND2x2_ASAP7_75t_L g327 ( .A(n_293), .B(n_297), .Y(n_327) );
AND2x2_ASAP7_75t_L g335 ( .A(n_294), .B(n_336), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_294), .A2(n_373), .B(n_433), .C(n_434), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g405 ( .A1(n_295), .A2(n_308), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_297), .B(n_324), .Y(n_364) );
AND2x2_ASAP7_75t_L g370 ( .A(n_297), .B(n_338), .Y(n_370) );
AND2x2_ASAP7_75t_L g404 ( .A(n_297), .B(n_306), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_298), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_SL g414 ( .A(n_298), .Y(n_414) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_302), .A2(n_330), .B1(n_332), .B2(n_337), .Y(n_329) );
OAI22xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_305), .B1(n_307), .B2(n_308), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_304), .A2(n_340), .B1(n_342), .B2(n_343), .Y(n_339) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_309), .A2(n_411), .B1(n_413), .B2(n_415), .C(n_419), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B(n_318), .C(n_339), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OR2x2_ASAP7_75t_L g380 ( .A(n_316), .B(n_333), .Y(n_380) );
INVx1_ASAP7_75t_L g431 ( .A(n_316), .Y(n_431) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_317), .A2(n_319), .B1(n_323), .B2(n_326), .C(n_329), .Y(n_318) );
INVx2_ASAP7_75t_SL g373 ( .A(n_317), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g438 ( .A(n_320), .Y(n_438) );
AND2x2_ASAP7_75t_L g362 ( .A(n_321), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g347 ( .A(n_322), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g409 ( .A(n_325), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_333), .B(n_435), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_337), .A2(n_349), .B(n_351), .C(n_353), .Y(n_348) );
INVx1_ASAP7_75t_L g426 ( .A(n_340), .Y(n_426) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_344), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx2_ASAP7_75t_L g357 ( .A(n_347), .Y(n_357) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI222xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_360), .B1(n_361), .B2(n_364), .C1(n_365), .C2(n_367), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g393 ( .A(n_357), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_360), .B(n_414), .Y(n_413) );
NAND2xp33_ASAP7_75t_SL g391 ( .A(n_361), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g366 ( .A(n_363), .Y(n_366) );
AND2x2_ASAP7_75t_L g430 ( .A(n_363), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g396 ( .A(n_366), .B(n_393), .Y(n_396) );
INVx1_ASAP7_75t_L g425 ( .A(n_367), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B(n_374), .C(n_379), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_373), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
AOI322xp5_ASAP7_75t_L g424 ( .A1(n_376), .A2(n_404), .A3(n_409), .B1(n_425), .B2(n_426), .C1(n_427), .C2(n_430), .Y(n_424) );
AND2x2_ASAP7_75t_L g411 ( .A(n_377), .B(n_412), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_382), .B2(n_384), .Y(n_379) );
INVxp33_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B1(n_391), .B2(n_394), .C(n_395), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
NAND5xp2_ASAP7_75t_L g398 ( .A(n_399), .B(n_410), .C(n_424), .D(n_432), .E(n_436), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_404), .B(n_405), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp33_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_412), .A2(n_437), .B(n_438), .C(n_439), .Y(n_436) );
AOI31xp33_ASAP7_75t_L g419 ( .A1(n_414), .A2(n_420), .A3(n_421), .B(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g437 ( .A(n_435), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_443), .B(n_447), .C(n_732), .Y(n_446) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g728 ( .A(n_449), .Y(n_728) );
AND3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_642), .C(n_691), .Y(n_449) );
NOR3xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_549), .C(n_587), .Y(n_450) );
OAI222xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_482), .B1(n_524), .B2(n_530), .C1(n_544), .C2(n_547), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_464), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_453), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_453), .B(n_592), .Y(n_683) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g560 ( .A(n_454), .B(n_473), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_454), .B(n_465), .Y(n_568) );
AND2x2_ASAP7_75t_L g603 ( .A(n_454), .B(n_580), .Y(n_603) );
OR2x2_ASAP7_75t_L g627 ( .A(n_454), .B(n_465), .Y(n_627) );
OR2x2_ASAP7_75t_L g635 ( .A(n_454), .B(n_534), .Y(n_635) );
AND2x2_ASAP7_75t_L g638 ( .A(n_454), .B(n_473), .Y(n_638) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g532 ( .A(n_455), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g546 ( .A(n_455), .B(n_473), .Y(n_546) );
AND2x2_ASAP7_75t_L g596 ( .A(n_455), .B(n_534), .Y(n_596) );
AND2x2_ASAP7_75t_L g609 ( .A(n_455), .B(n_465), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_455), .B(n_695), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_464), .A2(n_635), .B(n_636), .C(n_639), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_464), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_464), .B(n_579), .Y(n_701) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .Y(n_464) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_465), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g559 ( .A(n_465), .Y(n_559) );
AND2x2_ASAP7_75t_L g586 ( .A(n_465), .B(n_580), .Y(n_586) );
INVx1_ASAP7_75t_SL g594 ( .A(n_465), .Y(n_594) );
AND2x2_ASAP7_75t_L g617 ( .A(n_465), .B(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g695 ( .A(n_465), .Y(n_695) );
BUFx2_ASAP7_75t_L g531 ( .A(n_473), .Y(n_531) );
INVx1_ASAP7_75t_L g593 ( .A(n_473), .Y(n_593) );
INVx3_ASAP7_75t_L g618 ( .A(n_473), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_482), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_503), .Y(n_482) );
INVx1_ASAP7_75t_L g614 ( .A(n_483), .Y(n_614) );
OAI32xp33_ASAP7_75t_L g620 ( .A1(n_483), .A2(n_559), .A3(n_621), .B1(n_622), .B2(n_623), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_483), .A2(n_625), .B1(n_628), .B2(n_633), .Y(n_624) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g562 ( .A(n_484), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g640 ( .A(n_484), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g710 ( .A(n_484), .B(n_656), .Y(n_710) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
AND2x2_ASAP7_75t_L g525 ( .A(n_485), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g555 ( .A(n_485), .Y(n_555) );
INVx1_ASAP7_75t_L g574 ( .A(n_485), .Y(n_574) );
OR2x2_ASAP7_75t_L g582 ( .A(n_485), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g589 ( .A(n_485), .B(n_563), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_485), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g610 ( .A(n_485), .B(n_528), .Y(n_610) );
INVx3_ASAP7_75t_L g632 ( .A(n_485), .Y(n_632) );
AND2x2_ASAP7_75t_L g657 ( .A(n_485), .B(n_529), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_485), .B(n_622), .Y(n_705) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
INVx2_ASAP7_75t_L g529 ( .A(n_494), .Y(n_529) );
AND2x2_ASAP7_75t_L g661 ( .A(n_494), .B(n_504), .Y(n_661) );
INVx2_ASAP7_75t_L g703 ( .A(n_503), .Y(n_703) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
INVx1_ASAP7_75t_L g548 ( .A(n_504), .Y(n_548) );
AND2x2_ASAP7_75t_L g575 ( .A(n_504), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_504), .B(n_529), .Y(n_583) );
AND2x2_ASAP7_75t_L g641 ( .A(n_504), .B(n_564), .Y(n_641) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g527 ( .A(n_505), .Y(n_527) );
AND2x2_ASAP7_75t_L g554 ( .A(n_505), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g563 ( .A(n_505), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_505), .B(n_529), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_512), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_511), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_515), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g576 ( .A(n_515), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_515), .B(n_529), .Y(n_622) );
AND2x2_ASAP7_75t_L g631 ( .A(n_515), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g656 ( .A(n_515), .Y(n_656) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g528 ( .A(n_516), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g564 ( .A(n_516), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_524), .A2(n_534), .B1(n_693), .B2(n_696), .Y(n_692) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
OAI21xp5_ASAP7_75t_SL g715 ( .A1(n_526), .A2(n_637), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_527), .B(n_632), .Y(n_649) );
INVx1_ASAP7_75t_L g674 ( .A(n_527), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_528), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g601 ( .A(n_528), .B(n_554), .Y(n_601) );
INVx2_ASAP7_75t_L g557 ( .A(n_529), .Y(n_557) );
INVx1_ASAP7_75t_L g607 ( .A(n_529), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g698 ( .A1(n_530), .A2(n_682), .B1(n_699), .B2(n_702), .C(n_704), .Y(n_698) );
OR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g569 ( .A(n_531), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_531), .B(n_580), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_532), .B(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g623 ( .A(n_532), .B(n_569), .Y(n_623) );
INVx3_ASAP7_75t_SL g664 ( .A(n_532), .Y(n_664) );
AND2x2_ASAP7_75t_L g608 ( .A(n_533), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g637 ( .A(n_533), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_533), .B(n_546), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_533), .B(n_592), .Y(n_678) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g580 ( .A(n_534), .Y(n_580) );
OAI322xp33_ASAP7_75t_L g675 ( .A1(n_534), .A2(n_606), .A3(n_628), .B1(n_676), .B2(n_678), .C1(n_679), .C2(n_680), .Y(n_675) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_545), .A2(n_548), .B(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_SL g625 ( .A(n_546), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g647 ( .A(n_546), .B(n_559), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_546), .B(n_586), .Y(n_662) );
INVxp67_ASAP7_75t_L g613 ( .A(n_548), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g619 ( .A1(n_548), .A2(n_620), .B(n_624), .C(n_634), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_558), .B1(n_561), .B2(n_565), .C(n_570), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g573 ( .A(n_557), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g690 ( .A(n_557), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_558), .A2(n_707), .B1(n_712), .B2(n_713), .C(n_715), .Y(n_706) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_559), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g606 ( .A(n_559), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_559), .B(n_637), .Y(n_644) );
AND2x2_ASAP7_75t_L g686 ( .A(n_559), .B(n_664), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_560), .B(n_585), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_560), .A2(n_572), .B1(n_682), .B2(n_683), .Y(n_681) );
OR2x2_ASAP7_75t_L g712 ( .A(n_560), .B(n_580), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g689 ( .A(n_563), .Y(n_689) );
AND2x2_ASAP7_75t_L g714 ( .A(n_563), .B(n_657), .Y(n_714) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_SL g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g578 ( .A(n_568), .B(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_577), .B1(n_581), .B2(n_584), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g645 ( .A(n_573), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_573), .B(n_613), .Y(n_680) );
AOI322xp5_ASAP7_75t_L g604 ( .A1(n_575), .A2(n_605), .A3(n_607), .B1(n_608), .B2(n_610), .C1(n_611), .C2(n_615), .Y(n_604) );
INVxp67_ASAP7_75t_L g598 ( .A(n_576), .Y(n_598) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_578), .A2(n_583), .B1(n_600), .B2(n_602), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_579), .B(n_592), .Y(n_679) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_580), .B(n_618), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_580), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g676 ( .A(n_582), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NAND3xp33_ASAP7_75t_SL g587 ( .A(n_588), .B(n_604), .C(n_619), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_595), .B2(n_597), .C(n_599), .Y(n_588) );
AND2x2_ASAP7_75t_L g595 ( .A(n_591), .B(n_596), .Y(n_595) );
INVx3_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g605 ( .A(n_596), .B(n_606), .Y(n_605) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_598), .Y(n_677) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_603), .B(n_617), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_606), .B(n_664), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_607), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g682 ( .A(n_610), .Y(n_682) );
AND2x2_ASAP7_75t_L g697 ( .A(n_610), .B(n_674), .Y(n_697) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g691 ( .A1(n_621), .A2(n_692), .B(n_698), .C(n_706), .Y(n_691) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g660 ( .A(n_631), .B(n_661), .Y(n_660) );
NAND2x1_ASAP7_75t_SL g702 ( .A(n_632), .B(n_703), .Y(n_702) );
CKINVDCx16_ASAP7_75t_R g672 ( .A(n_635), .Y(n_672) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g667 ( .A(n_641), .Y(n_667) );
AND2x2_ASAP7_75t_L g671 ( .A(n_641), .B(n_657), .Y(n_671) );
NOR5xp2_ASAP7_75t_L g642 ( .A(n_643), .B(n_658), .C(n_675), .D(n_681), .E(n_684), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_646), .B2(n_648), .C(n_650), .Y(n_643) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_647), .B(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g673 ( .A(n_657), .B(n_674), .Y(n_673) );
OAI221xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_662), .B1(n_663), .B2(n_665), .C(n_668), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g711 ( .A(n_671), .Y(n_711) );
AOI211xp5_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_687), .B(n_689), .C(n_690), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
CKINVDCx14_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
CKINVDCx14_ASAP7_75t_R g726 ( .A(n_723), .Y(n_726) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx3_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
endmodule