module fake_netlist_6_4338_n_1725 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1725);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1725;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_66),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_27),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_84),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_78),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_67),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_31),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_28),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_123),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_90),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_110),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_17),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_10),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_89),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_44),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_114),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_77),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_43),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_101),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_18),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_4),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_97),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_44),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_46),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_103),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_61),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_65),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_50),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_85),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_34),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_7),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_36),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_137),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_25),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_7),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_138),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_45),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_56),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_68),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_33),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_43),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_24),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_106),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_129),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_38),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_25),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_105),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_39),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_17),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_38),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_73),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_14),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_80),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_20),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_71),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_29),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_11),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_93),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_36),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_41),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_0),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_48),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_95),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_72),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_98),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_99),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_63),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_113),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_26),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_30),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_50),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_116),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_124),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_39),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_94),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_145),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_142),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_55),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_2),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_131),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_28),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_75),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_108),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_57),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_54),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_51),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_60),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_121),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_22),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_32),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_23),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_52),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_37),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_76),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_119),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_23),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_136),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_14),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_70),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_6),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_37),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_3),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_12),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_62),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_19),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_52),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_143),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_53),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_26),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_40),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_40),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_45),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_10),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_24),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_74),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_16),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_196),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_156),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_280),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_196),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_196),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_231),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_231),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_169),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_161),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_161),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_212),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_178),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_178),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_181),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_158),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_255),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_181),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_159),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_185),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_185),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_192),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_160),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_192),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_163),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_255),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_164),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_206),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_232),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_259),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_165),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_206),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_207),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_207),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_211),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_215),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_167),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_223),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_215),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_220),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_168),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_220),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_221),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_171),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_172),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_221),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_259),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_173),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_230),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_230),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_241),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_175),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_241),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_243),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_243),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_252),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_252),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_176),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_277),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_254),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_177),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

NOR2x1_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_166),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_371),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_332),
.B(n_308),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_312),
.A2(n_276),
.B1(n_306),
.B2(n_238),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_166),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_318),
.A2(n_254),
.B1(n_216),
.B2(n_228),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_313),
.B(n_319),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_327),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_344),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_380),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_319),
.B(n_205),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_341),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_311),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_341),
.B(n_179),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_318),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_331),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_341),
.B(n_205),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_379),
.A2(n_236),
.B1(n_301),
.B2(n_293),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_346),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_157),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_346),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_346),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_320),
.B(n_208),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_350),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_357),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_329),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_320),
.B(n_208),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_350),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_330),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_366),
.B(n_217),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_366),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_330),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_335),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_326),
.B(n_180),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_354),
.B(n_223),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_322),
.B(n_326),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_334),
.B(n_287),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_336),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_322),
.B(n_217),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_338),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_340),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_326),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_438),
.B(n_342),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_418),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_438),
.B(n_347),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_407),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_418),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_420),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_409),
.B(n_356),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_421),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_413),
.B(n_360),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_364),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_333),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_421),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_385),
.B(n_367),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_413),
.B(n_377),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_443),
.B(n_287),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_420),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_191),
.Y(n_471)
);

CKINVDCx11_ASAP7_75t_R g472 ( 
.A(n_400),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_420),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_399),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_421),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_443),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_444),
.B(n_287),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_420),
.Y(n_479)
);

AO22x2_ASAP7_75t_L g480 ( 
.A1(n_395),
.A2(n_301),
.B1(n_293),
.B2(n_290),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_424),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_444),
.B(n_287),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_SL g484 ( 
.A(n_440),
.B(n_345),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_420),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_424),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_407),
.Y(n_492)
);

AND2x2_ASAP7_75t_SL g493 ( 
.A(n_393),
.B(n_229),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g494 ( 
.A(n_387),
.B(n_184),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_416),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_411),
.B(n_247),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_411),
.B(n_187),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_393),
.B(n_343),
.C(n_333),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_416),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_385),
.B(n_188),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_416),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_432),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_439),
.B(n_396),
.Y(n_506)
);

OAI22xp33_ASAP7_75t_SL g507 ( 
.A1(n_391),
.A2(n_266),
.B1(n_281),
.B2(n_273),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_416),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_396),
.B(n_189),
.Y(n_510)
);

BUFx6f_ASAP7_75t_SL g511 ( 
.A(n_431),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_L g512 ( 
.A1(n_395),
.A2(n_345),
.B1(n_359),
.B2(n_244),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_404),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_432),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_396),
.B(n_343),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_433),
.Y(n_521)
);

BUFx8_ASAP7_75t_SL g522 ( 
.A(n_400),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_L g524 ( 
.A(n_393),
.B(n_190),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_404),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_431),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_391),
.B(n_370),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

INVx8_ASAP7_75t_L g531 ( 
.A(n_406),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_406),
.B(n_193),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_406),
.A2(n_373),
.B1(n_370),
.B2(n_288),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_423),
.B(n_428),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_412),
.B(n_194),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_423),
.B(n_199),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_412),
.B(n_373),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_423),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_386),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_428),
.A2(n_290),
.B1(n_288),
.B2(n_285),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_428),
.A2(n_442),
.B1(n_417),
.B2(n_427),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_422),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_410),
.A2(n_239),
.B1(n_245),
.B2(n_307),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_422),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_410),
.B(n_284),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_422),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_442),
.B(n_337),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_410),
.A2(n_258),
.B1(n_174),
.B2(n_197),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_442),
.B(n_337),
.Y(n_551)
);

NAND3xp33_ASAP7_75t_L g552 ( 
.A(n_427),
.B(n_246),
.C(n_229),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_382),
.Y(n_553)
);

INVx8_ASAP7_75t_L g554 ( 
.A(n_422),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_427),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_417),
.A2(n_225),
.B1(n_203),
.B2(n_253),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_429),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_382),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_429),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_384),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_429),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_384),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_425),
.B(n_202),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_390),
.B(n_162),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_390),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_383),
.B(n_204),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_398),
.B(n_170),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_387),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_L g570 ( 
.A(n_429),
.B(n_209),
.Y(n_570)
);

AND3x2_ASAP7_75t_L g571 ( 
.A(n_398),
.B(n_256),
.C(n_246),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_429),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_425),
.B(n_213),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_429),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_414),
.A2(n_309),
.B1(n_285),
.B2(n_277),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_429),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_402),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_408),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_386),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_414),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_392),
.B(n_214),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_392),
.B(n_224),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_402),
.B(n_223),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_441),
.B(n_227),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_415),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_419),
.A2(n_234),
.B1(n_218),
.B2(n_305),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_408),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_441),
.B(n_235),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_408),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_408),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_415),
.A2(n_426),
.B1(n_436),
.B2(n_435),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_408),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_426),
.A2(n_309),
.B1(n_257),
.B2(n_260),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_493),
.B(n_441),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_493),
.B(n_441),
.Y(n_595)
);

CKINVDCx14_ASAP7_75t_R g596 ( 
.A(n_472),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_529),
.B(n_242),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_537),
.B(n_182),
.Y(n_598)
);

BUFx8_ASAP7_75t_L g599 ( 
.A(n_577),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_464),
.B(n_399),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_493),
.A2(n_257),
.B1(n_256),
.B2(n_295),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_539),
.B(n_445),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_462),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_560),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_539),
.B(n_441),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_539),
.B(n_441),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_506),
.B(n_441),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_534),
.B(n_445),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_525),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_506),
.B(n_441),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_496),
.B(n_445),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_471),
.B(n_445),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_484),
.A2(n_524),
.B1(n_477),
.B2(n_517),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_531),
.B(n_248),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_531),
.B(n_445),
.Y(n_617)
);

BUFx8_ASAP7_75t_L g618 ( 
.A(n_577),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_562),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_558),
.B(n_445),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_498),
.A2(n_260),
.B1(n_295),
.B2(n_281),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_498),
.B(n_183),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_566),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_464),
.B(n_419),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_558),
.B(n_446),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_525),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_542),
.B(n_249),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_457),
.B(n_430),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_580),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_462),
.B(n_419),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_446),
.B(n_445),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_446),
.B(n_445),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_446),
.B(n_383),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_463),
.B(n_186),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_531),
.A2(n_271),
.B1(n_262),
.B2(n_264),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_467),
.A2(n_251),
.B1(n_299),
.B2(n_291),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_551),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_551),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_531),
.B(n_451),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_L g643 ( 
.A1(n_583),
.A2(n_266),
.B1(n_271),
.B2(n_262),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_585),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_451),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_453),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_531),
.B(n_383),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_480),
.A2(n_264),
.B1(n_270),
.B2(n_269),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_548),
.B(n_250),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_453),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_497),
.B(n_548),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_466),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_546),
.B(n_261),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_532),
.B(n_536),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_555),
.B(n_383),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_555),
.B(n_383),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_513),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_466),
.B(n_394),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_522),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_483),
.B(n_394),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_510),
.B(n_195),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_483),
.B(n_394),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_535),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_481),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_491),
.Y(n_666)
);

AOI221xp5_ASAP7_75t_L g667 ( 
.A1(n_512),
.A2(n_233),
.B1(n_198),
.B2(n_200),
.C(n_201),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_491),
.B(n_274),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_474),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_492),
.A2(n_282),
.B1(n_270),
.B2(n_273),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_571),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_492),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_495),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_447),
.B(n_210),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_495),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_500),
.B(n_394),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_500),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_533),
.B(n_226),
.C(n_303),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_502),
.B(n_503),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_502),
.B(n_269),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_503),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_569),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_505),
.B(n_394),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_505),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_509),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_509),
.B(n_434),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_518),
.B(n_434),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_518),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_523),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_523),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_507),
.A2(n_430),
.B(n_434),
.C(n_369),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_526),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_526),
.B(n_388),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_527),
.B(n_388),
.Y(n_694)
);

BUFx6f_ASAP7_75t_SL g695 ( 
.A(n_569),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_450),
.A2(n_403),
.B1(n_388),
.B2(n_381),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_527),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_520),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_480),
.A2(n_223),
.B1(n_403),
.B2(n_349),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_520),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_449),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_456),
.B(n_339),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_567),
.B(n_403),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_452),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_452),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_507),
.B(n_408),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_454),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_454),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_458),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_481),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_565),
.B(n_408),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_591),
.A2(n_219),
.B1(n_302),
.B2(n_300),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_568),
.B(n_408),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_455),
.B(n_473),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_458),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_538),
.B(n_386),
.Y(n_716)
);

NOR2x1p5_ASAP7_75t_L g717 ( 
.A(n_553),
.B(n_222),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_459),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_494),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_455),
.B(n_381),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_544),
.B(n_237),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_455),
.B(n_381),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_481),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_501),
.A2(n_240),
.B1(n_265),
.B2(n_267),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_455),
.B(n_381),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_456),
.B(n_339),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_473),
.B(n_389),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_541),
.B(n_348),
.Y(n_728)
);

INVx8_ASAP7_75t_L g729 ( 
.A(n_553),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_473),
.B(n_389),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_473),
.B(n_389),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_460),
.B(n_58),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_469),
.B(n_268),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_485),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_586),
.A2(n_272),
.B1(n_275),
.B2(n_278),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_478),
.B(n_279),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_511),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_552),
.A2(n_405),
.B(n_401),
.C(n_397),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_461),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_552),
.A2(n_405),
.B(n_401),
.C(n_397),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_487),
.B(n_389),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_461),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_487),
.B(n_397),
.Y(n_743)
);

BUFx8_ASAP7_75t_L g744 ( 
.A(n_553),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_456),
.B(n_348),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_511),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_480),
.A2(n_593),
.B1(n_575),
.B2(n_511),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_482),
.B(n_283),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_487),
.B(n_397),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_SL g750 ( 
.A1(n_586),
.A2(n_286),
.B1(n_289),
.B2(n_292),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_487),
.B(n_401),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_538),
.B(n_386),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_559),
.B(n_386),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_485),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_559),
.B(n_386),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_549),
.B(n_351),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_556),
.B(n_351),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_456),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_489),
.B(n_401),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_468),
.B(n_352),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_561),
.B(n_386),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_554),
.A2(n_386),
.B(n_405),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_485),
.Y(n_763)
);

XOR2x2_ASAP7_75t_L g764 ( 
.A(n_733),
.B(n_581),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_596),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_700),
.B(n_659),
.Y(n_766)
);

BUFx4f_ASAP7_75t_L g767 ( 
.A(n_729),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_651),
.B(n_489),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_669),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_598),
.B(n_489),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_669),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_700),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_621),
.A2(n_582),
.B(n_588),
.C(n_584),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_657),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_700),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_615),
.A2(n_570),
.B1(n_563),
.B2(n_573),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_598),
.B(n_489),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_645),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_646),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_650),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_636),
.B(n_499),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_729),
.B(n_569),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_636),
.B(n_499),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_652),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_666),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_672),
.Y(n_786)
);

AO21x1_ASAP7_75t_L g787 ( 
.A1(n_595),
.A2(n_574),
.B(n_561),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_729),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_600),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_603),
.B(n_641),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_594),
.A2(n_554),
.B(n_479),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_640),
.B(n_499),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_601),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_647),
.A2(n_554),
.B(n_479),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_610),
.Y(n_795)
);

BUFx8_ASAP7_75t_L g796 ( 
.A(n_695),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_640),
.B(n_499),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_601),
.B(n_530),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_702),
.B(n_569),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_673),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_675),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_677),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_681),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_621),
.A2(n_355),
.B1(n_358),
.B2(n_361),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_684),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_599),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_685),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_700),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_625),
.A2(n_574),
.B1(n_572),
.B2(n_576),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_648),
.A2(n_622),
.B1(n_628),
.B2(n_699),
.Y(n_810)
);

AND2x2_ASAP7_75t_SL g811 ( 
.A(n_648),
.B(n_543),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_624),
.B(n_353),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_654),
.A2(n_545),
.B1(n_530),
.B2(n_572),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_688),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_689),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_698),
.A2(n_545),
.B1(n_530),
.B2(n_576),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_604),
.B(n_530),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_659),
.B(n_543),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_692),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_660),
.B(n_353),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_697),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_605),
.B(n_545),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_611),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_726),
.B(n_355),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_745),
.B(n_358),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_758),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_627),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_739),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_619),
.B(n_545),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_595),
.A2(n_543),
.B1(n_547),
.B2(n_550),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_623),
.B(n_547),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_695),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_626),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_630),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_739),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_739),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_629),
.B(n_361),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_635),
.B(n_547),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_638),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_632),
.A2(n_554),
.B(n_479),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_644),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_599),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_622),
.B(n_550),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_608),
.B(n_550),
.Y(n_844)
);

NOR2x2_ASAP7_75t_L g845 ( 
.A(n_760),
.B(n_578),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_664),
.B(n_589),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_612),
.B(n_589),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_744),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_760),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_618),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_747),
.B(n_634),
.Y(n_851)
);

OAI22xp33_ASAP7_75t_L g852 ( 
.A1(n_757),
.A2(n_362),
.B1(n_365),
.B2(n_368),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_665),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_747),
.B(n_461),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_614),
.B(n_461),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_703),
.B(n_589),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_739),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_737),
.B(n_578),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_699),
.A2(n_362),
.B1(n_365),
.B2(n_368),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_737),
.B(n_587),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_742),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_613),
.B(n_461),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_679),
.B(n_470),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_710),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_742),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_693),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_694),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_597),
.B(n_589),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_668),
.A2(n_592),
.B1(n_590),
.B2(n_587),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_658),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_744),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_735),
.B(n_592),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_662),
.B(n_459),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_671),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_756),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_631),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_742),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_723),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_661),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_742),
.B(n_470),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_682),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_663),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_719),
.B(n_369),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_633),
.A2(n_554),
.B(n_479),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_728),
.A2(n_735),
.B1(n_721),
.B2(n_706),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_676),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_746),
.B(n_587),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_683),
.Y(n_888)
);

INVx5_ASAP7_75t_L g889 ( 
.A(n_746),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_690),
.Y(n_890)
);

AO22x1_ASAP7_75t_L g891 ( 
.A1(n_733),
.A2(n_372),
.B1(n_374),
.B2(n_375),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_736),
.B(n_748),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_711),
.B(n_470),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_618),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_701),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_SL g896 ( 
.A1(n_736),
.A2(n_372),
.B1(n_374),
.B2(n_375),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_704),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_728),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_748),
.B(n_376),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_606),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_705),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_620),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_734),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_754),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_763),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_607),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_609),
.A2(n_504),
.B(n_465),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_707),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_SL g909 ( 
.A(n_717),
.B(n_470),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_662),
.B(n_590),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_708),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_696),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_709),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_715),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_732),
.B(n_376),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_609),
.B(n_465),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_674),
.B(n_590),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_674),
.B(n_592),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_649),
.B(n_470),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_653),
.B(n_475),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_668),
.B(n_475),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_616),
.B(n_59),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_678),
.B(n_479),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_718),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_667),
.B(n_378),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_680),
.B(n_476),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_680),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_643),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_686),
.Y(n_929)
);

NAND2x1p5_ASAP7_75t_L g930 ( 
.A(n_642),
.B(n_557),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_712),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_SL g932 ( 
.A1(n_750),
.A2(n_378),
.B1(n_564),
.B2(n_557),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_706),
.A2(n_514),
.B1(n_476),
.B2(n_508),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_687),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_655),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_656),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_724),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_713),
.B(n_488),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_643),
.B(n_557),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_642),
.A2(n_557),
.B1(n_564),
.B2(n_515),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_720),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_670),
.B(n_0),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_602),
.B(n_515),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_602),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_637),
.A2(n_557),
.B1(n_564),
.B2(n_514),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_617),
.A2(n_564),
.B(n_528),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_714),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_716),
.B(n_564),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_877),
.A2(n_617),
.B(n_751),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_877),
.A2(n_730),
.B(n_722),
.Y(n_950)
);

AO21x2_ASAP7_75t_L g951 ( 
.A1(n_843),
.A2(n_893),
.B(n_777),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_SL g952 ( 
.A(n_892),
.B(n_691),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_789),
.B(n_639),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_885),
.B(n_716),
.C(n_761),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_875),
.A2(n_931),
.B(n_937),
.C(n_812),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_877),
.A2(n_725),
.B(n_727),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_836),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_836),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_826),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_780),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_866),
.B(n_731),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_SL g962 ( 
.A1(n_917),
.A2(n_762),
.B(n_749),
.C(n_759),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_877),
.A2(n_743),
.B(n_741),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_925),
.A2(n_740),
.B(n_738),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_791),
.A2(n_761),
.B(n_755),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_867),
.B(n_755),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_810),
.A2(n_753),
.B(n_752),
.C(n_508),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_786),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_781),
.A2(n_753),
.B(n_752),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_789),
.B(n_504),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_899),
.B(n_516),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_775),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_764),
.A2(n_516),
.B1(n_488),
.B2(n_521),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_876),
.B(n_490),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_783),
.A2(n_528),
.B(n_579),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_799),
.B(n_519),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_786),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_824),
.B(n_490),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_801),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_771),
.B(n_1),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_769),
.B(n_9),
.Y(n_981)
);

OA21x2_ASAP7_75t_L g982 ( 
.A1(n_787),
.A2(n_521),
.B(n_519),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_769),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_825),
.B(n_486),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_801),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_774),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_790),
.B(n_486),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_934),
.B(n_486),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_770),
.A2(n_528),
.B(n_540),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_R g990 ( 
.A(n_765),
.B(n_100),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_768),
.A2(n_528),
.B(n_579),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_810),
.A2(n_885),
.B1(n_811),
.B2(n_939),
.Y(n_992)
);

BUFx8_ASAP7_75t_SL g993 ( 
.A(n_842),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_825),
.B(n_405),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_788),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_776),
.A2(n_528),
.B1(n_540),
.B2(n_579),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_811),
.A2(n_528),
.B1(n_13),
.B2(n_15),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_894),
.B(n_579),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_883),
.B(n_9),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_898),
.B(n_15),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_938),
.A2(n_847),
.B(n_893),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_794),
.A2(n_540),
.B(n_448),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_SL g1003 ( 
.A1(n_917),
.A2(n_96),
.B(n_155),
.C(n_154),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_836),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_836),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_807),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_773),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_1007)
);

INVxp67_ASAP7_75t_SL g1008 ( 
.A(n_857),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_853),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_833),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_856),
.A2(n_540),
.B(n_448),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_775),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_900),
.B(n_21),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_840),
.A2(n_448),
.B(n_102),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_851),
.A2(n_448),
.B1(n_30),
.B2(n_35),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_900),
.B(n_21),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_788),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_795),
.B(n_35),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_884),
.A2(n_104),
.B(n_148),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_851),
.A2(n_152),
.B(n_92),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_870),
.B(n_91),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_910),
.A2(n_107),
.B(n_140),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_833),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_910),
.A2(n_88),
.B(n_133),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_872),
.A2(n_42),
.B(n_46),
.C(n_47),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_848),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_837),
.B(n_87),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_806),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_912),
.A2(n_42),
.B1(n_47),
.B2(n_49),
.Y(n_1029)
);

NAND2xp33_ASAP7_75t_R g1030 ( 
.A(n_922),
.B(n_117),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_879),
.B(n_111),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_882),
.B(n_118),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_795),
.B(n_49),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_871),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_834),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_942),
.A2(n_51),
.B(n_53),
.C(n_64),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_912),
.A2(n_69),
.B1(n_79),
.B2(n_81),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_782),
.B(n_83),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_827),
.B(n_120),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_939),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_886),
.B(n_128),
.Y(n_1041)
);

NAND2x1p5_ASAP7_75t_L g1042 ( 
.A(n_889),
.B(n_130),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_837),
.B(n_144),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_827),
.B(n_849),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_873),
.A2(n_862),
.B(n_855),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_855),
.A2(n_862),
.B(n_918),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_806),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_857),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_853),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_874),
.B(n_823),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_932),
.A2(n_854),
.B1(n_798),
.B2(n_872),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_864),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_918),
.A2(n_927),
.B(n_923),
.C(n_888),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_854),
.A2(n_821),
.B1(n_805),
.B2(n_819),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_SL g1055 ( 
.A(n_793),
.B(n_896),
.C(n_881),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_906),
.B(n_935),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_909),
.A2(n_915),
.B1(n_923),
.B2(n_803),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_844),
.A2(n_818),
.B(n_863),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_820),
.B(n_834),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_864),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_857),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_796),
.Y(n_1062)
);

INVx3_ASAP7_75t_SL g1063 ( 
.A(n_832),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_928),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_878),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_778),
.A2(n_815),
.B1(n_800),
.B2(n_814),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_863),
.A2(n_919),
.B(n_846),
.C(n_909),
.Y(n_1067)
);

BUFx8_ASAP7_75t_L g1068 ( 
.A(n_850),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_889),
.B(n_839),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_841),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_845),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_852),
.A2(n_890),
.B(n_802),
.C(n_779),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_784),
.A2(n_785),
.B1(n_859),
.B2(n_841),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_857),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_782),
.B(n_889),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_844),
.A2(n_818),
.B(n_797),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_792),
.A2(n_868),
.B(n_919),
.Y(n_1077)
);

NOR2xp67_ASAP7_75t_SL g1078 ( 
.A(n_889),
.B(n_865),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_845),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_767),
.B(n_772),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_906),
.B(n_935),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_915),
.A2(n_928),
.B1(n_887),
.B2(n_860),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_921),
.A2(n_830),
.B(n_880),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_878),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_880),
.A2(n_941),
.B(n_936),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_905),
.Y(n_1086)
);

INVxp67_ASAP7_75t_SL g1087 ( 
.A(n_865),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_941),
.A2(n_936),
.B(n_946),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_929),
.B(n_902),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_793),
.B(n_859),
.C(n_891),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_R g1091 ( 
.A(n_767),
.B(n_772),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_1038),
.B(n_782),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_992),
.A2(n_846),
.A3(n_809),
.B(n_944),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1077),
.A2(n_916),
.B(n_920),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_1004),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1088),
.A2(n_907),
.B(n_930),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_959),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_986),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_965),
.A2(n_930),
.B(n_838),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_960),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_983),
.B(n_820),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1090),
.A2(n_895),
.B(n_897),
.C(n_908),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_955),
.A2(n_901),
.B(n_913),
.C(n_911),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1029),
.A2(n_804),
.B(n_852),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1051),
.A2(n_804),
.B1(n_766),
.B2(n_933),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1058),
.A2(n_1085),
.B(n_1076),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_995),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_1067),
.A2(n_869),
.B(n_831),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1071),
.B(n_820),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_SL g1110 ( 
.A1(n_1020),
.A2(n_829),
.B(n_822),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_972),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1055),
.A2(n_924),
.B1(n_914),
.B2(n_911),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1001),
.A2(n_865),
.B(n_817),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1083),
.A2(n_813),
.B(n_933),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_999),
.B(n_924),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1056),
.B(n_902),
.Y(n_1116)
);

AO21x1_ASAP7_75t_L g1117 ( 
.A1(n_1051),
.A2(n_1054),
.B(n_997),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_1046),
.A2(n_816),
.B(n_914),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1045),
.A2(n_943),
.B(n_940),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_1007),
.A2(n_926),
.B(n_905),
.C(n_808),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_997),
.A2(n_766),
.B1(n_913),
.B2(n_865),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1015),
.A2(n_945),
.B1(n_947),
.B2(n_835),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_SL g1123 ( 
.A1(n_1020),
.A2(n_922),
.B(n_947),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1053),
.A2(n_887),
.B(n_860),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1059),
.B(n_858),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_1078),
.Y(n_1126)
);

OAI22x1_ASAP7_75t_L g1127 ( 
.A1(n_1082),
.A2(n_858),
.B1(n_887),
.B2(n_860),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1072),
.A2(n_858),
.B(n_903),
.C(n_904),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_1054),
.A2(n_947),
.A3(n_948),
.B(n_861),
.Y(n_1129)
);

CKINVDCx6p67_ASAP7_75t_R g1130 ( 
.A(n_1063),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_1021),
.A2(n_828),
.B(n_835),
.C(n_861),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_957),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_968),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_952),
.A2(n_903),
.B(n_904),
.C(n_948),
.Y(n_1134)
);

OAI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1030),
.A2(n_828),
.B1(n_1079),
.B2(n_1071),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_964),
.A2(n_969),
.B(n_952),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1081),
.B(n_970),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_949),
.A2(n_950),
.B(n_956),
.Y(n_1138)
);

INVxp67_ASAP7_75t_SL g1139 ( 
.A(n_1089),
.Y(n_1139)
);

NOR4xp25_ASAP7_75t_L g1140 ( 
.A(n_1025),
.B(n_1036),
.C(n_1040),
.D(n_1013),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1017),
.Y(n_1141)
);

NOR2x1_ASAP7_75t_SL g1142 ( 
.A(n_1004),
.B(n_1038),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_967),
.A2(n_1073),
.A3(n_1032),
.B(n_1031),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1081),
.B(n_961),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_977),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_971),
.A2(n_962),
.B(n_951),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_963),
.A2(n_1014),
.B(n_975),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1028),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_961),
.B(n_966),
.Y(n_1149)
);

NAND3x1_ASAP7_75t_L g1150 ( 
.A(n_981),
.B(n_1018),
.C(n_1033),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_966),
.B(n_985),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1002),
.A2(n_989),
.B(n_991),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_979),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_SL g1154 ( 
.A1(n_1021),
.A2(n_1032),
.B(n_1031),
.Y(n_1154)
);

AOI211x1_ASAP7_75t_L g1155 ( 
.A1(n_1066),
.A2(n_1073),
.B(n_1016),
.C(n_953),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1066),
.B(n_987),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_957),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1006),
.B(n_1010),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1023),
.B(n_1035),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1009),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_957),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_951),
.A2(n_978),
.B(n_1041),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_1044),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1041),
.A2(n_1004),
.B(n_1057),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1000),
.B(n_980),
.C(n_1024),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1047),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1050),
.B(n_974),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1011),
.A2(n_1019),
.B(n_982),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_SL g1169 ( 
.A1(n_1022),
.A2(n_1040),
.B(n_1037),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1062),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1070),
.B(n_1050),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1075),
.A2(n_1042),
.B(n_1038),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_982),
.A2(n_988),
.B(n_1069),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_994),
.B(n_1084),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1027),
.A2(n_1043),
.B1(n_976),
.B2(n_984),
.C(n_1039),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1064),
.B(n_1091),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_954),
.A2(n_973),
.B(n_1086),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1004),
.A2(n_996),
.B(n_1008),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1049),
.A2(n_1065),
.A3(n_1060),
.B(n_1052),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1042),
.A2(n_972),
.B(n_1012),
.Y(n_1180)
);

AO31x2_ASAP7_75t_L g1181 ( 
.A1(n_1003),
.A2(n_1087),
.A3(n_958),
.B(n_1048),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_990),
.B(n_1034),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1012),
.B(n_1075),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_958),
.Y(n_1184)
);

NOR2xp67_ASAP7_75t_L g1185 ( 
.A(n_1026),
.B(n_958),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_SL g1186 ( 
.A1(n_1080),
.A2(n_1005),
.B(n_1048),
.C(n_1061),
.Y(n_1186)
);

BUFx10_ASAP7_75t_L g1187 ( 
.A(n_1005),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1005),
.A2(n_1048),
.B(n_1061),
.C(n_1074),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1061),
.A2(n_1074),
.B(n_998),
.C(n_1068),
.Y(n_1189)
);

AO21x2_ASAP7_75t_L g1190 ( 
.A1(n_1074),
.A2(n_998),
.B(n_1068),
.Y(n_1190)
);

OAI22x1_ASAP7_75t_L g1191 ( 
.A1(n_993),
.A2(n_892),
.B1(n_477),
.B2(n_615),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_998),
.B(n_892),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_992),
.A2(n_601),
.B1(n_810),
.B2(n_885),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_992),
.A2(n_892),
.B1(n_764),
.B2(n_1090),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_960),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1077),
.A2(n_531),
.B(n_843),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1056),
.B(n_892),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_992),
.A2(n_892),
.B(n_477),
.C(n_615),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1088),
.A2(n_965),
.B(n_1058),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_957),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_986),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_992),
.A2(n_892),
.B(n_477),
.C(n_615),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1056),
.B(n_892),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_983),
.B(n_789),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_972),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_992),
.A2(n_438),
.B1(n_583),
.B2(n_615),
.Y(n_1206)
);

NAND2xp33_ASAP7_75t_R g1207 ( 
.A(n_959),
.B(n_387),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_992),
.A2(n_997),
.B1(n_1090),
.B2(n_1051),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_959),
.B(n_669),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1071),
.B(n_327),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_992),
.A2(n_1051),
.A3(n_787),
.B(n_1053),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_992),
.A2(n_1051),
.B(n_1046),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_992),
.B(n_892),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_992),
.B(n_866),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_SL g1215 ( 
.A(n_1028),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_992),
.A2(n_601),
.B1(n_810),
.B2(n_885),
.Y(n_1216)
);

O2A1O1Ixp5_ASAP7_75t_SL g1217 ( 
.A1(n_992),
.A2(n_997),
.B(n_440),
.C(n_501),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_992),
.B(n_866),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1088),
.A2(n_965),
.B(n_1058),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1077),
.A2(n_531),
.B(n_843),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_SL g1221 ( 
.A1(n_1007),
.A2(n_992),
.B(n_1053),
.C(n_1031),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1088),
.A2(n_965),
.B(n_1058),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1067),
.A2(n_1046),
.B(n_1045),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_992),
.B(n_866),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_992),
.A2(n_1051),
.B(n_1046),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1059),
.B(n_898),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1088),
.A2(n_965),
.B(n_1058),
.Y(n_1227)
);

CKINVDCx8_ASAP7_75t_R g1228 ( 
.A(n_959),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1197),
.B(n_1203),
.Y(n_1229)
);

AO21x2_ASAP7_75t_L g1230 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1212),
.Y(n_1230)
);

AOI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1206),
.A2(n_1194),
.B1(n_1216),
.B2(n_1193),
.C(n_1140),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1132),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1139),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1208),
.B(n_1144),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1100),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1133),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1150),
.A2(n_1202),
.B1(n_1198),
.B2(n_1193),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1201),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1152),
.A2(n_1138),
.B(n_1147),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1153),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1212),
.A2(n_1225),
.B(n_1154),
.Y(n_1241)
);

INVxp67_ASAP7_75t_SL g1242 ( 
.A(n_1204),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1220),
.A2(n_1216),
.B(n_1213),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_R g1244 ( 
.A(n_1097),
.B(n_1182),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1134),
.A2(n_1214),
.B(n_1224),
.C(n_1218),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_1168),
.B(n_1222),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1208),
.B(n_1144),
.Y(n_1247)
);

BUFx2_ASAP7_75t_SL g1248 ( 
.A(n_1215),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1137),
.B(n_1167),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1199),
.A2(n_1219),
.B(n_1227),
.Y(n_1250)
);

AOI221xp5_ASAP7_75t_L g1251 ( 
.A1(n_1140),
.A2(n_1104),
.B1(n_1191),
.B2(n_1221),
.C(n_1225),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1165),
.A2(n_1217),
.B(n_1164),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1172),
.B(n_1155),
.Y(n_1253)
);

CKINVDCx8_ASAP7_75t_R g1254 ( 
.A(n_1226),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1132),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1106),
.A2(n_1096),
.B(n_1113),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1115),
.B(n_1149),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1149),
.B(n_1116),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1095),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1130),
.Y(n_1260)
);

AOI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1094),
.A2(n_1178),
.B(n_1169),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1119),
.A2(n_1114),
.B(n_1173),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1210),
.B(n_1163),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1107),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1207),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1129),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1214),
.B(n_1218),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1136),
.A2(n_1180),
.B(n_1124),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1165),
.B(n_1175),
.Y(n_1269)
);

AOI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1104),
.A2(n_1117),
.B1(n_1136),
.B2(n_1105),
.C(n_1109),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1098),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1101),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1187),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1105),
.A2(n_1135),
.B1(n_1175),
.B2(n_1156),
.C(n_1102),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1171),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1095),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1195),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1192),
.A2(n_1226),
.B1(n_1127),
.B2(n_1125),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1110),
.A2(n_1123),
.B(n_1131),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1111),
.B(n_1205),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1190),
.B(n_1142),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1092),
.A2(n_1209),
.B1(n_1112),
.B2(n_1176),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1160),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1228),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1129),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1141),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1124),
.A2(n_1223),
.B(n_1118),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1112),
.A2(n_1103),
.B(n_1122),
.C(n_1121),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1128),
.A2(n_1151),
.B(n_1122),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1151),
.B(n_1174),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1174),
.B(n_1145),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1223),
.A2(n_1118),
.B(n_1121),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1108),
.A2(n_1177),
.B(n_1159),
.Y(n_1293)
);

OAI221xp5_ASAP7_75t_L g1294 ( 
.A1(n_1092),
.A2(n_1185),
.B1(n_1189),
.B2(n_1166),
.C(n_1183),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1120),
.A2(n_1092),
.B(n_1126),
.C(n_1158),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1111),
.B(n_1205),
.Y(n_1296)
);

NAND2x1p5_ASAP7_75t_L g1297 ( 
.A(n_1177),
.B(n_1161),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1148),
.B(n_1184),
.C(n_1188),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1190),
.Y(n_1299)
);

OAI22x1_ASAP7_75t_L g1300 ( 
.A1(n_1211),
.A2(n_1143),
.B1(n_1093),
.B2(n_1181),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1143),
.A2(n_1211),
.B(n_1181),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1132),
.B(n_1157),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1143),
.A2(n_1211),
.B(n_1181),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1186),
.A2(n_1093),
.B(n_1187),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1093),
.A2(n_1157),
.B(n_1161),
.Y(n_1305)
);

AOI22x1_ASAP7_75t_L g1306 ( 
.A1(n_1200),
.A2(n_892),
.B1(n_1191),
.B2(n_1154),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1215),
.A2(n_1206),
.B(n_892),
.C(n_1202),
.Y(n_1307)
);

CKINVDCx6p67_ASAP7_75t_R g1308 ( 
.A(n_1170),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1200),
.A2(n_1117),
.A3(n_1216),
.B(n_1193),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1201),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1194),
.B(n_1208),
.Y(n_1311)
);

AOI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1164),
.A2(n_1146),
.B(n_1196),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1095),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1225),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1193),
.A2(n_1216),
.B(n_992),
.C(n_1202),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1100),
.Y(n_1316)
);

AO21x1_ASAP7_75t_L g1317 ( 
.A1(n_1193),
.A2(n_1216),
.B(n_992),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1179),
.Y(n_1318)
);

AO21x2_ASAP7_75t_L g1319 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1225),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1201),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1212),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1204),
.Y(n_1322)
);

CKINVDCx16_ASAP7_75t_R g1323 ( 
.A(n_1207),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1206),
.A2(n_892),
.B(n_1202),
.C(n_1198),
.Y(n_1324)
);

CKINVDCx8_ASAP7_75t_R g1325 ( 
.A(n_1097),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1212),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1225),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1198),
.A2(n_892),
.B(n_1202),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1152),
.A2(n_1138),
.B(n_1147),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1095),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1198),
.A2(n_892),
.B(n_1202),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1179),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1100),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1197),
.B(n_1203),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_SL g1335 ( 
.A1(n_1142),
.A2(n_1123),
.B(n_1154),
.Y(n_1335)
);

OAI221xp5_ASAP7_75t_L g1336 ( 
.A1(n_1194),
.A2(n_484),
.B1(n_438),
.B2(n_477),
.C(n_764),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1197),
.B(n_1203),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1197),
.B(n_1203),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1179),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1179),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1152),
.A2(n_1138),
.B(n_1147),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1132),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1152),
.A2(n_1138),
.B(n_1147),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1194),
.A2(n_892),
.B1(n_764),
.B2(n_1206),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1198),
.A2(n_892),
.B(n_1202),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1198),
.A2(n_892),
.B(n_1202),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1152),
.A2(n_1138),
.B(n_1147),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1100),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1336),
.A2(n_1344),
.B1(n_1237),
.B2(n_1231),
.C(n_1251),
.Y(n_1349)
);

O2A1O1Ixp5_ASAP7_75t_L g1350 ( 
.A1(n_1269),
.A2(n_1252),
.B(n_1317),
.C(n_1243),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1272),
.B(n_1299),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1233),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1265),
.A2(n_1323),
.B1(n_1315),
.B2(n_1263),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1299),
.B(n_1281),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1249),
.B(n_1311),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1242),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1265),
.A2(n_1315),
.B1(n_1278),
.B2(n_1254),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1257),
.B(n_1334),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_SL g1359 ( 
.A1(n_1328),
.A2(n_1346),
.B(n_1345),
.C(n_1331),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1325),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1264),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1322),
.B(n_1234),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1254),
.A2(n_1294),
.B1(n_1270),
.B2(n_1253),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1235),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1292),
.A2(n_1303),
.B(n_1301),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1275),
.B(n_1258),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1253),
.A2(n_1298),
.B1(n_1282),
.B2(n_1288),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1324),
.A2(n_1307),
.B(n_1288),
.C(n_1274),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1290),
.B(n_1247),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1236),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1238),
.Y(n_1372)
);

NOR2xp67_ASAP7_75t_L g1373 ( 
.A(n_1271),
.B(n_1273),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1286),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1291),
.B(n_1267),
.Y(n_1375)
);

OAI31xp33_ASAP7_75t_L g1376 ( 
.A1(n_1269),
.A2(n_1320),
.A3(n_1238),
.B(n_1310),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_SL g1377 ( 
.A1(n_1306),
.A2(n_1317),
.B(n_1261),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1267),
.B(n_1283),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1310),
.B(n_1320),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1325),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1295),
.A2(n_1245),
.B(n_1304),
.C(n_1335),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1240),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1253),
.A2(n_1259),
.B(n_1313),
.Y(n_1383)
);

O2A1O1Ixp5_ASAP7_75t_L g1384 ( 
.A1(n_1312),
.A2(n_1305),
.B(n_1340),
.C(n_1339),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1232),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1286),
.Y(n_1386)
);

INVx3_ASAP7_75t_SL g1387 ( 
.A(n_1284),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1253),
.A2(n_1260),
.B1(n_1248),
.B2(n_1284),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1277),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1259),
.A2(n_1330),
.B(n_1313),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1241),
.A2(n_1348),
.B(n_1333),
.C(n_1316),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1241),
.B(n_1309),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_SL g1393 ( 
.A1(n_1260),
.A2(n_1273),
.B1(n_1244),
.B2(n_1302),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1280),
.A2(n_1296),
.B1(n_1289),
.B2(n_1297),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1292),
.A2(n_1303),
.B(n_1301),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1287),
.A2(n_1293),
.B(n_1343),
.Y(n_1396)
);

AOI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1300),
.A2(n_1230),
.B1(n_1319),
.B2(n_1314),
.C(n_1327),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1232),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1296),
.A2(n_1289),
.B1(n_1276),
.B2(n_1308),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1309),
.B(n_1289),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1302),
.B(n_1276),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_L g1402 ( 
.A(n_1259),
.B(n_1313),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1287),
.A2(n_1293),
.B(n_1239),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1232),
.B(n_1342),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1308),
.A2(n_1330),
.B1(n_1266),
.B2(n_1285),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1232),
.Y(n_1406)
);

AND2x2_ASAP7_75t_SL g1407 ( 
.A(n_1266),
.B(n_1285),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1239),
.A2(n_1347),
.B(n_1343),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1255),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1330),
.A2(n_1342),
.B1(n_1255),
.B2(n_1326),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1255),
.A2(n_1342),
.B1(n_1321),
.B2(n_1318),
.Y(n_1411)
);

OAI31xp33_ASAP7_75t_L g1412 ( 
.A1(n_1332),
.A2(n_1279),
.A3(n_1321),
.B(n_1268),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1255),
.B(n_1268),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1262),
.B(n_1256),
.Y(n_1414)
);

AOI221x1_ASAP7_75t_SL g1415 ( 
.A1(n_1262),
.A2(n_1256),
.B1(n_1246),
.B2(n_1250),
.C(n_1329),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1246),
.B(n_1329),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1341),
.A2(n_1336),
.B1(n_1344),
.B2(n_1150),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1233),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1336),
.A2(n_1344),
.B1(n_1150),
.B2(n_1194),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1336),
.A2(n_1344),
.B1(n_1150),
.B2(n_1194),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1257),
.B(n_1229),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1252),
.A2(n_1292),
.B(n_1301),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1367),
.B(n_1370),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1392),
.B(n_1400),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_1356),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1363),
.B(n_1422),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1354),
.B(n_1413),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1349),
.A2(n_1419),
.B1(n_1420),
.B2(n_1353),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1422),
.B(n_1407),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1422),
.B(n_1407),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1416),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1351),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1397),
.A2(n_1384),
.B(n_1350),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1369),
.A2(n_1360),
.B1(n_1417),
.B2(n_1368),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1350),
.A2(n_1369),
.B(n_1414),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1359),
.A2(n_1381),
.B(n_1364),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1365),
.B(n_1382),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1352),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1418),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1366),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1418),
.B(n_1412),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1355),
.B(n_1395),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1371),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1395),
.B(n_1396),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1411),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1395),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1396),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1389),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1394),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1403),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1378),
.B(n_1421),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1391),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1408),
.B(n_1405),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1399),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1408),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1385),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1377),
.A2(n_1415),
.B(n_1358),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1401),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1443),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1438),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1431),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1428),
.A2(n_1357),
.B1(n_1388),
.B2(n_1393),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1442),
.B(n_1372),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1448),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1426),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1442),
.B(n_1404),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1426),
.B(n_1376),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1425),
.B(n_1379),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1432),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1426),
.B(n_1442),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1443),
.Y(n_1472)
);

BUFx4f_ASAP7_75t_SL g1473 ( 
.A(n_1457),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1439),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1424),
.B(n_1379),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1439),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1425),
.B(n_1373),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1424),
.B(n_1386),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1448),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1429),
.B(n_1385),
.Y(n_1480)
);

NAND2x1p5_ASAP7_75t_L g1481 ( 
.A(n_1435),
.B(n_1401),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1437),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1423),
.B(n_1387),
.Y(n_1483)
);

INVx8_ASAP7_75t_L g1484 ( 
.A(n_1437),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1423),
.B(n_1398),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1463),
.A2(n_1434),
.B1(n_1436),
.B2(n_1455),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1465),
.A2(n_1456),
.B(n_1447),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1467),
.B(n_1430),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1483),
.A2(n_1434),
.B1(n_1436),
.B2(n_1446),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1460),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1463),
.A2(n_1428),
.B1(n_1435),
.B2(n_1455),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1461),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1468),
.A2(n_1453),
.B1(n_1446),
.B2(n_1445),
.C(n_1450),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1453),
.C(n_1458),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1474),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1484),
.B(n_1383),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1468),
.A2(n_1445),
.B1(n_1450),
.B2(n_1452),
.C(n_1449),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1461),
.Y(n_1498)
);

NAND2xp33_ASAP7_75t_R g1499 ( 
.A(n_1470),
.B(n_1361),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1467),
.B(n_1427),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1474),
.Y(n_1501)
);

OAI211xp5_ASAP7_75t_L g1502 ( 
.A1(n_1477),
.A2(n_1435),
.B(n_1433),
.C(n_1452),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1481),
.A2(n_1435),
.B(n_1433),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1469),
.A2(n_1427),
.B1(n_1435),
.B2(n_1459),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1460),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1462),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1473),
.Y(n_1507)
);

OR2x6_ASAP7_75t_L g1508 ( 
.A(n_1484),
.B(n_1441),
.Y(n_1508)
);

AOI211xp5_ASAP7_75t_L g1509 ( 
.A1(n_1477),
.A2(n_1387),
.B(n_1441),
.C(n_1454),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1472),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1467),
.B(n_1427),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1479),
.A2(n_1451),
.B(n_1447),
.Y(n_1512)
);

OAI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1481),
.A2(n_1441),
.B1(n_1433),
.B2(n_1374),
.C(n_1454),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1480),
.B(n_1427),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1475),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1472),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1471),
.B(n_1424),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1490),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1507),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1508),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1503),
.A2(n_1440),
.B(n_1444),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1505),
.Y(n_1523)
);

BUFx4f_ASAP7_75t_L g1524 ( 
.A(n_1496),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1507),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1505),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1512),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1512),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1486),
.B(n_1433),
.C(n_1458),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1506),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1507),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1510),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1492),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1508),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1489),
.B(n_1362),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1510),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1494),
.A2(n_1451),
.B(n_1447),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1493),
.B(n_1475),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1517),
.B(n_1471),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1516),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1508),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1516),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1508),
.B(n_1482),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1491),
.A2(n_1449),
.B(n_1433),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1512),
.Y(n_1545)
);

AND2x6_ASAP7_75t_SL g1546 ( 
.A(n_1496),
.B(n_1380),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1508),
.B(n_1482),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1487),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1488),
.B(n_1471),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1521),
.B(n_1488),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1538),
.B(n_1493),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1518),
.B(n_1519),
.Y(n_1552)
);

NAND5xp2_ASAP7_75t_L g1553 ( 
.A(n_1535),
.B(n_1491),
.C(n_1509),
.D(n_1497),
.E(n_1502),
.Y(n_1553)
);

INVx3_ASAP7_75t_SL g1554 ( 
.A(n_1531),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1518),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1521),
.B(n_1534),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1519),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1534),
.B(n_1500),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1541),
.B(n_1500),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_1517),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1539),
.B(n_1494),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1523),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1541),
.B(n_1511),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1523),
.B(n_1497),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1528),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1533),
.B(n_1495),
.Y(n_1566)
);

AOI221x1_ASAP7_75t_L g1567 ( 
.A1(n_1529),
.A2(n_1503),
.B1(n_1507),
.B2(n_1485),
.C(n_1390),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1528),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1526),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1528),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1544),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1526),
.B(n_1501),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1543),
.B(n_1506),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1532),
.B(n_1466),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1520),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1543),
.B(n_1547),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1532),
.B(n_1466),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_L g1578 ( 
.A(n_1520),
.B(n_1513),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1528),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1536),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1549),
.B(n_1543),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1549),
.B(n_1511),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1515),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1540),
.B(n_1476),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1543),
.B(n_1514),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1544),
.B(n_1464),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1529),
.A2(n_1513),
.B1(n_1509),
.B2(n_1504),
.C(n_1476),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1545),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1540),
.B(n_1464),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1542),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1547),
.B(n_1514),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1551),
.B(n_1520),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1525),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1578),
.B(n_1547),
.Y(n_1594)
);

NOR2x1p5_ASAP7_75t_L g1595 ( 
.A(n_1575),
.B(n_1525),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1575),
.B(n_1525),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1566),
.B(n_1475),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1566),
.B(n_1478),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1564),
.B(n_1542),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1564),
.B(n_1561),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1575),
.B(n_1556),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1556),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1557),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1557),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1555),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1555),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1554),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1562),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1556),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1553),
.B(n_1525),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1587),
.B(n_1531),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1562),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1561),
.B(n_1583),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1578),
.B(n_1547),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1554),
.B(n_1531),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1558),
.B(n_1524),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1569),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1587),
.A2(n_1531),
.B1(n_1524),
.B2(n_1496),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1569),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1554),
.B(n_1531),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1580),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1580),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1560),
.B(n_1478),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1571),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1590),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1620),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1620),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1610),
.B(n_1550),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1619),
.A2(n_1571),
.B1(n_1586),
.B2(n_1524),
.C(n_1531),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1610),
.B(n_1550),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1605),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1602),
.B(n_1550),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1625),
.B(n_1560),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1611),
.A2(n_1553),
.B(n_1567),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1606),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_L g1637 ( 
.A(n_1611),
.B(n_1590),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_L g1638 ( 
.A(n_1600),
.B(n_1567),
.C(n_1586),
.Y(n_1638)
);

INVx4_ASAP7_75t_L g1639 ( 
.A(n_1607),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1608),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1612),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1595),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1600),
.A2(n_1524),
.B1(n_1537),
.B2(n_1563),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1594),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1609),
.B(n_1558),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1618),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1622),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1593),
.A2(n_1617),
.B1(n_1613),
.B2(n_1601),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1596),
.B(n_1559),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1563),
.Y(n_1651)
);

AOI211x1_ASAP7_75t_L g1652 ( 
.A1(n_1635),
.A2(n_1616),
.B(n_1621),
.C(n_1615),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1637),
.B(n_1603),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1627),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1639),
.B(n_1617),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1651),
.B(n_1597),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1638),
.A2(n_1599),
.B(n_1594),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1639),
.B(n_1615),
.Y(n_1658)
);

AOI222xp33_ASAP7_75t_L g1659 ( 
.A1(n_1629),
.A2(n_1631),
.B1(n_1649),
.B2(n_1630),
.C1(n_1628),
.C2(n_1643),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1642),
.B(n_1585),
.Y(n_1660)
);

AO21x1_ASAP7_75t_L g1661 ( 
.A1(n_1644),
.A2(n_1604),
.B(n_1599),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1648),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1634),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1645),
.B(n_1633),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1648),
.A2(n_1598),
.B1(n_1573),
.B2(n_1576),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1644),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1632),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1649),
.B(n_1623),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_L g1669 ( 
.A(n_1636),
.B(n_1626),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1640),
.B(n_1624),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1660),
.B(n_1650),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1669),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1659),
.A2(n_1643),
.B1(n_1646),
.B2(n_1647),
.Y(n_1673)
);

NAND2x1_ASAP7_75t_L g1674 ( 
.A(n_1658),
.B(n_1641),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1655),
.B(n_1583),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1663),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1652),
.B(n_1582),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1666),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1659),
.A2(n_1537),
.B1(n_1614),
.B2(n_1576),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1661),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1662),
.B(n_1582),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1546),
.Y(n_1682)
);

OAI322xp33_ASAP7_75t_L g1683 ( 
.A1(n_1680),
.A2(n_1657),
.A3(n_1668),
.B1(n_1653),
.B2(n_1654),
.C1(n_1667),
.C2(n_1670),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1679),
.A2(n_1653),
.B(n_1670),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1679),
.A2(n_1665),
.B1(n_1656),
.B2(n_1573),
.Y(n_1685)
);

OAI221xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1673),
.A2(n_1614),
.B1(n_1576),
.B2(n_1573),
.C(n_1588),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1681),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_SL g1688 ( 
.A(n_1673),
.B(n_1581),
.C(n_1572),
.D(n_1492),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1678),
.B(n_1581),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1682),
.A2(n_1499),
.B1(n_1591),
.B2(n_1572),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1674),
.Y(n_1691)
);

OAI21xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1685),
.A2(n_1672),
.B(n_1677),
.Y(n_1692)
);

AOI211xp5_ASAP7_75t_L g1693 ( 
.A1(n_1683),
.A2(n_1676),
.B(n_1675),
.C(n_1671),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1691),
.A2(n_1579),
.B(n_1568),
.Y(n_1694)
);

A2O1A1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1684),
.A2(n_1530),
.B(n_1522),
.C(n_1565),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1686),
.A2(n_1530),
.B(n_1522),
.C(n_1565),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1694),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1693),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1692),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1696),
.B(n_1689),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1695),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1693),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1699),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1700),
.B(n_1690),
.Y(n_1704)
);

NOR4xp25_ASAP7_75t_L g1705 ( 
.A(n_1698),
.B(n_1687),
.C(n_1688),
.D(n_1588),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1702),
.B(n_1552),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1697),
.A2(n_1579),
.B1(n_1570),
.B2(n_1568),
.C(n_1588),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1703),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1704),
.B(n_1701),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1706),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1708),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1709),
.B1(n_1708),
.B2(n_1710),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1705),
.B(n_1707),
.Y(n_1713)
);

XNOR2x1_ASAP7_75t_L g1714 ( 
.A(n_1713),
.B(n_1546),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1714),
.A2(n_1570),
.B1(n_1579),
.B2(n_1568),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1715),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1570),
.B1(n_1565),
.B2(n_1584),
.Y(n_1717)
);

AOI21xp33_ASAP7_75t_L g1718 ( 
.A1(n_1716),
.A2(n_1552),
.B(n_1584),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1717),
.Y(n_1719)
);

OA22x2_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1548),
.B1(n_1545),
.B2(n_1527),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1718),
.A2(n_1406),
.B1(n_1409),
.B2(n_1577),
.Y(n_1721)
);

AOI22x1_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1591),
.B1(n_1548),
.B2(n_1585),
.Y(n_1722)
);

AOI322xp5_ASAP7_75t_L g1723 ( 
.A1(n_1720),
.A2(n_1548),
.A3(n_1577),
.B1(n_1574),
.B2(n_1498),
.C1(n_1591),
.C2(n_1545),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1722),
.A2(n_1574),
.B1(n_1589),
.B2(n_1545),
.Y(n_1724)
);

AOI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1724),
.A2(n_1723),
.B(n_1402),
.C(n_1589),
.Y(n_1725)
);


endmodule