module fake_ariane_1513_n_481 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_481);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_481;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_387;
wire n_406;
wire n_139;
wire n_391;
wire n_349;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_446;
wire n_143;
wire n_152;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_331;
wire n_401;
wire n_267;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_465;
wire n_247;
wire n_240;
wire n_369;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_478;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_390;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_464;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_409;
wire n_171;
wire n_384;
wire n_468;
wire n_182;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_480;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_65),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_31),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_5),
.Y(n_143)
);

INVxp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_7),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_49),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_88),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_46),
.B(n_10),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_47),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_23),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_83),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_119),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_25),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_57),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_108),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_110),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_16),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_41),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_12),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_71),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_34),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_39),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_33),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_4),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_93),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_103),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_94),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_58),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_48),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_50),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_80),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_63),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_86),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_68),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_45),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_35),
.B(n_26),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_8),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_22),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_28),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_121),
.B(n_78),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_53),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g216 ( 
.A(n_152),
.B(n_13),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_0),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_137),
.A2(n_1),
.B(n_3),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_138),
.A2(n_1),
.B(n_4),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_166),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_147),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_139),
.B(n_6),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_141),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_149),
.B(n_14),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_154),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_155),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_167),
.B(n_18),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_197),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_149),
.B(n_19),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_169),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_20),
.Y(n_244)
);

INVxp33_ASAP7_75t_SL g245 ( 
.A(n_158),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_144),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_158),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_170),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_211),
.B1(n_210),
.B2(n_171),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_164),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_168),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_172),
.Y(n_258)
);

OR2x2_ASAP7_75t_SL g259 ( 
.A(n_217),
.B(n_173),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_213),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_229),
.Y(n_263)
);

BUFx4f_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_181),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_213),
.B(n_142),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_174),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_175),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_176),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_148),
.B1(n_190),
.B2(n_206),
.Y(n_273)
);

AND3x4_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_207),
.C(n_198),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_212),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_178),
.Y(n_276)
);

BUFx4_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_214),
.B(n_164),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_180),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_231),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_241),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_240),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_236),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g290 ( 
.A(n_247),
.B(n_226),
.C(n_230),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_230),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_221),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_251),
.A2(n_224),
.B1(n_225),
.B2(n_239),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2x1p5_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_216),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_267),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_228),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_248),
.B(n_228),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_248),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_251),
.A2(n_203),
.B1(n_182),
.B2(n_194),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_221),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_253),
.A2(n_195),
.B1(n_185),
.B2(n_186),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

NAND2x1p5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_150),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_253),
.B(n_219),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_268),
.A2(n_189),
.B(n_193),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_250),
.A2(n_196),
.B(n_201),
.C(n_205),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_254),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

NAND2x1_ASAP7_75t_L g320 ( 
.A(n_253),
.B(n_164),
.Y(n_320)
);

BUFx12f_ASAP7_75t_SL g321 ( 
.A(n_277),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_151),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_242),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_286),
.A2(n_266),
.B1(n_202),
.B2(n_157),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_284),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_292),
.A2(n_312),
.B1(n_301),
.B2(n_305),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_290),
.A2(n_199),
.B1(n_163),
.B2(n_183),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_318),
.A2(n_161),
.B1(n_187),
.B2(n_188),
.Y(n_335)
);

BUFx4f_ASAP7_75t_SL g336 ( 
.A(n_294),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_191),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

NOR3xp33_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_192),
.C(n_262),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_272),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_310),
.A2(n_269),
.B(n_279),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_285),
.B(n_264),
.Y(n_347)
);

AOI222xp33_ASAP7_75t_L g348 ( 
.A1(n_324),
.A2(n_208),
.B1(n_242),
.B2(n_269),
.C1(n_27),
.C2(n_29),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_319),
.B(n_309),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_296),
.A2(n_289),
.B1(n_315),
.B2(n_311),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_208),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_21),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_295),
.A2(n_24),
.B1(n_30),
.B2(n_32),
.Y(n_355)
);

BUFx12f_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_36),
.B(n_37),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_134),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_320),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_317),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_330),
.Y(n_365)
);

AOI32xp33_ASAP7_75t_L g366 ( 
.A1(n_333),
.A2(n_317),
.A3(n_306),
.B1(n_51),
.B2(n_52),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

AO31x2_ASAP7_75t_L g368 ( 
.A1(n_332),
.A2(n_308),
.A3(n_54),
.B(n_55),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_56),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

AO21x2_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_64),
.B(n_67),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_69),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

OAI21x1_ASAP7_75t_L g375 ( 
.A1(n_344),
.A2(n_358),
.B(n_353),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_72),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_348),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_351),
.A2(n_77),
.B(n_82),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_133),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_90),
.Y(n_387)
);

AOI21x1_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_362),
.B(n_335),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

INVx8_ASAP7_75t_L g390 ( 
.A(n_369),
.Y(n_390)
);

AOI222xp33_ASAP7_75t_L g391 ( 
.A1(n_389),
.A2(n_356),
.B1(n_341),
.B2(n_354),
.C1(n_343),
.C2(n_350),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_327),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_327),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_377),
.A2(n_355),
.B1(n_340),
.B2(n_96),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_340),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_385),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_376),
.A2(n_340),
.B(n_355),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_131),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_91),
.B(n_92),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_382),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_97),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_366),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_364),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_400),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

AOI21xp33_ASAP7_75t_L g415 ( 
.A1(n_391),
.A2(n_379),
.B(n_387),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_398),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_405),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_407),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_410),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_387),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_407),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_404),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_366),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_391),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_420),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_421),
.Y(n_429)
);

NAND2x1_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_409),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_408),
.C(n_406),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_393),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

NAND2x1_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_401),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_419),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_390),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_367),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_394),
.B1(n_408),
.B2(n_406),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_413),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_424),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_442),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_441),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_426),
.Y(n_449)
);

NOR3xp33_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_370),
.C(n_402),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_443),
.B(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

OAI21xp33_ASAP7_75t_L g454 ( 
.A1(n_440),
.A2(n_370),
.B(n_401),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_410),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_439),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_446),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_444),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_438),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_429),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_454),
.A2(n_437),
.B1(n_435),
.B2(n_430),
.Y(n_462)
);

AOI32xp33_ASAP7_75t_L g463 ( 
.A1(n_450),
.A2(n_364),
.A3(n_367),
.B1(n_378),
.B2(n_403),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_461),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_459),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_457),
.B(n_456),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_451),
.Y(n_467)
);

OAI221xp5_ASAP7_75t_L g468 ( 
.A1(n_465),
.A2(n_463),
.B1(n_445),
.B2(n_460),
.C(n_462),
.Y(n_468)
);

NOR2x1_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_452),
.Y(n_469)
);

OAI221xp5_ASAP7_75t_L g470 ( 
.A1(n_467),
.A2(n_464),
.B1(n_455),
.B2(n_458),
.C(n_453),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_469),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_470),
.Y(n_472)
);

NAND4xp75_ASAP7_75t_L g473 ( 
.A(n_472),
.B(n_368),
.C(n_372),
.D(n_388),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_471),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_474),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_475),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_476),
.B(n_473),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_R g478 ( 
.A1(n_477),
.A2(n_106),
.B1(n_111),
.B2(n_112),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_478),
.A2(n_114),
.B1(n_117),
.B2(n_120),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_479),
.A2(n_122),
.B1(n_124),
.B2(n_127),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_481)
);


endmodule