module real_jpeg_16297_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_52;
wire n_10;
wire n_9;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_51;
wire n_14;
wire n_47;
wire n_11;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_1),
.B(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

OR2x4_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_22),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_4),
.B(n_12),
.Y(n_11)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_13),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_4),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_4),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_5),
.B(n_14),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_6),
.A2(n_47),
.B1(n_52),
.B2(n_55),
.Y(n_46)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_32),
.B1(n_34),
.B2(n_41),
.C(n_46),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

OAI22xp5_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_10)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_15),
.B(n_19),
.Y(n_13)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_17),
.A2(n_38),
.B(n_40),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

AND2x4_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

OR2x4_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);


endmodule