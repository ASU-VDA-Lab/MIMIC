module fake_jpeg_7933_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_8),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_43),
.B(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_46),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_32),
.B1(n_16),
.B2(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_19),
.B1(n_32),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_68),
.B1(n_22),
.B2(n_18),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_76),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_32),
.B1(n_20),
.B2(n_18),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_70),
.A2(n_16),
.B1(n_29),
.B2(n_30),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_39),
.B1(n_17),
.B2(n_33),
.Y(n_71)
);

AOI22x1_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_81),
.B1(n_17),
.B2(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_79),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_27),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_17),
.B1(n_33),
.B2(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_87),
.Y(n_116)
);

CKINVDCx9p33_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_48),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_95),
.B1(n_101),
.B2(n_115),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_97),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_20),
.B(n_59),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_81),
.B(n_36),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_38),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_102),
.B(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_104),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_110),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_30),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_29),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_36),
.C(n_54),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_120),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_132),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_123),
.B(n_25),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_46),
.B1(n_59),
.B2(n_52),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_144),
.B1(n_118),
.B2(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_133),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_81),
.B1(n_53),
.B2(n_84),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_136),
.B1(n_93),
.B2(n_91),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_81),
.B(n_25),
.C(n_27),
.D(n_31),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_31),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_23),
.Y(n_166)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_142),
.Y(n_179)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_140),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_85),
.B1(n_89),
.B2(n_69),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_17),
.Y(n_138)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_92),
.A2(n_69),
.B1(n_62),
.B2(n_82),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_0),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_147),
.B(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_33),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_64),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_92),
.C(n_100),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_154),
.C(n_173),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_150),
.A2(n_163),
.B1(n_178),
.B2(n_149),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_151),
.B(n_161),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_119),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_155),
.A2(n_157),
.B(n_165),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_169),
.B1(n_174),
.B2(n_177),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_142),
.A2(n_128),
.B1(n_129),
.B2(n_123),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_167),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_162),
.B(n_166),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_91),
.B1(n_104),
.B2(n_105),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_25),
.B(n_24),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_176),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_64),
.B1(n_26),
.B2(n_31),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_5),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_10),
.C(n_15),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_96),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_65),
.C(n_24),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_23),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_181),
.C(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_124),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_9),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_185),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_196),
.Y(n_212)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_201),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_140),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_197),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_146),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_199),
.B(n_203),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_146),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_175),
.C(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

BUFx8_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_10),
.B(n_15),
.C(n_14),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_6),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_7),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_156),
.B1(n_169),
.B2(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_135),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_218),
.C(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_168),
.C(n_165),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_222),
.C(n_224),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_236),
.Y(n_247)
);

AND2x4_ASAP7_75t_SL g222 ( 
.A(n_208),
.B(n_158),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_181),
.C(n_174),
.Y(n_223)
);

NAND2x1p5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_6),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_140),
.B1(n_135),
.B2(n_6),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_228),
.B1(n_200),
.B2(n_190),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_234),
.C(n_192),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_202),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_8),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_9),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_201),
.B1(n_186),
.B2(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_254),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_210),
.C(n_206),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_223),
.C(n_218),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_194),
.B1(n_187),
.B2(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_258),
.C(n_260),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_217),
.C(n_234),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_239),
.B(n_224),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_268),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_224),
.B1(n_226),
.B2(n_231),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_246),
.B1(n_226),
.B2(n_264),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_214),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_270),
.C(n_253),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_216),
.Y(n_275)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_276),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_244),
.B(n_240),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_238),
.B(n_235),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_266),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_261),
.B1(n_267),
.B2(n_259),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_270),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_282),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_281),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_244),
.C(n_237),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_237),
.B1(n_243),
.B2(n_251),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_205),
.B1(n_233),
.B2(n_204),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_243),
.C(n_251),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_182),
.C(n_230),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_283),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_287),
.A2(n_298),
.B(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

INVxp33_ASAP7_75t_SL g301 ( 
.A(n_291),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_SL g293 ( 
.A1(n_285),
.A2(n_228),
.B(n_198),
.C(n_203),
.Y(n_293)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_233),
.B1(n_205),
.B2(n_12),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_280),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_303),
.B(n_293),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_302),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_278),
.B(n_286),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_294),
.C(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_307),
.C(n_292),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_10),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_14),
.C(n_11),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_293),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_313),
.A3(n_301),
.B1(n_306),
.B2(n_305),
.C1(n_14),
.C2(n_11),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_293),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_314),
.A2(n_316),
.B(n_305),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_310),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_315),
.Y(n_319)
);

AOI21x1_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_308),
.B(n_12),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_13),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_13),
.Y(n_323)
);


endmodule