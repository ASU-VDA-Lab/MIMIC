module fake_jpeg_12010_n_202 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_48),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_6),
.A2(n_33),
.B(n_18),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_7),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_39),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_95),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_88),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_0),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_68),
.B1(n_80),
.B2(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_77),
.B1(n_111),
.B2(n_98),
.Y(n_130)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_89),
.Y(n_102)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_76),
.B1(n_80),
.B2(n_68),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_106),
.B1(n_85),
.B2(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_74),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_76),
.B1(n_75),
.B2(n_79),
.Y(n_106)
);

CKINVDCx9p33_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_112),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_117),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_124),
.B1(n_29),
.B2(n_54),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_12),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_96),
.B1(n_79),
.B2(n_70),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_133),
.B1(n_77),
.B2(n_65),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_92),
.C(n_85),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_131),
.C(n_1),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_57),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_126),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_88),
.B1(n_67),
.B2(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_63),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_84),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_58),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_83),
.B(n_67),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_130),
.B(n_134),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_60),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_70),
.B1(n_83),
.B2(n_71),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_132),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_82),
.B1(n_81),
.B2(n_61),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_77),
.B1(n_62),
.B2(n_4),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_117),
.B(n_115),
.C(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_140),
.B1(n_146),
.B2(n_149),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_132),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_10),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_147),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_13),
.B(n_14),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_121),
.B(n_36),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_126),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_155),
.B1(n_35),
.B2(n_40),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_28),
.C(n_30),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_46),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_171),
.B1(n_153),
.B2(n_157),
.C(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_55),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_173),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_41),
.B(n_43),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_159),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_142),
.B1(n_136),
.B2(n_150),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_45),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_175),
.B(n_171),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_137),
.B1(n_148),
.B2(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_183),
.B1(n_168),
.B2(n_174),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_182),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_180),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_160),
.A2(n_166),
.B1(n_162),
.B2(n_174),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_184),
.B(n_183),
.CI(n_181),
.CON(n_187),
.SN(n_187)
);

NOR3xp33_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_184),
.C(n_170),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_191),
.C(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_182),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_161),
.C(n_182),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_190),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_191),
.C(n_188),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_176),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_186),
.A3(n_187),
.B1(n_164),
.B2(n_162),
.C1(n_158),
.C2(n_51),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_200),
.B(n_175),
.C(n_158),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_49),
.Y(n_202)
);


endmodule