module fake_jpeg_26003_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_L g12 ( 
.A1(n_1),
.A2(n_0),
.B(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_6),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_1),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.C(n_24),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_6),
.B1(n_14),
.B2(n_9),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_16),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_18),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_20),
.B1(n_26),
.B2(n_19),
.Y(n_29)
);


endmodule