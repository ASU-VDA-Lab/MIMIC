module fake_netlist_5_2268_n_1680 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1680);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1680;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_12),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVxp33_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_36),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_6),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_108),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_44),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_65),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_83),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_80),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_93),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_67),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_70),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_103),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_47),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_41),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_21),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_43),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_29),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_35),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_66),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_25),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_56),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_73),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_91),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_84),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_28),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_34),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_128),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_104),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_28),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_39),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_54),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_55),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_19),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_19),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_25),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_145),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_31),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_52),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_75),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_43),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_15),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_53),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_120),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_22),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_82),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_16),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_139),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_96),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_125),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_76),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_64),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_4),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_30),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_34),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_59),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_133),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_33),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_129),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_14),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_35),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_20),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_79),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_69),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_151),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_71),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_20),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_68),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_94),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_130),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_50),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_6),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_45),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_10),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_23),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_4),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_41),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_85),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_17),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_131),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_117),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_150),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_11),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_3),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_90),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_15),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_57),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_119),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_49),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_46),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_126),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_89),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_16),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_86),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_113),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_140),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_27),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_87),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_8),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_143),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_78),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_101),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_42),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_42),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_121),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_72),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_8),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_138),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_7),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_63),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_127),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_98),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_37),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_61),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_88),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_58),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_39),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_74),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_7),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_110),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_26),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_199),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_191),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_175),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_175),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_194),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_156),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_178),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_213),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_196),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_161),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_194),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_187),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_178),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_186),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_164),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_278),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_165),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_201),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_197),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_182),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_289),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_198),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_204),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_208),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_225),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_201),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_290),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_234),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_226),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_205),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_226),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_210),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_245),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_246),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_186),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_219),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_202),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_240),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_188),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_246),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_245),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_264),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_264),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_270),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_248),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_254),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_242),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_259),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_199),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_270),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_269),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_273),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_283),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_250),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_298),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_202),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_273),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_222),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_257),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_258),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_250),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_222),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_261),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_275),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_314),
.B(n_275),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_373),
.Y(n_389)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_308),
.A2(n_300),
.B(n_211),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_361),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_311),
.A2(n_256),
.B1(n_281),
.B2(n_252),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_317),
.B(n_280),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_262),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_313),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_322),
.Y(n_405)
);

CKINVDCx8_ASAP7_75t_R g406 ( 
.A(n_344),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_310),
.A2(n_287),
.B1(n_277),
.B2(n_271),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_325),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

NAND2x1p5_ASAP7_75t_L g411 ( 
.A(n_329),
.B(n_280),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_342),
.B(n_262),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_325),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_328),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_351),
.B(n_297),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_333),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_211),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_353),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_300),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_297),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_320),
.A2(n_287),
.B1(n_277),
.B2(n_288),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_381),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_331),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_337),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_338),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_157),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_321),
.B(n_167),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_340),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_363),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_309),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_309),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_324),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_333),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_330),
.A2(n_288),
.B1(n_305),
.B2(n_303),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_158),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_316),
.B(n_252),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_384),
.B(n_159),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_400),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

BUFx4f_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_389),
.B(n_357),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_388),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_398),
.B(n_336),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_L g460 ( 
.A1(n_405),
.A2(n_209),
.B1(n_218),
.B2(n_294),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_412),
.A2(n_307),
.B1(n_297),
.B2(n_368),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_388),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_434),
.Y(n_464)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_417),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_404),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_397),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_385),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_384),
.B(n_345),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_404),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_R g471 ( 
.A(n_448),
.B(n_345),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_404),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_162),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_447),
.B(n_347),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_446),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_451),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_347),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_450),
.B(n_352),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_430),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_419),
.A2(n_334),
.B1(n_163),
.B2(n_173),
.Y(n_484)
);

OAI21xp33_ASAP7_75t_SL g485 ( 
.A1(n_383),
.A2(n_180),
.B(n_171),
.Y(n_485)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_403),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_407),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_352),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_430),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_384),
.B(n_354),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_446),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_184),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_437),
.Y(n_497)
);

AND3x2_ASAP7_75t_L g498 ( 
.A(n_448),
.B(n_244),
.C(n_355),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_385),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_439),
.B(n_354),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_414),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_400),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_396),
.B(n_364),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_411),
.B(n_364),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_385),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_433),
.B(n_378),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_396),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_400),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_429),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_429),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_396),
.B(n_378),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_415),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_411),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_385),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_416),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_411),
.B(n_379),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_400),
.B(n_379),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_444),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_419),
.B(n_192),
.Y(n_529)
);

AND3x2_ASAP7_75t_L g530 ( 
.A(n_419),
.B(n_274),
.C(n_306),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_387),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_395),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_418),
.B(n_323),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_387),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_436),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_408),
.B(n_332),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_400),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_401),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_L g540 ( 
.A1(n_424),
.A2(n_266),
.B1(n_263),
.B2(n_267),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_387),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_438),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_401),
.B(n_155),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_401),
.B(n_402),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_401),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_387),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_419),
.A2(n_216),
.B1(n_220),
.B2(n_302),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_401),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_401),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_402),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_387),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_L g552 ( 
.A(n_417),
.B(n_199),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_387),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_438),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_402),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_441),
.B(n_223),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_406),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_441),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_402),
.B(n_166),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_386),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_402),
.B(n_168),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_402),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_393),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_442),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_393),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_422),
.B(n_231),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_422),
.B(n_255),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_422),
.Y(n_569)
);

BUFx6f_ASAP7_75t_SL g570 ( 
.A(n_422),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_443),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_390),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_395),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_386),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_386),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_394),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_394),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_445),
.B(n_260),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_386),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_420),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_417),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_427),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_391),
.B(n_177),
.Y(n_584)
);

BUFx6f_ASAP7_75t_SL g585 ( 
.A(n_391),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_431),
.B(n_272),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_392),
.B(n_440),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_392),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_431),
.B(n_206),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_440),
.B(n_341),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_390),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_390),
.A2(n_295),
.B1(n_285),
.B2(n_301),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_431),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_427),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_417),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_435),
.B(n_346),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_399),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_399),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_435),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_520),
.B(n_282),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_520),
.B(n_199),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_480),
.B(n_286),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_490),
.B(n_299),
.C(n_170),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_462),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_476),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_462),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_L g607 ( 
.A(n_526),
.B(n_199),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_495),
.Y(n_608)
);

OAI221xp5_ASAP7_75t_L g609 ( 
.A1(n_461),
.A2(n_221),
.B1(n_435),
.B2(n_292),
.C(n_425),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_523),
.B(n_592),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_513),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_573),
.B(n_410),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_513),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_573),
.B(n_591),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_515),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_476),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_591),
.B(n_410),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_454),
.B(n_421),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_455),
.B(n_199),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_494),
.B(n_467),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_516),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_455),
.B(n_199),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_458),
.B(n_169),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_494),
.B(n_475),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_473),
.B(n_406),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_501),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_455),
.B(n_239),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_464),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_569),
.B(n_239),
.Y(n_630)
);

INVx8_ASAP7_75t_L g631 ( 
.A(n_585),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_477),
.B(n_479),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_512),
.A2(n_428),
.B(n_426),
.C(n_425),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_483),
.B(n_421),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_491),
.B(n_426),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_536),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_502),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_488),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_481),
.A2(n_349),
.B1(n_376),
.B2(n_369),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_492),
.B(n_428),
.Y(n_643)
);

A2O1A1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_452),
.A2(n_228),
.B(n_183),
.C(n_189),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_554),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_597),
.A2(n_281),
.B1(n_256),
.B2(n_239),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_504),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_497),
.B(n_160),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_569),
.B(n_239),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_557),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_504),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_511),
.B(n_193),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_597),
.A2(n_239),
.B1(n_190),
.B2(n_188),
.Y(n_653)
);

O2A1O1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_529),
.A2(n_358),
.B(n_367),
.C(n_360),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_558),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_474),
.B(n_169),
.C(n_170),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

INVxp33_ASAP7_75t_L g658 ( 
.A(n_488),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_452),
.B(n_195),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_452),
.B(n_564),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_567),
.B(n_200),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_469),
.B(n_172),
.Y(n_662)
);

NAND2x1_ASAP7_75t_L g663 ( 
.A(n_459),
.B(n_417),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_560),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_510),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_493),
.B(n_239),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_571),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_572),
.B(n_203),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_456),
.B(n_172),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_510),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_518),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_598),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_505),
.B(n_239),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_518),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_517),
.B(n_207),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_543),
.B(n_212),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_559),
.B(n_214),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_598),
.A2(n_188),
.B1(n_190),
.B2(n_167),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_496),
.B(n_215),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_503),
.A2(n_243),
.B(n_217),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_L g681 ( 
.A1(n_456),
.A2(n_359),
.B1(n_284),
.B2(n_279),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_496),
.B(n_224),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_496),
.B(n_561),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_560),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_519),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_589),
.B(n_227),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_519),
.Y(n_687)
);

INVxp33_ASAP7_75t_L g688 ( 
.A(n_533),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_514),
.B(n_249),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_466),
.B(n_247),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_460),
.A2(n_190),
.B1(n_167),
.B2(n_230),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_466),
.B(n_251),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_596),
.B(n_176),
.C(n_174),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_478),
.B(n_174),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_470),
.B(n_253),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_575),
.B(n_265),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_470),
.B(n_472),
.Y(n_697)
);

AND2x4_ASAP7_75t_SL g698 ( 
.A(n_528),
.B(n_230),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_527),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_587),
.A2(n_237),
.B(n_229),
.C(n_304),
.Y(n_700)
);

AND2x2_ASAP7_75t_SL g701 ( 
.A(n_552),
.B(n_230),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_527),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_472),
.B(n_268),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_489),
.B(n_296),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_489),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_507),
.B(n_176),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_481),
.A2(n_233),
.B1(n_179),
.B2(n_284),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_522),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_SL g710 ( 
.A1(n_532),
.A2(n_574),
.B1(n_486),
.B2(n_537),
.Y(n_710)
);

AND2x6_ASAP7_75t_L g711 ( 
.A(n_538),
.B(n_132),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_593),
.B(n_423),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_599),
.B(n_423),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_474),
.B(n_279),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_522),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_500),
.B(n_276),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_544),
.A2(n_538),
.B(n_539),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_539),
.B(n_423),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_548),
.B(n_549),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_548),
.B(n_549),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_473),
.B(n_0),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_555),
.A2(n_423),
.B(n_417),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_588),
.B(n_276),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_525),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_555),
.B(n_423),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_570),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_507),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_556),
.B(n_236),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_581),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_525),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_583),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_562),
.B(n_423),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_562),
.B(n_181),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_485),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_583),
.B(n_144),
.Y(n_735)
);

NAND2x1_ASAP7_75t_L g736 ( 
.A(n_459),
.B(n_142),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_SL g737 ( 
.A(n_465),
.B(n_2),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_594),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_588),
.B(n_141),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_556),
.A2(n_3),
.B1(n_9),
.B2(n_11),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_594),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_471),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_588),
.B(n_135),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_457),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_473),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_584),
.B(n_106),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_508),
.B(n_105),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_465),
.B(n_102),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_577),
.B(n_100),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_577),
.B(n_97),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_577),
.B(n_95),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_457),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_540),
.B(n_13),
.C(n_14),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_453),
.B(n_77),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_453),
.B(n_62),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_570),
.A2(n_51),
.B1(n_48),
.B2(n_21),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_453),
.A2(n_17),
.B(n_18),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_556),
.B(n_18),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_465),
.B(n_22),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_506),
.B(n_23),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_463),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_463),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_529),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_556),
.B(n_24),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_704),
.B(n_487),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_727),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_624),
.B(n_616),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_672),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_706),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_629),
.B(n_563),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_639),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_629),
.B(n_563),
.Y(n_772)
);

INVx5_ASAP7_75t_L g773 ( 
.A(n_711),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_614),
.B(n_565),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_683),
.B(n_565),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_605),
.B(n_699),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_688),
.B(n_486),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_757),
.A2(n_566),
.B(n_568),
.C(n_586),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_631),
.B(n_473),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_741),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_616),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_646),
.A2(n_484),
.B1(n_547),
.B2(n_579),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_707),
.Y(n_783)
);

INVx6_ASAP7_75t_L g784 ( 
.A(n_631),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_615),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_610),
.A2(n_506),
.B(n_545),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_619),
.A2(n_566),
.B(n_568),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_613),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_613),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_621),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_702),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_622),
.Y(n_792)
);

AOI21xp33_ASAP7_75t_L g793 ( 
.A1(n_602),
.A2(n_579),
.B(n_586),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_694),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_701),
.A2(n_579),
.B1(n_585),
.B2(n_578),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_636),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_642),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_645),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_742),
.B(n_557),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_SL g800 ( 
.A1(n_710),
.A2(n_579),
.B1(n_528),
.B2(n_498),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_726),
.B(n_530),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_624),
.B(n_468),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_613),
.B(n_595),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_612),
.B(n_578),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_617),
.B(n_535),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_655),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_664),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_716),
.B(n_535),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_SL g809 ( 
.A(n_681),
.B(n_585),
.C(n_31),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_726),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_752),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_762),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_618),
.B(n_576),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_716),
.B(n_545),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_658),
.B(n_545),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_701),
.A2(n_580),
.B1(n_552),
.B2(n_576),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_618),
.B(n_667),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_650),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_631),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_746),
.B(n_509),
.Y(n_821)
);

CKINVDCx11_ASAP7_75t_R g822 ( 
.A(n_626),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_745),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_604),
.B(n_509),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_626),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_736),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_669),
.B(n_580),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_606),
.B(n_509),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_611),
.B(n_580),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_660),
.B(n_535),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_608),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_620),
.Y(n_832)
);

AND2x6_ASAP7_75t_L g833 ( 
.A(n_657),
.B(n_459),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_657),
.B(n_575),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_714),
.A2(n_482),
.B(n_468),
.C(n_551),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_686),
.B(n_482),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_625),
.B(n_482),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_714),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_684),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_669),
.B(n_575),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_729),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_731),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_633),
.B(n_468),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_632),
.B(n_634),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_L g845 ( 
.A(n_656),
.B(n_760),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_738),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_R g847 ( 
.A(n_684),
.B(n_551),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_635),
.B(n_551),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_761),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_643),
.B(n_506),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_656),
.B(n_595),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_747),
.A2(n_550),
.B1(n_575),
.B2(n_553),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_600),
.B(n_550),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_646),
.B(n_595),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_627),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_637),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_721),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_626),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_676),
.B(n_550),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_728),
.B(n_575),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_711),
.Y(n_861)
);

AND2x6_ASAP7_75t_L g862 ( 
.A(n_758),
.B(n_764),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_747),
.A2(n_499),
.B1(n_553),
.B2(n_546),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_697),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_698),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_693),
.B(n_582),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_673),
.A2(n_499),
.B1(n_553),
.B2(n_546),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_673),
.A2(n_499),
.B1(n_553),
.B2(n_546),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_679),
.B(n_582),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_663),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_638),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_711),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_681),
.B(n_499),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_640),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_647),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_678),
.B(n_29),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_603),
.B(n_499),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_728),
.B(n_521),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_720),
.A2(n_521),
.B(n_553),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_651),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_665),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_670),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_671),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_666),
.B(n_546),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_619),
.A2(n_546),
.B(n_541),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_674),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_641),
.B(n_32),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_659),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_685),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_711),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_721),
.Y(n_891)
);

NOR2x1_ASAP7_75t_L g892 ( 
.A(n_739),
.B(n_541),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_721),
.Y(n_893)
);

BUFx8_ASAP7_75t_L g894 ( 
.A(n_711),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_687),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_709),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_678),
.B(n_32),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_715),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_708),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_719),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_724),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_609),
.A2(n_541),
.B1(n_531),
.B2(n_521),
.Y(n_902)
);

O2A1O1Ixp5_ASAP7_75t_L g903 ( 
.A1(n_666),
.A2(n_541),
.B(n_531),
.C(n_521),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_754),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_682),
.B(n_465),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_623),
.A2(n_541),
.B(n_531),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_730),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_623),
.B(n_531),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_628),
.B(n_531),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_739),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_719),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_753),
.A2(n_521),
.B1(n_534),
.B2(n_582),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_758),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_628),
.B(n_582),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_755),
.B(n_582),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_SL g916 ( 
.A1(n_717),
.A2(n_465),
.B(n_534),
.C(n_37),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_662),
.B(n_534),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_718),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_743),
.B(n_534),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_712),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_675),
.B(n_534),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_743),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_675),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_748),
.B(n_38),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_661),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_668),
.B(n_40),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_601),
.B(n_40),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_601),
.B(n_677),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_764),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_676),
.B(n_677),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_733),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_733),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_648),
.B(n_652),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_630),
.A2(n_649),
.B1(n_703),
.B2(n_705),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_690),
.B(n_695),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_692),
.B(n_689),
.Y(n_936)
);

INVx8_ASAP7_75t_L g937 ( 
.A(n_644),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_713),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_723),
.B(n_654),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_753),
.A2(n_630),
.B1(n_649),
.B2(n_759),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_725),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_732),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_759),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_691),
.B(n_653),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_735),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_607),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_766),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_811),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_786),
.A2(n_750),
.B(n_751),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_785),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_838),
.A2(n_756),
.B1(n_691),
.B2(n_653),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_925),
.B(n_696),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_SL g953 ( 
.A1(n_944),
.A2(n_748),
.B(n_749),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_811),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_853),
.A2(n_722),
.B(n_680),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_767),
.B(n_844),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_913),
.B(n_765),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_790),
.Y(n_958)
);

BUFx12f_ASAP7_75t_L g959 ( 
.A(n_822),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_783),
.B(n_734),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_819),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_850),
.A2(n_700),
.B(n_763),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_792),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_941),
.A2(n_740),
.B(n_737),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_775),
.A2(n_740),
.B(n_936),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_811),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_771),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_831),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_910),
.A2(n_940),
.B1(n_815),
.B2(n_899),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_819),
.B(n_777),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_775),
.A2(n_935),
.B(n_859),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_836),
.A2(n_933),
.B(n_805),
.Y(n_972)
);

CKINVDCx6p67_ASAP7_75t_R g973 ( 
.A(n_779),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_926),
.A2(n_939),
.B(n_845),
.C(n_887),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_862),
.A2(n_782),
.B1(n_943),
.B2(n_931),
.Y(n_975)
);

INVx3_ASAP7_75t_SL g976 ( 
.A(n_858),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_799),
.B(n_832),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_805),
.A2(n_808),
.B(n_908),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_778),
.A2(n_932),
.B(n_928),
.C(n_930),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_832),
.B(n_888),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_908),
.A2(n_909),
.B(n_830),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_888),
.B(n_864),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_788),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_796),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_818),
.B(n_797),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_SL g986 ( 
.A(n_923),
.B(n_922),
.C(n_809),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_782),
.A2(n_876),
.B(n_897),
.C(n_927),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_798),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_781),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_909),
.A2(n_830),
.B(n_821),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_823),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_928),
.A2(n_930),
.B(n_793),
.C(n_787),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_784),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_779),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_806),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_788),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_818),
.B(n_770),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_794),
.B(n_929),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_791),
.B(n_910),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_770),
.B(n_772),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_927),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_779),
.Y(n_1002)
);

BUFx8_ASAP7_75t_L g1003 ( 
.A(n_820),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_784),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_776),
.B(n_816),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_821),
.A2(n_802),
.B(n_914),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_857),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_840),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_878),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_814),
.B(n_891),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_914),
.A2(n_804),
.B(n_787),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_772),
.B(n_862),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_862),
.B(n_827),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_SL g1014 ( 
.A(n_861),
.B(n_872),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_862),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_814),
.B(n_860),
.Y(n_1016)
);

AO32x1_ASAP7_75t_L g1017 ( 
.A1(n_945),
.A2(n_768),
.A3(n_769),
.B1(n_849),
.B2(n_846),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_841),
.B(n_842),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_893),
.B(n_878),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_873),
.A2(n_937),
.B1(n_924),
.B2(n_860),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_800),
.B(n_865),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_937),
.A2(n_924),
.B1(n_854),
.B2(n_829),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_804),
.A2(n_774),
.B(n_906),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_825),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_934),
.A2(n_817),
.B1(n_892),
.B2(n_861),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_774),
.A2(n_885),
.B(n_884),
.Y(n_1026)
);

NOR2x1p5_ASAP7_75t_L g1027 ( 
.A(n_801),
.B(n_789),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_937),
.A2(n_829),
.B1(n_780),
.B2(n_813),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_890),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_773),
.A2(n_872),
.B1(n_795),
.B2(n_890),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_810),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_801),
.B(n_812),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_884),
.A2(n_869),
.B(n_905),
.Y(n_1033)
);

BUFx2_ASAP7_75t_SL g1034 ( 
.A(n_773),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_824),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_871),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_916),
.A2(n_843),
.B(n_835),
.C(n_938),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_807),
.B(n_839),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_855),
.B(n_856),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_918),
.B(n_882),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_911),
.B(n_900),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_894),
.B(n_890),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_918),
.B(n_875),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_773),
.A2(n_843),
.B1(n_902),
.B2(n_863),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_848),
.A2(n_879),
.B(n_919),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_834),
.Y(n_1046)
);

OAI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_912),
.A2(n_877),
.B(n_907),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_874),
.B(n_883),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_919),
.A2(n_915),
.B(n_837),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_903),
.A2(n_828),
.B(n_824),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_942),
.B(n_920),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_881),
.B(n_901),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_886),
.B(n_895),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_SL g1054 ( 
.A(n_894),
.B(n_773),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_904),
.A2(n_852),
.B1(n_898),
.B2(n_946),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_880),
.A2(n_896),
.B(n_889),
.C(n_921),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_834),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_828),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_904),
.A2(n_921),
.B(n_803),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_917),
.A2(n_851),
.B(n_904),
.C(n_866),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_917),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_833),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_898),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_870),
.A2(n_867),
.B(n_868),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_826),
.A2(n_870),
.B1(n_847),
.B2(n_833),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_833),
.B(n_826),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_833),
.Y(n_1067)
);

AND2x2_ASAP7_75t_SL g1068 ( 
.A(n_944),
.B(n_701),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_831),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_786),
.A2(n_455),
.B(n_573),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_811),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_R g1072 ( 
.A(n_925),
.B(n_557),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_767),
.B(n_844),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_785),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_831),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_811),
.B(n_814),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_838),
.A2(n_767),
.B(n_944),
.C(n_704),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_785),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_862),
.A2(n_944),
.B1(n_782),
.B2(n_838),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_785),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_838),
.B(n_704),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_788),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_786),
.A2(n_455),
.B(n_573),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_786),
.A2(n_455),
.B(n_573),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_785),
.Y(n_1085)
);

BUFx4_ASAP7_75t_SL g1086 ( 
.A(n_1004),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_1027),
.B(n_1076),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_956),
.B(n_1073),
.Y(n_1088)
);

AND2x6_ASAP7_75t_L g1089 ( 
.A(n_1062),
.B(n_1029),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1076),
.B(n_1016),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_950),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_958),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_977),
.B(n_997),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_963),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_SL g1095 ( 
.A1(n_974),
.A2(n_1059),
.B(n_987),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1068),
.A2(n_1079),
.B1(n_1000),
.B2(n_969),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_SL g1097 ( 
.A1(n_951),
.A2(n_1025),
.B(n_1044),
.C(n_1055),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_992),
.A2(n_979),
.A3(n_1045),
.B(n_1006),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_978),
.A2(n_1056),
.A3(n_1023),
.B(n_1064),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_971),
.A2(n_972),
.B(n_949),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_982),
.B(n_1001),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1070),
.A2(n_1083),
.B(n_1084),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_947),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_957),
.B(n_980),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_L g1105 ( 
.A(n_948),
.B(n_954),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_990),
.A2(n_1011),
.B(n_955),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1001),
.B(n_1005),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1062),
.Y(n_1108)
);

OA21x2_ASAP7_75t_L g1109 ( 
.A1(n_1050),
.A2(n_1026),
.B(n_962),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_SL g1110 ( 
.A1(n_964),
.A2(n_975),
.B(n_1037),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_965),
.A2(n_1079),
.B(n_1077),
.C(n_953),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1047),
.A2(n_960),
.B(n_964),
.C(n_986),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_989),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1049),
.A2(n_1065),
.B(n_981),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_985),
.B(n_1081),
.Y(n_1115)
);

AOI31xp67_ASAP7_75t_L g1116 ( 
.A1(n_1012),
.A2(n_1013),
.A3(n_1058),
.B(n_1017),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1020),
.A2(n_1008),
.B1(n_1022),
.B2(n_1018),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_970),
.B(n_1032),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1033),
.A2(n_1030),
.B(n_1041),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_993),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_998),
.B(n_989),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1047),
.A2(n_1060),
.B(n_1043),
.C(n_1040),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_984),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_993),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1065),
.A2(n_1014),
.B(n_1066),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_961),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1008),
.B(n_1035),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1072),
.B(n_952),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_999),
.B(n_991),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1021),
.B(n_1007),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_SL g1131 ( 
.A(n_967),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1031),
.B(n_1085),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_959),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1014),
.A2(n_1051),
.B(n_1063),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1010),
.B(n_1016),
.Y(n_1135)
);

CKINVDCx11_ASAP7_75t_R g1136 ( 
.A(n_976),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1038),
.A2(n_1052),
.B(n_1028),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_988),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_SL g1139 ( 
.A1(n_1054),
.A2(n_994),
.B1(n_1002),
.B2(n_1015),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_R g1140 ( 
.A(n_1042),
.B(n_1057),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_SL g1141 ( 
.A1(n_1035),
.A2(n_1080),
.B1(n_1078),
.B2(n_995),
.C(n_1074),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1063),
.A2(n_1053),
.B(n_1048),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_993),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1036),
.B(n_1019),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_948),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1061),
.A2(n_1024),
.B(n_1075),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1009),
.B(n_1046),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1039),
.B(n_1009),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_968),
.A2(n_1069),
.B(n_1067),
.C(n_1054),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1046),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_1003),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1034),
.A2(n_1017),
.B(n_973),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1003),
.Y(n_1153)
);

CKINVDCx11_ASAP7_75t_R g1154 ( 
.A(n_954),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_966),
.B(n_1071),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_R g1156 ( 
.A(n_966),
.B(n_1071),
.Y(n_1156)
);

CKINVDCx8_ASAP7_75t_R g1157 ( 
.A(n_1071),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1029),
.B(n_983),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1082),
.A2(n_971),
.B(n_972),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_996),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_996),
.Y(n_1161)
);

NOR2xp67_ASAP7_75t_SL g1162 ( 
.A(n_1082),
.B(n_727),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_992),
.A2(n_979),
.B(n_971),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_956),
.B(n_1073),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_957),
.B(n_977),
.Y(n_1165)
);

NOR2x1_ASAP7_75t_SL g1166 ( 
.A(n_1034),
.B(n_1063),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_956),
.B(n_1073),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_977),
.B(n_688),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1070),
.A2(n_1084),
.B(n_1083),
.Y(n_1169)
);

CKINVDCx14_ASAP7_75t_R g1170 ( 
.A(n_1072),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_989),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_965),
.B(n_910),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_992),
.A2(n_979),
.B(n_971),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1070),
.A2(n_1084),
.B(n_1083),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_992),
.A2(n_979),
.B(n_971),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_947),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_969),
.A2(n_1073),
.B1(n_956),
.B2(n_1068),
.Y(n_1177)
);

AOI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1011),
.A2(n_978),
.B(n_971),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_950),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_950),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_950),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_961),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_969),
.A2(n_1073),
.B1(n_956),
.B2(n_1068),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_956),
.A2(n_1073),
.B1(n_1068),
.B2(n_1079),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1070),
.A2(n_1084),
.B(n_1083),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_SL g1186 ( 
.A1(n_951),
.A2(n_897),
.B(n_876),
.Y(n_1186)
);

OR2x2_ASAP7_75t_L g1187 ( 
.A(n_970),
.B(n_487),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_965),
.B(n_910),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_956),
.B(n_1073),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_950),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_992),
.A2(n_979),
.B(n_971),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_971),
.A2(n_972),
.B(n_1000),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1044),
.A2(n_1025),
.A3(n_992),
.B(n_979),
.Y(n_1193)
);

INVx3_ASAP7_75t_SL g1194 ( 
.A(n_961),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_992),
.A2(n_979),
.B(n_971),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_950),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_957),
.B(n_977),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_957),
.B(n_977),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_956),
.B(n_1073),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_977),
.B(n_970),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_950),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_SL g1202 ( 
.A1(n_969),
.A2(n_757),
.B(n_747),
.C(n_666),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_998),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_950),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1062),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1070),
.A2(n_1084),
.B(n_1083),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_950),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_992),
.A2(n_979),
.B(n_971),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1070),
.A2(n_1084),
.B(n_1083),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_956),
.B(n_1073),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_L g1211 ( 
.A(n_970),
.B(n_727),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1070),
.A2(n_1084),
.B(n_1083),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1044),
.A2(n_1025),
.A3(n_992),
.B(n_979),
.Y(n_1213)
);

NAND2x1_ASAP7_75t_L g1214 ( 
.A(n_1063),
.B(n_833),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_959),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_956),
.A2(n_1073),
.B1(n_1068),
.B2(n_1079),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_961),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1062),
.Y(n_1218)
);

AO32x2_ASAP7_75t_L g1219 ( 
.A1(n_969),
.A2(n_951),
.A3(n_1044),
.B1(n_1025),
.B2(n_1030),
.Y(n_1219)
);

INVx5_ASAP7_75t_L g1220 ( 
.A(n_948),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1025),
.A2(n_969),
.B(n_1065),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1220),
.B(n_1143),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1088),
.A2(n_1199),
.B1(n_1210),
.B2(n_1164),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1185),
.A2(n_1209),
.B(n_1206),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1176),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1168),
.B(n_1200),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1158),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_SL g1228 ( 
.A(n_1143),
.Y(n_1228)
);

AO32x2_ASAP7_75t_L g1229 ( 
.A1(n_1096),
.A2(n_1184),
.A3(n_1216),
.B1(n_1177),
.B2(n_1183),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1112),
.A2(n_1122),
.B(n_1149),
.C(n_1189),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1182),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1221),
.B(n_1125),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1163),
.A2(n_1175),
.B(n_1173),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1134),
.B(n_1142),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_1096),
.A2(n_1216),
.A3(n_1184),
.B1(n_1117),
.B2(n_1141),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1091),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1092),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1167),
.A2(n_1093),
.B1(n_1115),
.B2(n_1186),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_R g1239 ( 
.A(n_1217),
.B(n_1126),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1123),
.Y(n_1240)
);

AOI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1172),
.A2(n_1188),
.B(n_1119),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1186),
.A2(n_1107),
.B1(n_1203),
.B2(n_1187),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1171),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1138),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_1121),
.B(n_1144),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_1089),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1101),
.B(n_1117),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1127),
.A2(n_1197),
.B1(n_1165),
.B2(n_1198),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1120),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1194),
.A2(n_1130),
.B1(n_1140),
.B2(n_1171),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1118),
.B(n_1104),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1111),
.B(n_1193),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1135),
.B(n_1129),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1179),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1193),
.B(n_1213),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1212),
.A2(n_1102),
.B(n_1114),
.Y(n_1256)
);

OAI222xp33_ASAP7_75t_L g1257 ( 
.A1(n_1139),
.A2(n_1219),
.B1(n_1207),
.B2(n_1196),
.C1(n_1180),
.C2(n_1181),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1113),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1090),
.B(n_1148),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1190),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1106),
.A2(n_1178),
.B(n_1192),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1154),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1201),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1204),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1132),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1128),
.B(n_1170),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1110),
.A2(n_1095),
.B1(n_1211),
.B2(n_1172),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1146),
.B(n_1087),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1163),
.A2(n_1175),
.B(n_1195),
.Y(n_1269)
);

AND2x4_ASAP7_75t_SL g1270 ( 
.A(n_1103),
.B(n_1147),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1157),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1173),
.A2(n_1191),
.B(n_1195),
.C(n_1208),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1147),
.B(n_1150),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1137),
.A2(n_1152),
.B(n_1109),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1086),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1193),
.B(n_1213),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1161),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1116),
.A2(n_1141),
.B(n_1214),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1155),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1108),
.A2(n_1205),
.B(n_1218),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1219),
.A2(n_1089),
.B(n_1213),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1156),
.Y(n_1282)
);

NOR3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1160),
.B(n_1133),
.C(n_1131),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1145),
.B(n_1124),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1219),
.A2(n_1089),
.B(n_1105),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1162),
.A2(n_1220),
.B(n_1145),
.C(n_1098),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1220),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1166),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1153),
.A2(n_1131),
.B1(n_1136),
.B2(n_1215),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1151),
.A2(n_862),
.B1(n_986),
.B2(n_1068),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1099),
.A2(n_1159),
.B(n_1169),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1098),
.A2(n_1159),
.B(n_1169),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1098),
.A2(n_1159),
.B(n_1169),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1182),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1097),
.A2(n_1202),
.B(n_1111),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1088),
.B(n_1164),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1107),
.B(n_1200),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1177),
.A2(n_862),
.B1(n_986),
.B2(n_1068),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1088),
.B(n_1164),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1158),
.Y(n_1300)
);

AOI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1172),
.A2(n_1188),
.B(n_1006),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1159),
.A2(n_1174),
.B(n_1169),
.Y(n_1302)
);

AOI21xp33_ASAP7_75t_L g1303 ( 
.A1(n_1177),
.A2(n_974),
.B(n_987),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1182),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1094),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1136),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1186),
.A2(n_974),
.B(n_939),
.C(n_838),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1159),
.A2(n_1174),
.B(n_1169),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1094),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1177),
.A2(n_862),
.B1(n_986),
.B2(n_1068),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1107),
.B(n_1200),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1186),
.A2(n_974),
.B(n_939),
.C(n_838),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1094),
.Y(n_1313)
);

OR2x6_ASAP7_75t_L g1314 ( 
.A(n_1221),
.B(n_1125),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1102),
.A2(n_1100),
.B(n_1114),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1094),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1094),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1186),
.B(n_716),
.C(n_939),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1094),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1159),
.A2(n_1174),
.B(n_1169),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1159),
.A2(n_1174),
.B(n_1169),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1168),
.B(n_688),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1094),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1220),
.B(n_993),
.Y(n_1324)
);

CKINVDCx11_ASAP7_75t_R g1325 ( 
.A(n_1215),
.Y(n_1325)
);

CKINVDCx8_ASAP7_75t_R g1326 ( 
.A(n_1182),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1088),
.A2(n_1167),
.B1(n_1189),
.B2(n_1164),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1248),
.B(n_1265),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1296),
.A2(n_1299),
.B1(n_1327),
.B2(n_1223),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1223),
.A2(n_1327),
.B1(n_1318),
.B2(n_1297),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1295),
.A2(n_1278),
.B(n_1274),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1259),
.B(n_1251),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1248),
.B(n_1311),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1238),
.B(n_1250),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1318),
.A2(n_1252),
.B1(n_1298),
.B2(n_1310),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_L g1336 ( 
.A1(n_1303),
.A2(n_1295),
.B(n_1307),
.C(n_1312),
.Y(n_1336)
);

AND2x2_ASAP7_75t_SL g1337 ( 
.A(n_1233),
.B(n_1269),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1269),
.A2(n_1238),
.B1(n_1245),
.B2(n_1226),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1286),
.A2(n_1324),
.B(n_1228),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1225),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1290),
.A2(n_1285),
.B1(n_1281),
.B2(n_1243),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1258),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1324),
.A2(n_1228),
.B(n_1285),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1303),
.A2(n_1230),
.B(n_1242),
.C(n_1257),
.Y(n_1344)
);

AOI221x1_ASAP7_75t_SL g1345 ( 
.A1(n_1322),
.A2(n_1253),
.B1(n_1268),
.B2(n_1244),
.C(n_1254),
.Y(n_1345)
);

NOR2x1_ASAP7_75t_SL g1346 ( 
.A(n_1232),
.B(n_1314),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1325),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1255),
.B(n_1276),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1273),
.B(n_1279),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1276),
.B(n_1267),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1243),
.A2(n_1246),
.B1(n_1237),
.B2(n_1260),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1257),
.A2(n_1314),
.B(n_1232),
.C(n_1234),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_SL g1353 ( 
.A1(n_1283),
.A2(n_1239),
.B(n_1246),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1240),
.B(n_1232),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_L g1355 ( 
.A1(n_1278),
.A2(n_1241),
.B(n_1301),
.C(n_1288),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1234),
.A2(n_1264),
.B(n_1263),
.C(n_1316),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1315),
.A2(n_1261),
.B(n_1256),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1309),
.A2(n_1317),
.B1(n_1323),
.B2(n_1313),
.C(n_1319),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1249),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1282),
.A2(n_1305),
.B(n_1284),
.C(n_1266),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1277),
.B(n_1300),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1270),
.B(n_1229),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1229),
.B(n_1287),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1235),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1326),
.A2(n_1289),
.B(n_1222),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1292),
.A2(n_1293),
.B(n_1291),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1271),
.B(n_1280),
.Y(n_1367)
);

OAI211xp5_ASAP7_75t_L g1368 ( 
.A1(n_1275),
.A2(n_1271),
.B(n_1262),
.C(n_1231),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1302),
.A2(n_1308),
.B(n_1321),
.C(n_1320),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_SL g1370 ( 
.A1(n_1271),
.A2(n_1262),
.B(n_1294),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1262),
.B(n_1304),
.Y(n_1371)
);

CKINVDCx6p67_ASAP7_75t_R g1372 ( 
.A(n_1306),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1224),
.B(n_1247),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1272),
.A2(n_939),
.B(n_1318),
.C(n_974),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1236),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1259),
.B(n_1251),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1223),
.B(n_1327),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1247),
.B(n_1238),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1303),
.A2(n_1318),
.B1(n_681),
.B2(n_951),
.C(n_460),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1265),
.B(n_1227),
.Y(n_1380)
);

CKINVDCx14_ASAP7_75t_R g1381 ( 
.A(n_1325),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1259),
.B(n_1251),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1297),
.B(n_970),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1265),
.B(n_1227),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_L g1385 ( 
.A1(n_1303),
.A2(n_1295),
.B(n_1318),
.C(n_1272),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1272),
.A2(n_969),
.B(n_1223),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1259),
.B(n_1251),
.Y(n_1387)
);

OA22x2_ASAP7_75t_L g1388 ( 
.A1(n_1285),
.A2(n_1186),
.B1(n_1238),
.B2(n_395),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1248),
.B(n_1265),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1307),
.A2(n_1312),
.B(n_512),
.C(n_951),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1272),
.A2(n_969),
.B(n_1223),
.Y(n_1391)
);

AOI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1303),
.A2(n_1318),
.B1(n_681),
.B2(n_951),
.C(n_460),
.Y(n_1392)
);

AOI31xp33_ASAP7_75t_L g1393 ( 
.A1(n_1318),
.A2(n_1139),
.A3(n_1290),
.B(n_1298),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1272),
.A2(n_1296),
.B1(n_1299),
.B2(n_1199),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1247),
.B(n_1238),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1322),
.B(n_688),
.Y(n_1396)
);

BUFx2_ASAP7_75t_SL g1397 ( 
.A(n_1228),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1295),
.A2(n_1278),
.B(n_1274),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1249),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1337),
.B(n_1331),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1331),
.B(n_1398),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1373),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1363),
.B(n_1364),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1375),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1379),
.B(n_1392),
.C(n_1390),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1346),
.B(n_1367),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1354),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1329),
.B(n_1377),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1348),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1388),
.B(n_1362),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1366),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1366),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1355),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1388),
.A2(n_1334),
.B1(n_1335),
.B2(n_1330),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1378),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1328),
.B(n_1389),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1378),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1329),
.B(n_1395),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1395),
.B(n_1394),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1350),
.Y(n_1420)
);

OR2x6_ASAP7_75t_L g1421 ( 
.A(n_1352),
.B(n_1386),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1385),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1350),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1369),
.B(n_1357),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1336),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1347),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1356),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1391),
.B(n_1343),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1338),
.B(n_1394),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1374),
.A2(n_1344),
.B(n_1338),
.Y(n_1430)
);

NAND3xp33_ASAP7_75t_L g1431 ( 
.A(n_1330),
.B(n_1393),
.C(n_1360),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1333),
.B(n_1341),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1341),
.B(n_1382),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1351),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1345),
.B(n_1383),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1351),
.A2(n_1335),
.B(n_1361),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1424),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1411),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1411),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1400),
.B(n_1376),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1406),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1431),
.B(n_1342),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1431),
.B(n_1380),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1402),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1402),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1412),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1404),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1400),
.B(n_1387),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1415),
.B(n_1358),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1406),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1401),
.B(n_1332),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1420),
.B(n_1349),
.Y(n_1452)
);

NOR2x1_ASAP7_75t_SL g1453 ( 
.A(n_1428),
.B(n_1397),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1405),
.A2(n_1396),
.B1(n_1381),
.B2(n_1384),
.Y(n_1454)
);

OAI221xp5_ASAP7_75t_L g1455 ( 
.A1(n_1454),
.A2(n_1414),
.B1(n_1405),
.B2(n_1430),
.C(n_1429),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1442),
.A2(n_1429),
.B1(n_1421),
.B2(n_1428),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1454),
.A2(n_1414),
.B1(n_1421),
.B2(n_1419),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1437),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1451),
.B(n_1420),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1442),
.A2(n_1421),
.B1(n_1428),
.B2(n_1419),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1451),
.B(n_1420),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_R g1462 ( 
.A(n_1443),
.B(n_1371),
.Y(n_1462)
);

AOI211xp5_ASAP7_75t_L g1463 ( 
.A1(n_1443),
.A2(n_1422),
.B(n_1435),
.C(n_1408),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1451),
.B(n_1450),
.Y(n_1464)
);

OAI221xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1454),
.A2(n_1421),
.B1(n_1408),
.B2(n_1418),
.C(n_1422),
.Y(n_1465)
);

OAI33xp33_ASAP7_75t_L g1466 ( 
.A1(n_1449),
.A2(n_1435),
.A3(n_1418),
.B1(n_1415),
.B2(n_1417),
.B3(n_1409),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1452),
.A2(n_1421),
.B1(n_1422),
.B2(n_1428),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1438),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1437),
.A2(n_1421),
.B1(n_1428),
.B2(n_1425),
.Y(n_1469)
);

NOR3xp33_ASAP7_75t_L g1470 ( 
.A(n_1449),
.B(n_1425),
.C(n_1427),
.Y(n_1470)
);

AND2x4_ASAP7_75t_SL g1471 ( 
.A(n_1437),
.B(n_1428),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1449),
.A2(n_1421),
.B1(n_1428),
.B2(n_1425),
.C(n_1432),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1444),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1447),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1447),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1452),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1437),
.A2(n_1410),
.B1(n_1434),
.B2(n_1417),
.C(n_1433),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1403),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1437),
.A2(n_1436),
.B1(n_1427),
.B2(n_1407),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1480)
);

NAND3xp33_ASAP7_75t_L g1481 ( 
.A(n_1437),
.B(n_1434),
.C(n_1413),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1444),
.Y(n_1482)
);

AOI222xp33_ASAP7_75t_L g1483 ( 
.A1(n_1453),
.A2(n_1410),
.B1(n_1433),
.B2(n_1426),
.C1(n_1368),
.C2(n_1423),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1440),
.A2(n_1436),
.B1(n_1432),
.B2(n_1410),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1445),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1450),
.B(n_1403),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1452),
.A2(n_1432),
.B1(n_1433),
.B2(n_1416),
.Y(n_1487)
);

INVx5_ASAP7_75t_L g1488 ( 
.A(n_1458),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1484),
.Y(n_1489)
);

INVxp67_ASAP7_75t_SL g1490 ( 
.A(n_1473),
.Y(n_1490)
);

AO21x1_ASAP7_75t_L g1491 ( 
.A1(n_1463),
.A2(n_1470),
.B(n_1457),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1471),
.Y(n_1492)
);

NOR2x1p5_ASAP7_75t_L g1493 ( 
.A(n_1481),
.B(n_1426),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1482),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1485),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1458),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1480),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1458),
.B(n_1441),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1458),
.B(n_1441),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1464),
.B(n_1458),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1466),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1471),
.Y(n_1502)
);

NOR3xp33_ASAP7_75t_L g1503 ( 
.A(n_1455),
.B(n_1399),
.C(n_1413),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1455),
.B(n_1440),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1468),
.A2(n_1446),
.B(n_1439),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1474),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1475),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1480),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1492),
.B(n_1459),
.Y(n_1509)
);

NAND5xp2_ASAP7_75t_L g1510 ( 
.A(n_1503),
.B(n_1465),
.C(n_1483),
.D(n_1463),
.E(n_1456),
.Y(n_1510)
);

OAI21xp33_ASAP7_75t_L g1511 ( 
.A1(n_1501),
.A2(n_1479),
.B(n_1457),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1505),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1505),
.Y(n_1513)
);

AOI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1501),
.A2(n_1465),
.B1(n_1477),
.B2(n_1484),
.C(n_1472),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1492),
.B(n_1459),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1492),
.B(n_1461),
.Y(n_1516)
);

NOR2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1492),
.B(n_1426),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1492),
.B(n_1471),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1506),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1508),
.B(n_1476),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1506),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1502),
.B(n_1461),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1502),
.B(n_1478),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1508),
.B(n_1477),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1494),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1497),
.B(n_1476),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1502),
.B(n_1478),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1491),
.A2(n_1467),
.B1(n_1487),
.B2(n_1460),
.C(n_1469),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1494),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1491),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1488),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1500),
.B(n_1486),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1500),
.B(n_1486),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1502),
.B(n_1441),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1504),
.B(n_1372),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1495),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1504),
.B(n_1445),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1505),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1497),
.B(n_1445),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1491),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1491),
.B(n_1490),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1507),
.Y(n_1544)
);

NOR4xp25_ASAP7_75t_SL g1545 ( 
.A(n_1490),
.B(n_1462),
.C(n_1489),
.D(n_1493),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1511),
.B(n_1503),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1526),
.B(n_1495),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1519),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1519),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1545),
.B(n_1493),
.Y(n_1550)
);

A2O1A1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1531),
.A2(n_1542),
.B(n_1529),
.C(n_1511),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1531),
.B(n_1488),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1521),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1531),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1542),
.B(n_1489),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1514),
.B(n_1440),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1521),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1545),
.B(n_1493),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1526),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1523),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1533),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1514),
.B(n_1440),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1517),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1524),
.B(n_1528),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1448),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1544),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

CKINVDCx16_ASAP7_75t_R g1571 ( 
.A(n_1536),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1533),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1534),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1525),
.B(n_1448),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1530),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1543),
.A2(n_1483),
.B(n_1467),
.Y(n_1576)
);

NAND2x2_ASAP7_75t_L g1577 ( 
.A(n_1517),
.B(n_1359),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1543),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1534),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1525),
.B(n_1448),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1559),
.Y(n_1581)
);

NAND3x1_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1538),
.C(n_1539),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1547),
.B(n_1537),
.Y(n_1584)
);

CKINVDCx16_ASAP7_75t_R g1585 ( 
.A(n_1571),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1510),
.Y(n_1586)
);

CKINVDCx16_ASAP7_75t_R g1587 ( 
.A(n_1571),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1566),
.B(n_1539),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1547),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1566),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1550),
.B(n_1518),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1555),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1565),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1556),
.B(n_1564),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1548),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1574),
.B(n_1580),
.Y(n_1596)
);

CKINVDCx16_ASAP7_75t_R g1597 ( 
.A(n_1565),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1554),
.B(n_1537),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1575),
.B(n_1530),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1549),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1575),
.B(n_1538),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1549),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1553),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1553),
.Y(n_1604)
);

AOI222xp33_ASAP7_75t_L g1605 ( 
.A1(n_1567),
.A2(n_1510),
.B1(n_1541),
.B2(n_1518),
.C1(n_1528),
.C2(n_1516),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1585),
.B(n_1578),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1563),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1584),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1586),
.B(n_1563),
.Y(n_1609)
);

OAI32xp33_ASAP7_75t_L g1610 ( 
.A1(n_1586),
.A2(n_1558),
.A3(n_1550),
.B1(n_1576),
.B2(n_1577),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1605),
.A2(n_1558),
.B1(n_1518),
.B2(n_1577),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1588),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1589),
.B(n_1562),
.Y(n_1613)
);

OAI322xp33_ASAP7_75t_L g1614 ( 
.A1(n_1594),
.A2(n_1561),
.A3(n_1557),
.B1(n_1560),
.B2(n_1570),
.C1(n_1568),
.C2(n_1569),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1591),
.B(n_1597),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1582),
.A2(n_1579),
.B1(n_1573),
.B2(n_1572),
.Y(n_1616)
);

OAI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1592),
.A2(n_1579),
.B1(n_1573),
.B2(n_1572),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1584),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1591),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1590),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1582),
.A2(n_1552),
.B(n_1557),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1581),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1583),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1608),
.B(n_1599),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1620),
.B(n_1593),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1615),
.B(n_1588),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1612),
.B(n_1598),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1608),
.B(n_1601),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1607),
.B(n_1562),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1621),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1609),
.B(n_1596),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1606),
.B(n_1518),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1621),
.B(n_1600),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1627),
.A2(n_1611),
.B1(n_1616),
.B2(n_1617),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1625),
.A2(n_1610),
.B1(n_1622),
.B2(n_1613),
.Y(n_1637)
);

AOI211xp5_ASAP7_75t_SL g1638 ( 
.A1(n_1625),
.A2(n_1623),
.B(n_1614),
.C(n_1619),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1629),
.B(n_1622),
.C(n_1624),
.Y(n_1639)
);

OAI211xp5_ASAP7_75t_L g1640 ( 
.A1(n_1626),
.A2(n_1604),
.B(n_1603),
.C(n_1602),
.Y(n_1640)
);

AOI321xp33_ASAP7_75t_L g1641 ( 
.A1(n_1634),
.A2(n_1631),
.A3(n_1628),
.B1(n_1633),
.B2(n_1630),
.C(n_1632),
.Y(n_1641)
);

AOI221x1_ASAP7_75t_L g1642 ( 
.A1(n_1635),
.A2(n_1570),
.B1(n_1560),
.B2(n_1568),
.C(n_1561),
.Y(n_1642)
);

OAI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1625),
.A2(n_1370),
.B(n_1532),
.C(n_1569),
.Y(n_1643)
);

NOR3x1_ASAP7_75t_L g1644 ( 
.A(n_1626),
.B(n_1532),
.C(n_1541),
.Y(n_1644)
);

NOR3xp33_ASAP7_75t_L g1645 ( 
.A(n_1626),
.B(n_1552),
.C(n_1532),
.Y(n_1645)
);

NAND2xp33_ASAP7_75t_L g1646 ( 
.A(n_1625),
.B(n_1496),
.Y(n_1646)
);

NAND4xp25_ASAP7_75t_L g1647 ( 
.A(n_1641),
.B(n_1552),
.C(n_1340),
.D(n_1535),
.Y(n_1647)
);

OAI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1637),
.A2(n_1527),
.B1(n_1488),
.B2(n_1520),
.C(n_1496),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1636),
.B(n_1639),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1642),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1638),
.A2(n_1552),
.B1(n_1488),
.B2(n_1527),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1646),
.B(n_1488),
.C(n_1496),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1649),
.B(n_1645),
.C(n_1640),
.Y(n_1653)
);

CKINVDCx14_ASAP7_75t_R g1654 ( 
.A(n_1650),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1648),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1651),
.B(n_1644),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1652),
.B(n_1643),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1647),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1653),
.B(n_1509),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1656),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1654),
.B(n_1509),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1655),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1658),
.A2(n_1535),
.B(n_1516),
.Y(n_1663)
);

OAI32xp33_ASAP7_75t_L g1664 ( 
.A1(n_1661),
.A2(n_1657),
.A3(n_1540),
.B1(n_1513),
.B2(n_1512),
.Y(n_1664)
);

NAND2xp33_ASAP7_75t_L g1665 ( 
.A(n_1662),
.B(n_1496),
.Y(n_1665)
);

NOR2x1p5_ASAP7_75t_L g1666 ( 
.A(n_1660),
.B(n_1520),
.Y(n_1666)
);

NOR2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1666),
.B(n_1659),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_L g1668 ( 
.A(n_1667),
.B(n_1665),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1668),
.B(n_1664),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1668),
.A2(n_1663),
.B1(n_1488),
.B2(n_1496),
.Y(n_1670)
);

OR3x2_ASAP7_75t_L g1671 ( 
.A(n_1669),
.B(n_1353),
.C(n_1365),
.Y(n_1671)
);

XNOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1670),
.B(n_1535),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1671),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1672),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1674),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1673),
.B(n_1522),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1513),
.B(n_1512),
.Y(n_1677)
);

XOR2xp5_ASAP7_75t_L g1678 ( 
.A(n_1677),
.B(n_1515),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1496),
.B1(n_1513),
.B2(n_1512),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1339),
.B(n_1496),
.C(n_1540),
.Y(n_1680)
);


endmodule