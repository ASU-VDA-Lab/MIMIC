module real_jpeg_22060_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_20),
.B1(n_21),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_1),
.A2(n_4),
.B1(n_30),
.B2(n_43),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_18),
.B(n_25),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_21),
.B(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_1),
.A2(n_2),
.B1(n_30),
.B2(n_81),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_1),
.A2(n_4),
.B(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_1),
.B(n_92),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_30),
.B(n_36),
.C(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_6),
.B1(n_28),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_4),
.A2(n_6),
.B1(n_28),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_8),
.B1(n_43),
.B2(n_55),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_7),
.A2(n_20),
.B1(n_21),
.B2(n_36),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_7),
.A2(n_35),
.B(n_81),
.C(n_85),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_98),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_96),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_67),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_67),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_52),
.C(n_59),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_14),
.A2(n_15),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_32),
.C(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_23),
.B1(n_26),
.B2(n_29),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_17),
.B(n_29),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_20),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_18),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_19),
.A2(n_21),
.B(n_30),
.C(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_25),
.A2(n_30),
.B(n_55),
.C(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_27),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_30),
.B(n_41),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_30),
.B(n_56),
.Y(n_117)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_34),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_37),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_37),
.B(n_103),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_38),
.B(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B(n_44),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_48),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_43),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_52),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_52),
.B(n_75),
.C(n_125),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_52),
.A2(n_59),
.B1(n_60),
.B2(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_77),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_81),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_74),
.A2(n_75),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_117),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_86),
.B2(n_95),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_94),
.B1(n_107),
.B2(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_107),
.C(n_132),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_135),
.B(n_140),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_129),
.B(n_134),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_120),
.B(n_128),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_112),
.B(n_119),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_111),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_107),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_107),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_110),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B(n_118),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_137),
.Y(n_140)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);


endmodule