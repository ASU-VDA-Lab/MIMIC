module fake_jpeg_2859_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_45),
.Y(n_60)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_33),
.B1(n_14),
.B2(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_58),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_36),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_46),
.C(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_57),
.B1(n_52),
.B2(n_58),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_37),
.B1(n_31),
.B2(n_29),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_70),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_53),
.B(n_51),
.C(n_47),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_44),
.B(n_59),
.C(n_47),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_65),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_81),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_84),
.C(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_59),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_27),
.C(n_32),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_2),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_102),
.C(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_99),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_103),
.B(n_37),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_71),
.C(n_24),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_6),
.B(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_2),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_6),
.C(n_7),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_37),
.B(n_4),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_113),
.B(n_8),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_26),
.C(n_21),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.C(n_115),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_19),
.C(n_17),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_3),
.B(n_4),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_3),
.C(n_5),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_101),
.B1(n_96),
.B2(n_8),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_121),
.B1(n_10),
.B2(n_11),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_107),
.C(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_114),
.B(n_108),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_119),
.B(n_10),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_119),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_127),
.C(n_124),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_9),
.C(n_12),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_13),
.Y(n_132)
);


endmodule