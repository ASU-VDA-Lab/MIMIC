module fake_jpeg_29076_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_4),
.B(n_11),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_63),
.B1(n_55),
.B2(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_51),
.Y(n_85)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_1),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_60),
.C(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_3),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_81),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_3),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_5),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_93),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_78),
.B1(n_65),
.B2(n_66),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_95),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_58),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_14),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_73),
.B(n_72),
.C(n_71),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_104),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_86),
.B1(n_62),
.B2(n_64),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_103),
.B1(n_108),
.B2(n_114),
.Y(n_124)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_86),
.B1(n_92),
.B2(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_65),
.B1(n_68),
.B2(n_54),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_53),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_113),
.C(n_6),
.Y(n_122)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_67),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_68),
.B1(n_61),
.B2(n_59),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_59),
.B1(n_6),
.B2(n_7),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_122),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_8),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_137),
.B(n_18),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_12),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_130),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_12),
.CON(n_129),
.SN(n_129)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_134),
.B(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_13),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_30),
.B(n_44),
.C(n_43),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_40),
.B(n_42),
.C(n_46),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_13),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_135),
.B1(n_126),
.B2(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_15),
.B(n_17),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_121),
.A2(n_115),
.B1(n_15),
.B2(n_21),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_144),
.Y(n_160)
);

AO21x2_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_22),
.B(n_26),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_143),
.B(n_148),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_27),
.B(n_29),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_37),
.B(n_39),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_136),
.C(n_118),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_120),
.C(n_134),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_140),
.Y(n_158)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_156),
.C(n_158),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_140),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_156),
.C(n_154),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_150),
.C(n_160),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_151),
.B(n_163),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_145),
.C(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_168),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_159),
.C(n_152),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_147),
.Y(n_171)
);


endmodule