module fake_jpeg_19309_n_318 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_13),
.Y(n_48)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_51),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_30),
.B1(n_16),
.B2(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_42),
.B1(n_35),
.B2(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_72),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_44),
.B(n_43),
.C(n_40),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_44),
.B(n_61),
.C(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_25),
.B1(n_24),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_35),
.B1(n_37),
.B2(n_51),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_44),
.Y(n_99)
);

NAND2x1p5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_36),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_59),
.B(n_35),
.C(n_29),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_79),
.B1(n_60),
.B2(n_58),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_60),
.B1(n_53),
.B2(n_42),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_49),
.B1(n_51),
.B2(n_62),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_88),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_79),
.B1(n_65),
.B2(n_74),
.Y(n_111)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_46),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_98),
.B(n_65),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_43),
.B1(n_30),
.B2(n_61),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_75),
.B1(n_78),
.B2(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_74),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_75),
.B(n_71),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_108),
.A2(n_18),
.B(n_15),
.Y(n_150)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_110),
.A2(n_111),
.B1(n_119),
.B2(n_124),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_15),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_77),
.B1(n_74),
.B2(n_49),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_93),
.B(n_57),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_122),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_78),
.B1(n_81),
.B2(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_81),
.B1(n_70),
.B2(n_27),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_81),
.B1(n_25),
.B2(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_96),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_82),
.B(n_80),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_89),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_70),
.C(n_31),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_92),
.C(n_94),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_142),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_92),
.B(n_98),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_150),
.B(n_155),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_140),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_85),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_137),
.B(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_147),
.Y(n_166)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_89),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_28),
.B(n_85),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_158),
.B(n_22),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_96),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_157),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_90),
.B(n_70),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_90),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_18),
.B(n_13),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_16),
.A3(n_24),
.B1(n_13),
.B2(n_22),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_124),
.B1(n_119),
.B2(n_121),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_14),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_164),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_19),
.Y(n_162)
);

OR2x4_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_20),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_163),
.A2(n_129),
.B(n_22),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_19),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_130),
.B1(n_115),
.B2(n_112),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_181),
.B1(n_194),
.B2(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_104),
.Y(n_171)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_190),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_111),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_139),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_178),
.B1(n_140),
.B2(n_160),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_112),
.B1(n_130),
.B2(n_113),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_112),
.B1(n_123),
.B2(n_107),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_116),
.B(n_106),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_106),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_81),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_27),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_195),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_149),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_148),
.B1(n_151),
.B2(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_132),
.A2(n_20),
.B1(n_27),
.B2(n_32),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_135),
.A2(n_8),
.B(n_10),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_150),
.C(n_138),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_166),
.B(n_171),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_198),
.A2(n_200),
.B1(n_210),
.B2(n_219),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_131),
.C(n_162),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_201),
.C(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_133),
.B1(n_141),
.B2(n_138),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_156),
.C(n_146),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_207),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_139),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_145),
.C(n_142),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_159),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_169),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_158),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_190),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_166),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_145),
.C(n_31),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_188),
.C(n_181),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_178),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_220),
.A2(n_177),
.B1(n_182),
.B2(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_236),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_202),
.B1(n_195),
.B2(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_167),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_233),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_183),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_170),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_240),
.C(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_241),
.B1(n_213),
.B2(n_219),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_211),
.B1(n_205),
.B2(n_206),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_239),
.Y(n_248)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_180),
.C(n_183),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_172),
.B1(n_168),
.B2(n_180),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_251),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_211),
.B(n_226),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_232),
.B(n_225),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_255),
.Y(n_263)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_210),
.C(n_168),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_184),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_189),
.C(n_170),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_189),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_240),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_179),
.B1(n_194),
.B2(n_32),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_19),
.B(n_8),
.C(n_10),
.D(n_9),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_273),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_223),
.B1(n_235),
.B2(n_227),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_256),
.B1(n_246),
.B2(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_272),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_23),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_31),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_19),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_267),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_264),
.B1(n_268),
.B2(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_276),
.B(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_278),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_256),
.B(n_254),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_279),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_257),
.C(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_286),
.C(n_17),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_248),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_287),
.B1(n_277),
.B2(n_286),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_249),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_9),
.B(n_7),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_9),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_257),
.C(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_29),
.B(n_32),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_293),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_29),
.B(n_17),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_17),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_299),
.A3(n_7),
.B1(n_1),
.B2(n_2),
.C1(n_3),
.C2(n_0),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_0),
.C(n_1),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_284),
.C(n_1),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_9),
.B(n_7),
.Y(n_298)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

AOI211xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_301),
.B(n_304),
.C(n_307),
.Y(n_310)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_303),
.B(n_302),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_290),
.A2(n_0),
.B(n_1),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_0),
.B(n_2),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_311),
.A3(n_295),
.B1(n_296),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_305),
.A2(n_291),
.B(n_295),
.Y(n_309)
);

OAI31xp33_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_310),
.A3(n_300),
.B(n_301),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_313),
.B(n_2),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_294),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_2),
.B(n_3),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_3),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_4),
.B(n_5),
.Y(n_318)
);


endmodule