module fake_jpeg_28059_n_258 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_30),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_23),
.B(n_24),
.C(n_16),
.Y(n_61)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_24),
.B(n_22),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_16),
.B(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_34),
.B1(n_32),
.B2(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_13),
.B1(n_22),
.B2(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_31),
.B1(n_29),
.B2(n_34),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_29),
.B1(n_28),
.B2(n_30),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_30),
.B1(n_26),
.B2(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_82),
.Y(n_105)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_47),
.B1(n_44),
.B2(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_81),
.B1(n_50),
.B2(n_46),
.Y(n_91)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_41),
.C(n_40),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_30),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_40),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_65),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_35),
.B(n_41),
.C(n_32),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_62),
.B(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_35),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_38),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_104),
.B(n_115),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_111),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_59),
.B1(n_50),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_58),
.B1(n_57),
.B2(n_45),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_19),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_108),
.B(n_114),
.Y(n_123)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_97),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_96),
.B(n_100),
.Y(n_134)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_103),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_73),
.C(n_77),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g104 ( 
.A1(n_68),
.A2(n_26),
.B(n_66),
.C(n_45),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_106),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_45),
.A3(n_19),
.B1(n_25),
.B2(n_14),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_14),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_57),
.B1(n_25),
.B2(n_14),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_25),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_82),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_25),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_131),
.Y(n_168)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_78),
.Y(n_127)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_132),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_69),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

OR2x4_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_71),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_143),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx2_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_133),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_73),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_76),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_89),
.A3(n_94),
.B1(n_114),
.B2(n_99),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_114),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_150),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_104),
.C(n_76),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_104),
.B1(n_97),
.B2(n_38),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_122),
.B1(n_126),
.B2(n_137),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_19),
.Y(n_152)
);

NOR4xp25_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_125),
.C(n_121),
.D(n_124),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_38),
.C(n_12),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_156),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_38),
.C(n_12),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_162),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_170),
.B(n_1),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_117),
.A2(n_1),
.B(n_2),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_38),
.C(n_12),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_38),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_175),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_119),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_177),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_119),
.B1(n_126),
.B2(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_168),
.B(n_123),
.CI(n_143),
.CON(n_180),
.SN(n_180)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_120),
.B1(n_134),
.B2(n_142),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_182),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_187),
.B(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_38),
.B1(n_12),
.B2(n_3),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_7),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_159),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_161),
.C(n_147),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_194),
.C(n_207),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_161),
.C(n_169),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_152),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_203),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_155),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_164),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_156),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_174),
.C(n_175),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_201),
.B(n_154),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_192),
.B1(n_178),
.B2(n_172),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_200),
.B1(n_186),
.B2(n_208),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_200),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_176),
.C(n_179),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_195),
.C(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_146),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_197),
.B(n_199),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_165),
.B1(n_166),
.B2(n_148),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_170),
.B1(n_187),
.B2(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_148),
.B1(n_162),
.B2(n_203),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_224),
.A2(n_221),
.B1(n_210),
.B2(n_209),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_210),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_212),
.B(n_217),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_238),
.B(n_2),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_10),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_237),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_209),
.B(n_167),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_167),
.B(n_7),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_239),
.A2(n_222),
.B1(n_224),
.B2(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_7),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_10),
.B(n_9),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_19),
.C(n_12),
.Y(n_246)
);

AOI31xp67_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_236),
.A3(n_19),
.B(n_4),
.Y(n_247)
);

OAI321xp33_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_242),
.B(n_3),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_2),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.C(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_254),
.C(n_4),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_4),
.C(n_5),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_5),
.Y(n_258)
);


endmodule