module fake_jpeg_26296_n_205 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_22),
.B1(n_12),
.B2(n_15),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_39),
.B1(n_12),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_12),
.B1(n_17),
.B2(n_13),
.Y(n_39)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_12),
.B1(n_23),
.B2(n_19),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_47),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_30),
.B(n_19),
.C(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_12),
.B1(n_23),
.B2(n_19),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_51),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_37),
.B1(n_40),
.B2(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_33),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_29),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_29),
.C(n_31),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_31),
.C(n_27),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_32),
.B1(n_21),
.B2(n_17),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_60),
.B1(n_37),
.B2(n_40),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_34),
.B(n_44),
.C(n_27),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_64),
.C(n_67),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_26),
.C(n_33),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_33),
.C(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_77),
.B1(n_50),
.B2(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_75),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_42),
.B1(n_41),
.B2(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_33),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_47),
.C(n_7),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_81),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_53),
.A3(n_58),
.B1(n_60),
.B2(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_24),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_87),
.B(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_89),
.B1(n_62),
.B2(n_63),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_73),
.B1(n_61),
.B2(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_74),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_44),
.C(n_55),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_64),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_91),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_97),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_62),
.C(n_67),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_92),
.C(n_24),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_108),
.B1(n_80),
.B2(n_88),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_76),
.B(n_63),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_85),
.B(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_55),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_111),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_103),
.B1(n_108),
.B2(n_98),
.Y(n_138)
);

NAND2x1_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_79),
.Y(n_111)
);

XOR2x1_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_124),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_16),
.B(n_20),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_92),
.B1(n_85),
.B2(n_16),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_119),
.C(n_122),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_65),
.C(n_54),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_20),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_96),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_65),
.C(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_95),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_136),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_134),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_94),
.B1(n_99),
.B2(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_123),
.B1(n_110),
.B2(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_98),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_142),
.B(n_20),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_140),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_114),
.B1(n_119),
.B2(n_112),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_18),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_120),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_65),
.B(n_20),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_154),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_126),
.B1(n_138),
.B2(n_132),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_147),
.B1(n_150),
.B2(n_20),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_127),
.C(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_20),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_130),
.C(n_136),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_142),
.C(n_21),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_21),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_139),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_158),
.Y(n_169)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_142),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_168),
.C(n_17),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_14),
.B1(n_18),
.B2(n_2),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_8),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_151),
.C(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_167),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_7),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_17),
.C(n_14),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_150),
.B(n_154),
.C(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_175),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_172),
.B(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_157),
.C(n_14),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_14),
.C(n_7),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_11),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_9),
.B(n_8),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_183),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_10),
.C(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_184),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_176),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_8),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_1),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_192),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_177),
.A3(n_169),
.B1(n_170),
.B2(n_9),
.C1(n_4),
.C2(n_0),
.Y(n_189)
);

AOI31xp67_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_1),
.A3(n_2),
.B(n_3),
.Y(n_197)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_197),
.B1(n_189),
.B2(n_3),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_182),
.C(n_2),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_196),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_1),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

AOI321xp33_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_R g203 ( 
.A1(n_201),
.A2(n_199),
.B1(n_5),
.B2(n_6),
.Y(n_203)
);

AOI21x1_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_4),
.B(n_5),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_202),
.Y(n_205)
);


endmodule