module fake_jpeg_25092_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_45),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_46),
.B(n_62),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_55),
.Y(n_104)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_21),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_18),
.B(n_15),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_19),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_15),
.C(n_13),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_39),
.C(n_30),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_12),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_74),
.B(n_11),
.Y(n_116)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_76),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_20),
.B1(n_37),
.B2(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_80),
.A2(n_94),
.B1(n_4),
.B2(n_5),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_41),
.B1(n_26),
.B2(n_24),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_77),
.B1(n_66),
.B2(n_65),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_41),
.B1(n_26),
.B2(n_24),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_98),
.B1(n_102),
.B2(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_90),
.B(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_52),
.B1(n_70),
.B2(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_33),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_0),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_10),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_27),
.B1(n_25),
.B2(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_116),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_23),
.B1(n_22),
.B2(n_40),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_47),
.A2(n_23),
.B(n_39),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_47),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_38),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_127),
.Y(n_190)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_135),
.Y(n_181)
);

INVx5_ASAP7_75t_SL g130 ( 
.A(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_132),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_122),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_10),
.B1(n_38),
.B2(n_2),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_10),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_50),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_136),
.B(n_141),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_82),
.A2(n_60),
.B1(n_73),
.B2(n_68),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_94),
.B1(n_86),
.B2(n_117),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_157),
.B1(n_117),
.B2(n_79),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_95),
.Y(n_141)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx11_ASAP7_75t_SL g191 ( 
.A(n_144),
.Y(n_191)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_80),
.A2(n_76),
.B(n_2),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_146),
.A2(n_152),
.B(n_157),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_81),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_83),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_88),
.A2(n_76),
.B(n_2),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_1),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_153),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_154),
.A2(n_125),
.B1(n_147),
.B2(n_130),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_158),
.Y(n_184)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_86),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_4),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_105),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_111),
.B(n_112),
.C(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_119),
.B1(n_6),
.B2(n_112),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_100),
.B(n_6),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_91),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_167),
.A2(n_170),
.B1(n_172),
.B2(n_180),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_113),
.B1(n_79),
.B2(n_114),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_137),
.B1(n_138),
.B2(n_155),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_91),
.CI(n_97),
.CON(n_173),
.SN(n_173)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_134),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_182),
.B1(n_202),
.B2(n_203),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_114),
.B1(n_99),
.B2(n_120),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_125),
.B1(n_148),
.B2(n_165),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_103),
.B1(n_113),
.B2(n_105),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_97),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_195),
.A2(n_196),
.B(n_200),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_112),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_152),
.B(n_112),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_144),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_137),
.B(n_142),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_205),
.B(n_208),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx13_ASAP7_75t_L g269 ( 
.A(n_206),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_235),
.B1(n_197),
.B2(n_169),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_123),
.Y(n_208)
);

OR2x4_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_142),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_210),
.A2(n_226),
.B(n_197),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_123),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_211),
.B(n_213),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_134),
.C(n_132),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_236),
.C(n_201),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

AO21x2_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_159),
.B(n_128),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_209),
.B(n_207),
.C(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_156),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_225),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_151),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_150),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_147),
.Y(n_230)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_233),
.Y(n_249)
);

BUFx24_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_130),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_129),
.B1(n_145),
.B2(n_143),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_178),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_131),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_239),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_143),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_176),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_172),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_241),
.A2(n_255),
.B(n_263),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_257),
.B1(n_226),
.B2(n_195),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_247),
.B(n_258),
.C(n_272),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_173),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_258),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_206),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_253),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_231),
.A2(n_200),
.B1(n_169),
.B2(n_173),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_201),
.C(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_189),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_233),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_229),
.C(n_226),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_215),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_273),
.B(n_296),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_231),
.B1(n_219),
.B2(n_227),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_280),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_245),
.A2(n_216),
.B1(n_217),
.B2(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_216),
.B1(n_235),
.B2(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_290),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_293),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_241),
.A2(n_195),
.B1(n_196),
.B2(n_187),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_196),
.B1(n_187),
.B2(n_193),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_292),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_212),
.B1(n_176),
.B2(n_205),
.Y(n_286)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_171),
.Y(n_289)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_166),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_294),
.Y(n_311)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_168),
.B(n_204),
.C(n_171),
.D(n_178),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_204),
.B1(n_183),
.B2(n_168),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_266),
.A2(n_263),
.B1(n_265),
.B2(n_256),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_183),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_297),
.B(n_262),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_247),
.C(n_272),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_295),
.C(n_255),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_289),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_309),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_279),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_308),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_253),
.Y(n_310)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_315),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_242),
.C(n_251),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_317),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_263),
.B1(n_266),
.B2(n_243),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_246),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_307),
.B(n_285),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_323),
.B(n_311),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_339),
.C(n_306),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_282),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_314),
.Y(n_347)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_298),
.B(n_292),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_327),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_319),
.A2(n_280),
.B1(n_278),
.B2(n_276),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_331),
.A2(n_333),
.B1(n_335),
.B2(n_340),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_305),
.A2(n_278),
.B1(n_257),
.B2(n_290),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_305),
.A2(n_268),
.B1(n_270),
.B2(n_291),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_299),
.B1(n_243),
.B2(n_320),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_304),
.A2(n_286),
.B1(n_263),
.B2(n_256),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_284),
.C(n_283),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_313),
.Y(n_342)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_299),
.B1(n_312),
.B2(n_320),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_343),
.A2(n_344),
.B1(n_350),
.B2(n_340),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_330),
.B(n_316),
.Y(n_346)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_348),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_306),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_351),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_318),
.B1(n_314),
.B2(n_311),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_354),
.C(n_355),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g356 ( 
.A(n_353),
.B(n_324),
.CI(n_333),
.CON(n_356),
.SN(n_356)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_309),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_259),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_364),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_343),
.A2(n_338),
.B(n_331),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_357),
.A2(n_345),
.B(n_327),
.Y(n_368)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_354),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_362),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_332),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_328),
.C(n_335),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_348),
.C(n_353),
.Y(n_369)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_347),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_365),
.A2(n_267),
.B1(n_269),
.B2(n_179),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_368),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_371),
.C(n_376),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_355),
.C(n_322),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_373),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_259),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_374),
.A2(n_356),
.B1(n_269),
.B2(n_171),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_359),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_357),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_358),
.C(n_360),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_362),
.Y(n_379)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_379),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_382),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_367),
.C(n_366),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_364),
.C(n_356),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_383),
.B(n_370),
.C(n_372),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_385),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_179),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_384),
.B(n_174),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_390),
.A2(n_380),
.B(n_174),
.Y(n_392)
);

A2O1A1O1Ixp25_ASAP7_75t_L g391 ( 
.A1(n_386),
.A2(n_378),
.B(n_379),
.C(n_380),
.D(n_188),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_392),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_393),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_387),
.C(n_388),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_389),
.Y(n_397)
);


endmodule