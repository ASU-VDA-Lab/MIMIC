module real_aes_7264_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_656;
wire n_746;
wire n_532;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_0), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_1), .A2(n_205), .B1(n_313), .B2(n_318), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_2), .Y(n_707) );
XOR2x2_ASAP7_75t_L g427 ( .A(n_3), .B(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_4), .A2(n_174), .B1(n_439), .B2(n_462), .Y(n_542) );
INVx1_ASAP7_75t_L g570 ( .A(n_5), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_6), .A2(n_62), .B1(n_431), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_7), .A2(n_181), .B1(n_498), .B2(n_598), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_8), .Y(n_658) );
INVx1_ASAP7_75t_L g536 ( .A(n_9), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_10), .A2(n_31), .B1(n_219), .B2(n_457), .C1(n_458), .C2(n_461), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_11), .A2(n_115), .B1(n_541), .B2(n_580), .C(n_582), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_12), .A2(n_251), .B1(n_572), .B2(n_822), .Y(n_821) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_13), .A2(n_173), .B1(n_289), .B2(n_443), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_14), .B(n_434), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_15), .A2(n_148), .B1(n_634), .B2(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_16), .A2(n_79), .B1(n_447), .B2(n_449), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_17), .A2(n_28), .B1(n_523), .B2(n_719), .C(n_787), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_18), .A2(n_136), .B1(n_664), .B2(n_665), .C(n_868), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_19), .A2(n_242), .B1(n_528), .B2(n_572), .C(n_575), .Y(n_571) );
INVx1_ASAP7_75t_L g583 ( .A(n_20), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_21), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_22), .A2(n_76), .B1(n_447), .B2(n_565), .C(n_566), .Y(n_564) );
XOR2x2_ASAP7_75t_L g467 ( .A(n_23), .B(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_24), .A2(n_82), .B1(n_523), .B2(n_524), .Y(n_522) );
AOI222xp33_ASAP7_75t_L g585 ( .A1(n_25), .A2(n_35), .B1(n_252), .B2(n_437), .C1(n_457), .C2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g610 ( .A(n_26), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_27), .A2(n_95), .B1(n_461), .B2(n_689), .Y(n_688) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_29), .A2(n_87), .B1(n_294), .B2(n_299), .Y(n_302) );
INVx1_ASAP7_75t_L g811 ( .A(n_29), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_30), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_32), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_33), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_34), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_36), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_37), .A2(n_182), .B1(n_460), .B2(n_612), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_38), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_39), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_40), .A2(n_41), .B1(n_431), .B2(n_434), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_42), .A2(n_55), .B1(n_565), .B2(n_601), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_43), .A2(n_203), .B1(n_325), .B2(n_443), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_44), .Y(n_659) );
AO22x2_ASAP7_75t_L g304 ( .A1(n_45), .A2(n_90), .B1(n_294), .B2(n_295), .Y(n_304) );
INVx1_ASAP7_75t_L g812 ( .A(n_45), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_46), .A2(n_134), .B1(n_552), .B2(n_553), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_47), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_48), .A2(n_51), .B1(n_409), .B2(n_490), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_49), .A2(n_121), .B1(n_392), .B2(n_447), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_50), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_52), .A2(n_152), .B1(n_494), .B2(n_603), .C(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_53), .A2(n_259), .B1(n_458), .B2(n_684), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_54), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_56), .B(n_431), .Y(n_623) );
INVx1_ASAP7_75t_L g531 ( .A(n_57), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_58), .B(n_366), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_59), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_60), .A2(n_236), .B1(n_501), .B2(n_502), .Y(n_500) );
AOI22xp5_ASAP7_75t_SL g595 ( .A1(n_61), .A2(n_256), .B1(n_596), .B2(n_598), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_63), .Y(n_647) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_64), .A2(n_195), .B1(n_694), .B2(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g788 ( .A(n_65), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_66), .Y(n_859) );
XOR2x2_ASAP7_75t_L g677 ( .A(n_67), .B(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_68), .A2(n_207), .B1(n_395), .B2(n_396), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_69), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_70), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_71), .B(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_72), .A2(n_258), .B1(n_359), .B2(n_460), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_73), .A2(n_202), .B1(n_289), .B2(n_395), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_74), .B(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_75), .A2(n_254), .B1(n_475), .B2(n_483), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_77), .Y(n_768) );
INVx1_ASAP7_75t_L g426 ( .A(n_78), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_80), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_81), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_83), .A2(n_161), .B1(n_400), .B2(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_84), .A2(n_157), .B1(n_367), .B2(n_621), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_85), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_86), .A2(n_100), .B1(n_553), .B2(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_88), .A2(n_178), .B1(n_662), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_89), .A2(n_149), .B1(n_395), .B2(n_445), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_91), .A2(n_211), .B1(n_453), .B2(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_92), .A2(n_201), .B1(n_318), .B2(n_603), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_93), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_94), .Y(n_777) );
INVx1_ASAP7_75t_L g278 ( .A(n_96), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_97), .A2(n_128), .B1(n_392), .B2(n_393), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_98), .B(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_99), .A2(n_140), .B1(n_699), .B2(n_722), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_101), .A2(n_815), .B1(n_816), .B2(n_834), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_101), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g633 ( .A1(n_102), .A2(n_183), .B1(n_454), .B2(n_634), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_103), .Y(n_710) );
INVx1_ASAP7_75t_L g276 ( .A(n_104), .Y(n_276) );
INVx1_ASAP7_75t_L g613 ( .A(n_105), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_106), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_107), .A2(n_180), .B1(n_339), .B2(n_498), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_108), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_109), .A2(n_153), .B1(n_400), .B2(n_453), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_110), .A2(n_237), .B1(n_443), .B2(n_445), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_111), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_112), .A2(n_189), .B1(n_487), .B2(n_489), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_113), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_114), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g833 ( .A1(n_116), .A2(n_150), .B1(n_260), .B2(n_359), .C1(n_457), .C2(n_586), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_117), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_118), .A2(n_167), .B1(n_437), .B2(n_460), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_119), .A2(n_133), .B1(n_216), .B2(n_421), .C1(n_671), .C2(n_672), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_120), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_122), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_123), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_124), .A2(n_129), .B1(n_437), .B2(n_438), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_125), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_126), .A2(n_563), .B1(n_587), .B2(n_588), .Y(n_562) );
INVx1_ASAP7_75t_L g587 ( .A(n_126), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_127), .A2(n_206), .B1(n_335), .B2(n_339), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_130), .A2(n_264), .B1(n_453), .B2(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g584 ( .A(n_131), .Y(n_584) );
AO22x2_ASAP7_75t_L g643 ( .A1(n_132), .A2(n_644), .B1(n_673), .B2(n_674), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_132), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_135), .Y(n_778) );
INVx1_ASAP7_75t_L g576 ( .A(n_137), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_138), .A2(n_175), .B1(n_725), .B2(n_726), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_139), .B(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_141), .A2(n_269), .B1(n_664), .B2(n_665), .C(n_666), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_142), .A2(n_250), .B1(n_421), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_143), .A2(n_193), .B1(n_492), .B2(n_494), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_144), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_145), .A2(n_168), .B1(n_598), .B2(n_828), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_146), .Y(n_305) );
INVx1_ASAP7_75t_L g567 ( .A(n_147), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_151), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_154), .Y(n_854) );
INVx2_ASAP7_75t_L g279 ( .A(n_155), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_156), .A2(n_244), .B1(n_367), .B2(n_473), .Y(n_472) );
AO22x1_ASAP7_75t_L g764 ( .A1(n_158), .A2(n_765), .B1(n_793), .B2(n_794), .Y(n_764) );
INVx1_ASAP7_75t_L g793 ( .A(n_158), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_159), .Y(n_770) );
AOI222xp33_ASAP7_75t_L g871 ( .A1(n_160), .A2(n_224), .B1(n_249), .B2(n_672), .C1(n_872), .C2(n_873), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_162), .Y(n_349) );
INVx1_ASAP7_75t_L g578 ( .A(n_163), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_164), .A2(n_218), .B1(n_497), .B2(n_498), .Y(n_496) );
AND2x6_ASAP7_75t_L g275 ( .A(n_165), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_165), .Y(n_805) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_166), .A2(n_230), .B1(n_294), .B2(n_295), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_169), .A2(n_227), .B1(n_479), .B2(n_665), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_170), .Y(n_344) );
INVx1_ASAP7_75t_L g635 ( .A(n_171), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_172), .A2(n_229), .B1(n_308), .B2(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_176), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_177), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_179), .A2(n_238), .B1(n_324), .B2(n_453), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_184), .A2(n_215), .B1(n_719), .B2(n_820), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_185), .A2(n_221), .B1(n_447), .B2(n_548), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_186), .B(n_434), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_187), .B(n_586), .Y(n_775) );
AO22x2_ASAP7_75t_L g298 ( .A1(n_188), .A2(n_246), .B1(n_294), .B2(n_299), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_190), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_191), .A2(n_247), .B1(n_530), .B2(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_192), .B(n_606), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_194), .A2(n_198), .B1(n_395), .B2(n_548), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_196), .A2(n_733), .B1(n_761), .B2(n_762), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_196), .Y(n_761) );
INVx1_ASAP7_75t_L g790 ( .A(n_197), .Y(n_790) );
INVx1_ASAP7_75t_L g519 ( .A(n_199), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_200), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_204), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_208), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_209), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_210), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_212), .Y(n_311) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_213), .A2(n_265), .B1(n_359), .B2(n_439), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_214), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_217), .A2(n_262), .B1(n_574), .B2(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_220), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_222), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_223), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_223), .A2(n_843), .B1(n_845), .B2(n_876), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_225), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_226), .A2(n_241), .B1(n_462), .B2(n_832), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_228), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_230), .B(n_810), .Y(n_809) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_231), .A2(n_271), .B(n_280), .C(n_813), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_232), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_233), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_234), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_235), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_239), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_240), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_243), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_245), .Y(n_782) );
INVx1_ASAP7_75t_L g808 ( .A(n_246), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_248), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_253), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_255), .A2(n_702), .B1(n_728), .B2(n_729), .Y(n_701) );
INVx1_ASAP7_75t_L g728 ( .A(n_255), .Y(n_728) );
INVx1_ASAP7_75t_L g294 ( .A(n_257), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_257), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_261), .B(n_367), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_263), .A2(n_285), .B1(n_383), .B2(n_384), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_263), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_266), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_267), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_268), .B(n_479), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_276), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_277), .A2(n_803), .B(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_640), .B1(n_798), .B2(n_799), .C(n_800), .Y(n_280) );
INVx1_ASAP7_75t_L g798 ( .A(n_281), .Y(n_798) );
AOI22xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_560), .B1(n_561), .B2(n_639), .Y(n_281) );
INVx1_ASAP7_75t_L g639 ( .A(n_282), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_385), .B1(n_558), .B2(n_559), .Y(n_282) );
INVx2_ASAP7_75t_L g558 ( .A(n_283), .Y(n_558) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g384 ( .A(n_285), .Y(n_384) );
AND2x2_ASAP7_75t_SL g285 ( .A(n_286), .B(n_342), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_322), .Y(n_286) );
OAI221xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_305), .B1(n_306), .B2(n_311), .C(n_312), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_289), .Y(n_565) );
BUFx3_ASAP7_75t_L g725 ( .A(n_289), .Y(n_725) );
BUFx3_ASAP7_75t_L g820 ( .A(n_289), .Y(n_820) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_SL g392 ( .A(n_290), .Y(n_392) );
INVx2_ASAP7_75t_L g493 ( .A(n_290), .Y(n_493) );
BUFx2_ASAP7_75t_SL g523 ( .A(n_290), .Y(n_523) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_300), .Y(n_290) );
AND2x6_ASAP7_75t_L g315 ( .A(n_291), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g325 ( .A(n_291), .B(n_326), .Y(n_325) );
AND2x6_ASAP7_75t_L g355 ( .A(n_291), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_297), .Y(n_291) );
AND2x2_ASAP7_75t_L g310 ( .A(n_292), .B(n_298), .Y(n_310) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_293), .B(n_298), .Y(n_321) );
AND2x2_ASAP7_75t_L g331 ( .A(n_293), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g363 ( .A(n_293), .B(n_302), .Y(n_363) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g299 ( .A(n_296), .Y(n_299) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g332 ( .A(n_298), .Y(n_332) );
INVx1_ASAP7_75t_L g362 ( .A(n_298), .Y(n_362) );
AND2x4_ASAP7_75t_L g309 ( .A(n_300), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g319 ( .A(n_300), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_300), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g444 ( .A(n_300), .B(n_331), .Y(n_444) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
OR2x2_ASAP7_75t_L g317 ( .A(n_301), .B(n_304), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_301), .B(n_304), .Y(n_326) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g356 ( .A(n_302), .B(n_304), .Y(n_356) );
AND2x2_ASAP7_75t_L g361 ( .A(n_303), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g375 ( .A(n_303), .Y(n_375) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_306), .A2(n_493), .B1(n_647), .B2(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_309), .Y(n_406) );
INVx2_ASAP7_75t_L g448 ( .A(n_309), .Y(n_448) );
BUFx3_ASAP7_75t_L g501 ( .A(n_309), .Y(n_501) );
BUFx3_ASAP7_75t_L g553 ( .A(n_309), .Y(n_553) );
INVx1_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_310), .B(n_326), .Y(n_352) );
AND2x4_ASAP7_75t_L g433 ( .A(n_310), .B(n_316), .Y(n_433) );
AND2x6_ASAP7_75t_L g435 ( .A(n_310), .B(n_326), .Y(n_435) );
INVx1_ASAP7_75t_L g789 ( .A(n_313), .Y(n_789) );
INVx4_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g393 ( .A(n_314), .Y(n_393) );
INVx4_ASAP7_75t_L g453 ( .A(n_314), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_314), .A2(n_323), .B1(n_655), .B2(n_656), .Y(n_654) );
INVx2_ASAP7_75t_SL g699 ( .A(n_314), .Y(n_699) );
INVx11_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx11_ASAP7_75t_L g488 ( .A(n_315), .Y(n_488) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g347 ( .A(n_317), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_SL g409 ( .A(n_319), .Y(n_409) );
INVx1_ASAP7_75t_L g450 ( .A(n_319), .Y(n_450) );
BUFx3_ASAP7_75t_L g494 ( .A(n_319), .Y(n_494) );
BUFx2_ASAP7_75t_L g530 ( .A(n_319), .Y(n_530) );
BUFx3_ASAP7_75t_L g634 ( .A(n_319), .Y(n_634) );
BUFx3_ASAP7_75t_L g662 ( .A(n_319), .Y(n_662) );
BUFx3_ASAP7_75t_L g822 ( .A(n_319), .Y(n_822) );
AND2x2_ASAP7_75t_L g548 ( .A(n_320), .B(n_375), .Y(n_548) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x6_ASAP7_75t_L g340 ( .A(n_321), .B(n_341), .Y(n_340) );
OAI221xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_327), .B1(n_328), .B2(n_333), .C(n_334), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx6_ASAP7_75t_L g401 ( .A(n_325), .Y(n_401) );
BUFx3_ASAP7_75t_L g454 ( .A(n_325), .Y(n_454) );
BUFx3_ASAP7_75t_L g574 ( .A(n_325), .Y(n_574) );
AND2x2_ASAP7_75t_L g338 ( .A(n_326), .B(n_331), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_326), .B(n_331), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_328), .A2(n_398), .B1(n_399), .B2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g577 ( .A(n_329), .Y(n_577) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g382 ( .A(n_332), .Y(n_382) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g395 ( .A(n_337), .Y(n_395) );
BUFx3_ASAP7_75t_L g499 ( .A(n_337), .Y(n_499) );
INVx4_ASAP7_75t_L g597 ( .A(n_337), .Y(n_597) );
INVx5_ASAP7_75t_L g629 ( .A(n_337), .Y(n_629) );
INVx3_ASAP7_75t_L g828 ( .A(n_337), .Y(n_828) );
INVx8_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g396 ( .A(n_340), .Y(n_396) );
INVx6_ASAP7_75t_SL g445 ( .A(n_340), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_340), .A2(n_567), .B1(n_568), .B2(n_570), .Y(n_566) );
INVx1_ASAP7_75t_L g440 ( .A(n_341), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_353), .C(n_370), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B1(n_349), .B2(n_350), .Y(n_343) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g769 ( .A(n_346), .Y(n_769) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g424 ( .A(n_347), .Y(n_424) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_347), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_350), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_350), .A2(n_424), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g708 ( .A(n_351), .Y(n_708) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g740 ( .A(n_352), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B1(n_358), .B2(n_364), .C(n_365), .Y(n_353) );
OAI21xp5_ASAP7_75t_SL g470 ( .A1(n_354), .A2(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx4_ASAP7_75t_L g416 ( .A(n_355), .Y(n_416) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_355), .Y(n_457) );
BUFx3_ASAP7_75t_L g514 ( .A(n_355), .Y(n_514) );
INVx2_ASAP7_75t_L g618 ( .A(n_355), .Y(n_618) );
INVx1_ASAP7_75t_L g380 ( .A(n_356), .Y(n_380) );
AND2x4_ASAP7_75t_L g462 ( .A(n_356), .B(n_382), .Y(n_462) );
OAI221xp5_ASAP7_75t_SL g709 ( .A1(n_358), .A2(n_609), .B1(n_710), .B2(n_711), .C(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g742 ( .A(n_359), .Y(n_742) );
BUFx4f_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_360), .Y(n_421) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_360), .Y(n_437) );
BUFx2_ASAP7_75t_L g612 ( .A(n_360), .Y(n_612) );
BUFx6f_ASAP7_75t_L g875 ( .A(n_360), .Y(n_875) );
AND2x4_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g369 ( .A(n_362), .Y(n_369) );
AND2x4_ASAP7_75t_L g368 ( .A(n_363), .B(n_369), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_363), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g439 ( .A(n_363), .B(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
BUFx3_ASAP7_75t_L g672 ( .A(n_367), .Y(n_672) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx12f_ASAP7_75t_L g460 ( .A(n_368), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_376), .B2(n_377), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_372), .A2(n_377), .B1(n_748), .B2(n_749), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_372), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx3_ASAP7_75t_SL g413 ( .A(n_373), .Y(n_413) );
INVx4_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g518 ( .A(n_374), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_374), .A2(n_379), .B1(n_869), .B2(n_870), .Y(n_868) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g779 ( .A(n_378), .Y(n_779) );
CKINVDCx16_ASAP7_75t_R g378 ( .A(n_379), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_379), .A2(n_412), .B1(n_413), .B2(n_414), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_379), .A2(n_517), .B1(n_518), .B2(n_519), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_379), .A2(n_518), .B1(n_583), .B2(n_584), .Y(n_582) );
BUFx2_ASAP7_75t_L g669 ( .A(n_379), .Y(n_669) );
OR2x6_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g559 ( .A(n_385), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_463), .B1(n_464), .B2(n_557), .Y(n_385) );
INVx1_ASAP7_75t_L g557 ( .A(n_386), .Y(n_557) );
XOR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_427), .Y(n_386) );
XOR2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_426), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_410), .Y(n_388) );
NOR3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_397), .C(n_403), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g497 ( .A(n_401), .Y(n_497) );
INVx2_ASAP7_75t_L g722 ( .A(n_401), .Y(n_722) );
INVx2_ASAP7_75t_L g792 ( .A(n_401), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_407), .B2(n_408), .Y(n_403) );
INVx4_ASAP7_75t_L g603 ( .A(n_405), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g751 ( .A1(n_405), .A2(n_752), .B1(n_753), .B2(n_754), .C(n_755), .Y(n_751) );
INVx4_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_408), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_575) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_415), .C(n_422), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_413), .A2(n_669), .B1(n_714), .B2(n_715), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B1(n_418), .B2(n_419), .C(n_420), .Y(n_415) );
BUFx2_ASAP7_75t_L g609 ( .A(n_416), .Y(n_609) );
INVx4_ASAP7_75t_L g872 ( .A(n_416), .Y(n_872) );
OAI222xp33_ASAP7_75t_L g741 ( .A1(n_418), .A2(n_742), .B1(n_743), .B2(n_744), .C1(n_745), .C2(n_746), .Y(n_741) );
XOR2x2_ASAP7_75t_L g466 ( .A(n_427), .B(n_467), .Y(n_466) );
NAND4xp75_ASAP7_75t_L g428 ( .A(n_429), .B(n_441), .C(n_451), .D(n_456), .Y(n_428) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_430), .B(n_436), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx5_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
INVx2_ASAP7_75t_L g541 ( .A(n_432), .Y(n_541) );
INVx4_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx4f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
INVx1_ASAP7_75t_SL g581 ( .A(n_435), .Y(n_581) );
BUFx2_ASAP7_75t_L g665 ( .A(n_435), .Y(n_665) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_437), .Y(n_684) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVx1_ASAP7_75t_L g690 ( .A(n_439), .Y(n_690) );
BUFx2_ASAP7_75t_L g832 ( .A(n_439), .Y(n_832) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_446), .Y(n_441) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx3_ASAP7_75t_L g490 ( .A(n_444), .Y(n_490) );
BUFx3_ASAP7_75t_L g524 ( .A(n_444), .Y(n_524) );
BUFx3_ASAP7_75t_L g546 ( .A(n_444), .Y(n_546) );
BUFx2_ASAP7_75t_L g502 ( .A(n_445), .Y(n_502) );
BUFx2_ASAP7_75t_L g598 ( .A(n_445), .Y(n_598) );
BUFx2_ASAP7_75t_L g695 ( .A(n_445), .Y(n_695) );
BUFx4f_ASAP7_75t_SL g785 ( .A(n_445), .Y(n_785) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
INVx2_ASAP7_75t_SL g681 ( .A(n_457), .Y(n_681) );
INVx2_ASAP7_75t_L g744 ( .A(n_457), .Y(n_744) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx4f_ASAP7_75t_SL g586 ( .A(n_460), .Y(n_586) );
BUFx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_462), .Y(n_475) );
BUFx2_ASAP7_75t_SL g621 ( .A(n_462), .Y(n_621) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_503), .B2(n_556), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_484), .Y(n_468) );
NOR2xp33_ASAP7_75t_SL g469 ( .A(n_470), .B(n_476), .Y(n_469) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .C(n_482), .Y(n_476) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_479), .Y(n_664) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_495), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_491), .Y(n_485) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx4_ASAP7_75t_L g528 ( .A(n_488), .Y(n_528) );
INVx2_ASAP7_75t_L g601 ( .A(n_488), .Y(n_601) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_488), .Y(n_826) );
INVx5_ASAP7_75t_SL g864 ( .A(n_488), .Y(n_864) );
BUFx4f_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g760 ( .A(n_490), .Y(n_760) );
INVxp67_ASAP7_75t_L g849 ( .A(n_492), .Y(n_849) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g552 ( .A(n_493), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_500), .Y(n_495) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_501), .Y(n_726) );
INVx1_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
AO22x1_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_532), .B2(n_555), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
XOR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_531), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_520), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .C(n_516), .Y(n_507) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_515), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g535 ( .A1(n_513), .A2(n_536), .B(n_537), .Y(n_535) );
OAI221xp5_ASAP7_75t_L g771 ( .A1(n_513), .A2(n_772), .B1(n_773), .B2(n_774), .C(n_775), .Y(n_771) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_518), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_526), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
INVx1_ASAP7_75t_L g752 ( .A(n_523), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
INVx3_ASAP7_75t_SL g555 ( .A(n_532), .Y(n_555) );
XOR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_554), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_534), .B(n_543), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .C(n_542), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_549), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
INVx1_ASAP7_75t_L g720 ( .A(n_546), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g866 ( .A(n_553), .Y(n_866) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
OA22x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_589), .B1(n_590), .B2(n_638), .Y(n_561) );
INVx1_ASAP7_75t_L g638 ( .A(n_562), .Y(n_638) );
INVx1_ASAP7_75t_L g588 ( .A(n_563), .Y(n_588) );
AND4x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_571), .C(n_579), .D(n_585), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_568), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_568), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_568), .A2(n_652), .B1(n_853), .B2(n_854), .Y(n_852) );
BUFx2_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_577), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_577), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g606 ( .A(n_581), .Y(n_606) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_614), .B1(n_636), .B2(n_637), .Y(n_590) );
INVx2_ASAP7_75t_SL g636 ( .A(n_591), .Y(n_636) );
XOR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_613), .Y(n_591) );
NOR4xp75_ASAP7_75t_L g592 ( .A(n_593), .B(n_599), .C(n_604), .D(n_608), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_595), .Y(n_593) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVxp67_ASAP7_75t_L g652 ( .A(n_598), .Y(n_652) );
NAND2x1_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_605), .B(n_607), .Y(n_604) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g671 ( .A(n_609), .Y(n_671) );
INVx1_ASAP7_75t_L g637 ( .A(n_614), .Y(n_637) );
XOR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_635), .Y(n_614) );
NAND2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_626), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_622), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_619), .B(n_620), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .C(n_625), .Y(n_622) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_629), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx2_ASAP7_75t_L g851 ( .A(n_634), .Y(n_851) );
INVx1_ASAP7_75t_L g799 ( .A(n_640), .Y(n_799) );
AOI22xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_731), .B1(n_796), .B2(n_797), .Y(n_640) );
INVx1_ASAP7_75t_L g796 ( .A(n_641), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_675), .B2(n_676), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g674 ( .A(n_644), .Y(n_674) );
AND4x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_653), .C(n_663), .D(n_670), .Y(n_644) );
NOR2xp33_ASAP7_75t_SL g645 ( .A(n_646), .B(n_649), .Y(n_645) );
NOR2xp33_ASAP7_75t_SL g653 ( .A(n_654), .B(n_657), .Y(n_653) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI22xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_700), .B1(n_701), .B2(n_730), .Y(n_676) );
INVx1_ASAP7_75t_L g730 ( .A(n_677), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_691), .C(n_696), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_685), .Y(n_679) );
OAI21xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B(n_683), .Y(n_680) );
INVx2_ASAP7_75t_SL g773 ( .A(n_684), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .C(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g729 ( .A(n_702), .Y(n_729) );
AND2x2_ASAP7_75t_SL g702 ( .A(n_703), .B(n_716), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_709), .C(n_713), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_706), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_708), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_723), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_721), .Y(n_717) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g858 ( .A(n_722), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
CKINVDCx14_ASAP7_75t_R g797 ( .A(n_731), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_763), .B1(n_764), .B2(n_795), .Y(n_731) );
INVx1_ASAP7_75t_L g795 ( .A(n_732), .Y(n_795) );
INVx1_ASAP7_75t_L g762 ( .A(n_733), .Y(n_762) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_750), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_741), .C(n_747), .Y(n_734) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_756), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g794 ( .A(n_765), .Y(n_794) );
AND3x1_ASAP7_75t_L g765 ( .A(n_766), .B(n_780), .C(n_786), .Y(n_765) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_771), .C(n_776), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_787) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
NOR2x1_ASAP7_75t_L g801 ( .A(n_802), .B(n_806), .Y(n_801) );
OR2x2_ASAP7_75t_SL g879 ( .A(n_802), .B(n_807), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_803), .Y(n_837) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_804), .B(n_839), .Y(n_842) );
CKINVDCx16_ASAP7_75t_R g839 ( .A(n_805), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
OAI322xp33_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_835), .A3(n_838), .B1(n_840), .B2(n_843), .C1(n_844), .C2(n_877), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
NAND4xp75_ASAP7_75t_SL g817 ( .A(n_818), .B(n_823), .C(n_829), .D(n_833), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_821), .Y(n_818) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_827), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND2x2_ASAP7_75t_SL g829 ( .A(n_830), .B(n_831), .Y(n_829) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
CKINVDCx16_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g876 ( .A(n_845), .Y(n_876) );
AND4x1_ASAP7_75t_L g845 ( .A(n_846), .B(n_855), .C(n_867), .D(n_871), .Y(n_845) );
NOR2xp33_ASAP7_75t_SL g846 ( .A(n_847), .B(n_852), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B1(n_850), .B2(n_851), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_862), .B1(n_865), .B2(n_866), .Y(n_860) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx4_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_878), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_879), .Y(n_878) );
endmodule