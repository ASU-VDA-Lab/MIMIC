module fake_ariane_541_n_87 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_87);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_87;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_67;
wire n_34;
wire n_69;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_49;
wire n_20;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_23;
wire n_61;
wire n_22;
wire n_43;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_13),
.B(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_8),
.A2(n_12),
.B1(n_7),
.B2(n_11),
.Y(n_29)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_3),
.B(n_5),
.Y(n_30)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_9),
.A2(n_5),
.B(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_6),
.B1(n_3),
.B2(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_6),
.Y(n_38)
);

NOR2xp67_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_25),
.Y(n_41)
);

AOI221x1_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_25),
.C(n_27),
.Y(n_42)
);

AO31x2_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_26),
.A3(n_29),
.B(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_33),
.B1(n_26),
.B2(n_28),
.Y(n_44)
);

AO31x2_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_26),
.A3(n_29),
.B(n_32),
.Y(n_45)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_21),
.B(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

AOI21x1_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_25),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_23),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

OA21x2_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_21),
.B(n_20),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_43),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_45),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_45),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_47),
.B(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_53),
.B1(n_34),
.B2(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_53),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_47),
.B(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_53),
.B1(n_34),
.B2(n_30),
.Y(n_66)
);

AOI221xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_28),
.B1(n_54),
.B2(n_53),
.C(n_25),
.Y(n_67)
);

OAI221xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_30),
.B1(n_31),
.B2(n_48),
.C(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_55),
.Y(n_70)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_25),
.A3(n_43),
.B1(n_57),
.B2(n_55),
.Y(n_71)
);

OAI321xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_65),
.A3(n_48),
.B1(n_63),
.B2(n_64),
.C(n_57),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_52),
.B(n_30),
.Y(n_73)
);

NAND4xp25_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_43),
.C(n_30),
.D(n_31),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_30),
.B(n_31),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_43),
.C(n_30),
.Y(n_76)
);

AOI222xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_24),
.B1(n_31),
.B2(n_52),
.C1(n_60),
.C2(n_70),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_73),
.B(n_60),
.Y(n_78)
);

AOI211xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_31),
.B(n_24),
.C(n_52),
.Y(n_79)
);

NAND4xp75_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_31),
.C(n_60),
.D(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_75),
.B1(n_79),
.B2(n_74),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_24),
.B1(n_60),
.B2(n_81),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_84),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_80),
.B(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_86),
.Y(n_87)
);


endmodule