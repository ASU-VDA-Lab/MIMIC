module real_aes_8246_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_1), .A2(n_143), .B(n_146), .C(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g209 ( .A(n_2), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_3), .A2(n_138), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_4), .B(n_219), .Y(n_532) );
AOI21xp33_ASAP7_75t_L g220 ( .A1(n_5), .A2(n_138), .B(n_221), .Y(n_220) );
AND2x6_ASAP7_75t_L g143 ( .A(n_6), .B(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_7), .A2(n_189), .B(n_190), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_41), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_9), .A2(n_31), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_9), .Y(n_128) );
INVx1_ASAP7_75t_L g467 ( .A(n_10), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_11), .B(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g226 ( .A(n_12), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_13), .B(n_179), .Y(n_488) );
INVx1_ASAP7_75t_L g164 ( .A(n_14), .Y(n_164) );
INVx1_ASAP7_75t_L g197 ( .A(n_15), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_16), .A2(n_152), .B(n_198), .C(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_17), .B(n_219), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_18), .B(n_154), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_19), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_20), .B(n_568), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_21), .A2(n_178), .B(n_212), .C(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_22), .B(n_219), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_23), .B(n_179), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_24), .A2(n_194), .B(n_196), .C(n_198), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_25), .B(n_179), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_26), .Y(n_517) );
INVx1_ASAP7_75t_L g506 ( .A(n_27), .Y(n_506) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_28), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_29), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_30), .B(n_179), .Y(n_210) );
INVx1_ASAP7_75t_L g127 ( .A(n_31), .Y(n_127) );
INVx1_ASAP7_75t_L g564 ( .A(n_32), .Y(n_564) );
INVx1_ASAP7_75t_L g236 ( .A(n_33), .Y(n_236) );
INVx2_ASAP7_75t_L g141 ( .A(n_34), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_35), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_36), .A2(n_178), .B(n_227), .C(n_530), .Y(n_529) );
INVxp67_ASAP7_75t_L g565 ( .A(n_37), .Y(n_565) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_38), .A2(n_143), .B(n_146), .C(n_149), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_39), .A2(n_146), .B(n_505), .C(n_510), .Y(n_504) );
CKINVDCx14_ASAP7_75t_R g528 ( .A(n_40), .Y(n_528) );
INVx1_ASAP7_75t_L g234 ( .A(n_42), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_43), .A2(n_156), .B(n_224), .C(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_44), .B(n_179), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_45), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_46), .Y(n_561) );
INVx1_ASAP7_75t_L g495 ( .A(n_47), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_48), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_49), .B(n_138), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_50), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_51), .A2(n_146), .B1(n_212), .B2(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_52), .Y(n_166) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_53), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_54), .A2(n_224), .B(n_225), .C(n_227), .Y(n_223) );
CKINVDCx14_ASAP7_75t_R g464 ( .A(n_55), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_56), .Y(n_274) );
INVx1_ASAP7_75t_L g222 ( .A(n_57), .Y(n_222) );
INVx1_ASAP7_75t_L g144 ( .A(n_58), .Y(n_144) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
INVx1_ASAP7_75t_SL g531 ( .A(n_60), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_61), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_62), .B(n_219), .Y(n_499) );
INVx1_ASAP7_75t_L g520 ( .A(n_63), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_SL g244 ( .A1(n_64), .A2(n_154), .B(n_227), .C(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g246 ( .A(n_65), .Y(n_246) );
INVx1_ASAP7_75t_L g107 ( .A(n_66), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_67), .A2(n_138), .B(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_68), .A2(n_102), .B1(n_115), .B2(n_738), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_69), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_70), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_71), .A2(n_138), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g267 ( .A(n_72), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_73), .A2(n_189), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g474 ( .A(n_74), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_75), .Y(n_503) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_76), .A2(n_77), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_76), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_77), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_78), .A2(n_143), .B(n_146), .C(n_269), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_79), .A2(n_138), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g477 ( .A(n_80), .Y(n_477) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_81), .A2(n_126), .B1(n_129), .B2(n_725), .C1(n_726), .C2(n_730), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_82), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g161 ( .A(n_83), .Y(n_161) );
INVx1_ASAP7_75t_L g486 ( .A(n_84), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_85), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_86), .A2(n_143), .B(n_146), .C(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g110 ( .A(n_87), .Y(n_110) );
OR2x2_ASAP7_75t_L g123 ( .A(n_87), .B(n_111), .Y(n_123) );
OR2x2_ASAP7_75t_L g724 ( .A(n_87), .B(n_112), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_88), .A2(n_146), .B(n_519), .C(n_522), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_89), .B(n_172), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_90), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_91), .A2(n_143), .B(n_146), .C(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_92), .Y(n_184) );
INVx1_ASAP7_75t_L g243 ( .A(n_93), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_94), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_95), .B(n_151), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_96), .B(n_168), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_97), .B(n_168), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_98), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_99), .A2(n_138), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g498 ( .A(n_100), .Y(n_498) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx12_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g739 ( .A(n_105), .Y(n_739) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_SL g730 ( .A(n_108), .Y(n_730) );
INVx3_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
NOR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g454 ( .A(n_110), .B(n_112), .Y(n_454) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_125), .B1(n_731), .B2(n_732), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g731 ( .A(n_118), .Y(n_731) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_121), .A2(n_733), .B(n_737), .Y(n_732) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_124), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_123), .Y(n_737) );
INVx1_ASAP7_75t_L g725 ( .A(n_126), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_454), .B1(n_455), .B2(n_724), .Y(n_129) );
INVx2_ASAP7_75t_L g727 ( .A(n_130), .Y(n_727) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_423), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_316), .C(n_389), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_201), .B(n_248), .C(n_300), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
AND2x2_ASAP7_75t_L g264 ( .A(n_135), .B(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g283 ( .A(n_135), .Y(n_283) );
INVx2_ASAP7_75t_L g298 ( .A(n_135), .Y(n_298) );
INVx1_ASAP7_75t_L g328 ( .A(n_135), .Y(n_328) );
AND2x2_ASAP7_75t_L g378 ( .A(n_135), .B(n_299), .Y(n_378) );
AOI32xp33_ASAP7_75t_L g405 ( .A1(n_135), .A2(n_333), .A3(n_406), .B1(n_408), .B2(n_409), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_135), .B(n_254), .Y(n_411) );
AND2x2_ASAP7_75t_L g438 ( .A(n_135), .B(n_281), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_135), .B(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_165), .Y(n_135) );
AOI21xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_145), .B(n_158), .Y(n_136) );
BUFx2_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_139), .B(n_143), .Y(n_206) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g509 ( .A(n_140), .Y(n_509) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g213 ( .A(n_141), .Y(n_213) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx3_ASAP7_75t_L g152 ( .A(n_142), .Y(n_152) );
INVx1_ASAP7_75t_L g154 ( .A(n_142), .Y(n_154) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
INVx4_ASAP7_75t_SL g199 ( .A(n_143), .Y(n_199) );
BUFx3_ASAP7_75t_L g510 ( .A(n_143), .Y(n_510) );
INVx5_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_155), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_151), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_151), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_151), .A2(n_194), .B1(n_564), .B2(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_152), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_152), .B(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_152), .B(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_155), .A2(n_270), .B(n_271), .Y(n_269) );
O2A1O1Ixp5_ASAP7_75t_L g485 ( .A1(n_155), .A2(n_486), .B(n_487), .C(n_488), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_155), .A2(n_487), .B(n_520), .C(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
INVx1_ASAP7_75t_L g272 ( .A(n_158), .Y(n_272) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_204), .B(n_214), .Y(n_203) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_159), .A2(n_231), .B(n_238), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_159), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_161), .B(n_162), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx3_ASAP7_75t_L g219 ( .A(n_167), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_167), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_167), .B(n_512), .Y(n_511) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_167), .A2(n_516), .B(n_523), .Y(n_515) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_168), .A2(n_241), .B(n_247), .Y(n_240) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_168), .Y(n_471) );
AND2x2_ASAP7_75t_L g327 ( .A(n_169), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g349 ( .A(n_169), .Y(n_349) );
AND2x2_ASAP7_75t_L g434 ( .A(n_169), .B(n_264), .Y(n_434) );
AND2x2_ASAP7_75t_L g437 ( .A(n_169), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_186), .Y(n_169) );
INVx2_ASAP7_75t_L g256 ( .A(n_170), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_170), .B(n_281), .Y(n_287) );
AND2x2_ASAP7_75t_L g297 ( .A(n_170), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g333 ( .A(n_170), .Y(n_333) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_183), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_171), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g568 ( .A(n_171), .Y(n_568) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g185 ( .A(n_172), .Y(n_185) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_172), .A2(n_188), .B(n_200), .Y(n_187) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_172), .A2(n_462), .B(n_468), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_172), .A2(n_206), .B(n_503), .C(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_182), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_180), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_178), .B(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g224 ( .A(n_179), .Y(n_224) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx3_ASAP7_75t_L g227 ( .A(n_181), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_185), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_185), .B(n_274), .Y(n_273) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_185), .A2(n_482), .B(n_489), .Y(n_481) );
AND2x2_ASAP7_75t_L g275 ( .A(n_186), .B(n_256), .Y(n_275) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g257 ( .A(n_187), .Y(n_257) );
AND2x2_ASAP7_75t_L g299 ( .A(n_187), .B(n_281), .Y(n_299) );
AND2x2_ASAP7_75t_L g368 ( .A(n_187), .B(n_265), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .C(n_199), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_192), .A2(n_199), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_192), .A2(n_199), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g463 ( .A1(n_192), .A2(n_199), .B(n_464), .C(n_465), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_192), .A2(n_199), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_192), .A2(n_199), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_192), .A2(n_199), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_SL g560 ( .A1(n_192), .A2(n_199), .B(n_561), .C(n_562), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_194), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_194), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_194), .B(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g233 ( .A1(n_195), .A2(n_234), .B1(n_235), .B2(n_236), .Y(n_233) );
INVx2_ASAP7_75t_L g235 ( .A(n_195), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_199), .A2(n_206), .B1(n_232), .B2(n_237), .Y(n_231) );
INVx1_ASAP7_75t_L g522 ( .A(n_199), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_216), .Y(n_201) );
OR2x2_ASAP7_75t_L g262 ( .A(n_202), .B(n_230), .Y(n_262) );
INVx1_ASAP7_75t_L g341 ( .A(n_202), .Y(n_341) );
AND2x2_ASAP7_75t_L g355 ( .A(n_202), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_202), .B(n_229), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_202), .B(n_353), .Y(n_407) );
AND2x2_ASAP7_75t_L g415 ( .A(n_202), .B(n_416), .Y(n_415) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
AND2x2_ASAP7_75t_L g322 ( .A(n_203), .B(n_230), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_206), .A2(n_267), .B(n_268), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_206), .A2(n_483), .B(n_484), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_206), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_216), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g449 ( .A(n_216), .Y(n_449) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_229), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_217), .B(n_293), .Y(n_315) );
OR2x2_ASAP7_75t_L g344 ( .A(n_217), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g376 ( .A(n_217), .B(n_356), .Y(n_376) );
INVx1_ASAP7_75t_SL g396 ( .A(n_217), .Y(n_396) );
AND2x2_ASAP7_75t_L g400 ( .A(n_217), .B(n_261), .Y(n_400) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_218), .B(n_229), .Y(n_253) );
AND2x2_ASAP7_75t_L g260 ( .A(n_218), .B(n_240), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_218), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g303 ( .A(n_218), .B(n_285), .Y(n_303) );
INVx1_ASAP7_75t_SL g310 ( .A(n_218), .Y(n_310) );
BUFx2_ASAP7_75t_L g321 ( .A(n_218), .Y(n_321) );
AND2x2_ASAP7_75t_L g337 ( .A(n_218), .B(n_252), .Y(n_337) );
AND2x2_ASAP7_75t_L g352 ( .A(n_218), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g416 ( .A(n_218), .B(n_230), .Y(n_416) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_228), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_229), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g340 ( .A(n_229), .B(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_229), .A2(n_358), .B1(n_361), .B2(n_364), .C(n_369), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_229), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_240), .Y(n_229) );
INVx3_ASAP7_75t_L g285 ( .A(n_230), .Y(n_285) );
INVx2_ASAP7_75t_L g487 ( .A(n_235), .Y(n_487) );
BUFx2_ASAP7_75t_L g295 ( .A(n_240), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_240), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g326 ( .A(n_240), .Y(n_326) );
OR2x2_ASAP7_75t_L g345 ( .A(n_240), .B(n_285), .Y(n_345) );
INVx3_ASAP7_75t_L g353 ( .A(n_240), .Y(n_353) );
AND2x2_ASAP7_75t_L g356 ( .A(n_240), .B(n_285), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_254), .B1(n_258), .B2(n_263), .C(n_276), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_251), .B(n_325), .Y(n_450) );
OR2x2_ASAP7_75t_L g453 ( .A(n_251), .B(n_284), .Y(n_453) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_252), .A2(n_277), .B1(n_284), .B2(n_286), .C(n_289), .Y(n_276) );
AND2x2_ASAP7_75t_L g293 ( .A(n_252), .B(n_285), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_252), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_252), .B(n_309), .Y(n_308) );
NAND2x1_ASAP7_75t_L g351 ( .A(n_252), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g403 ( .A(n_252), .B(n_345), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_254), .A2(n_363), .B1(n_392), .B2(n_394), .Y(n_391) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI322xp5_ASAP7_75t_L g300 ( .A1(n_255), .A2(n_264), .A3(n_301), .B1(n_304), .B2(n_307), .C1(n_311), .C2(n_314), .Y(n_300) );
OR2x2_ASAP7_75t_L g312 ( .A(n_255), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_256), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g291 ( .A(n_256), .B(n_265), .Y(n_291) );
INVx1_ASAP7_75t_L g306 ( .A(n_256), .Y(n_306) );
AND2x2_ASAP7_75t_L g372 ( .A(n_256), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g282 ( .A(n_257), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g373 ( .A(n_257), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_257), .B(n_281), .Y(n_447) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_261), .B(n_396), .Y(n_395) );
INVx3_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g347 ( .A(n_262), .B(n_294), .Y(n_347) );
OR2x2_ASAP7_75t_L g444 ( .A(n_262), .B(n_295), .Y(n_444) );
INVx1_ASAP7_75t_L g425 ( .A(n_263), .Y(n_425) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_275), .Y(n_263) );
INVx4_ASAP7_75t_L g313 ( .A(n_264), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_264), .B(n_332), .Y(n_338) );
INVx2_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_272), .B(n_273), .Y(n_265) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_272), .A2(n_558), .B(n_566), .Y(n_557) );
INVx1_ASAP7_75t_L g575 ( .A(n_272), .Y(n_575) );
INVx1_ASAP7_75t_L g363 ( .A(n_275), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_275), .B(n_335), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_277), .A2(n_351), .B(n_354), .Y(n_350) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g335 ( .A(n_281), .Y(n_335) );
INVx1_ASAP7_75t_L g362 ( .A(n_281), .Y(n_362) );
INVx1_ASAP7_75t_L g288 ( .A(n_282), .Y(n_288) );
AND2x2_ASAP7_75t_L g290 ( .A(n_282), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g386 ( .A(n_283), .B(n_372), .Y(n_386) );
AND2x2_ASAP7_75t_L g408 ( .A(n_283), .B(n_368), .Y(n_408) );
BUFx2_ASAP7_75t_L g360 ( .A(n_285), .Y(n_360) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AOI32xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_292), .A3(n_293), .B1(n_294), .B2(n_296), .Y(n_289) );
INVx1_ASAP7_75t_L g370 ( .A(n_290), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_290), .A2(n_418), .B1(n_419), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_293), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_293), .B(n_352), .Y(n_393) );
AND2x2_ASAP7_75t_L g440 ( .A(n_293), .B(n_325), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_294), .B(n_341), .Y(n_388) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g441 ( .A(n_296), .Y(n_441) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g366 ( .A(n_297), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_299), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g413 ( .A(n_299), .B(n_333), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_299), .B(n_328), .Y(n_420) );
INVx1_ASAP7_75t_SL g402 ( .A(n_301), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_302), .B(n_353), .Y(n_380) );
NOR4xp25_ASAP7_75t_L g426 ( .A(n_302), .B(n_325), .C(n_427), .D(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_303), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_L g383 ( .A(n_306), .Y(n_383) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_309), .A2(n_400), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g325 ( .A(n_310), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g374 ( .A(n_313), .Y(n_374) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND4xp25_ASAP7_75t_SL g316 ( .A(n_317), .B(n_342), .C(n_357), .D(n_377), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_323), .B(n_327), .C(n_329), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g409 ( .A(n_322), .B(n_352), .Y(n_409) );
AND2x2_ASAP7_75t_L g418 ( .A(n_322), .B(n_396), .Y(n_418) );
INVx3_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_325), .B(n_360), .Y(n_422) );
AND2x2_ASAP7_75t_L g334 ( .A(n_328), .B(n_335), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_336), .B1(n_338), .B2(n_339), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
AND2x2_ASAP7_75t_L g432 ( .A(n_332), .B(n_378), .Y(n_432) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_334), .B(n_383), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_335), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .B(n_348), .C(n_350), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_343), .A2(n_378), .B1(n_379), .B2(n_381), .C(n_384), .Y(n_377) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_351), .A2(n_436), .B1(n_439), .B2(n_441), .C(n_442), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_352), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_360), .B(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_365), .A2(n_385), .B1(n_387), .B2(n_388), .Y(n_384) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B(n_375), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_374), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_385), .A2(n_411), .B1(n_449), .B2(n_450), .C(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
OAI211xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_391), .B(n_397), .C(n_417), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_401), .C(n_410), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_404), .C(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g429 ( .A(n_407), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g451 ( .A1(n_408), .A2(n_434), .B(n_452), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_414), .Y(n_410) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_420), .A2(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_435), .C(n_448), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B(n_431), .C(n_433), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
CKINVDCx14_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g729 ( .A(n_454), .Y(n_729) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_456), .A2(n_724), .B1(n_727), .B2(n_728), .Y(n_726) );
XOR2xp5_ASAP7_75t_L g733 ( .A(n_456), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_654), .Y(n_456) );
NAND5xp2_ASAP7_75t_L g457 ( .A(n_458), .B(n_569), .C(n_601), .D(n_618), .E(n_641), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_500), .B1(n_533), .B2(n_537), .C(n_541), .Y(n_458) );
INVx1_ASAP7_75t_L g681 ( .A(n_459), .Y(n_681) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_479), .Y(n_459) );
AND3x2_ASAP7_75t_L g656 ( .A(n_460), .B(n_481), .C(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_469), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_461), .B(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g548 ( .A(n_461), .Y(n_548) );
AND2x2_ASAP7_75t_L g552 ( .A(n_461), .B(n_491), .Y(n_552) );
INVx2_ASAP7_75t_L g578 ( .A(n_461), .Y(n_578) );
OR2x2_ASAP7_75t_L g589 ( .A(n_461), .B(n_492), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_461), .B(n_480), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_461), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g668 ( .A(n_461), .B(n_492), .Y(n_668) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_469), .Y(n_551) );
AND2x2_ASAP7_75t_L g609 ( .A(n_469), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_469), .B(n_480), .Y(n_628) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g540 ( .A(n_470), .B(n_480), .Y(n_540) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_470), .Y(n_547) );
AND2x2_ASAP7_75t_L g595 ( .A(n_470), .B(n_492), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_470), .B(n_479), .C(n_578), .Y(n_620) );
AND2x2_ASAP7_75t_L g685 ( .A(n_470), .B(n_481), .Y(n_685) );
AND2x2_ASAP7_75t_L g719 ( .A(n_470), .B(n_480), .Y(n_719) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_478), .Y(n_470) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_471), .A2(n_493), .B(n_499), .Y(n_492) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_471), .A2(n_526), .B(n_532), .Y(n_525) );
INVxp67_ASAP7_75t_L g549 ( .A(n_479), .Y(n_549) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_491), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_480), .B(n_578), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_480), .B(n_609), .Y(n_617) );
AND2x2_ASAP7_75t_L g667 ( .A(n_480), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g695 ( .A(n_480), .Y(n_695) );
INVx4_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g602 ( .A(n_481), .B(n_595), .Y(n_602) );
BUFx3_ASAP7_75t_L g634 ( .A(n_481), .Y(n_634) );
INVx2_ASAP7_75t_L g610 ( .A(n_491), .Y(n_610) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_492), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_500), .A2(n_670), .B1(n_672), .B2(n_673), .Y(n_669) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_513), .Y(n_500) );
AND2x2_ASAP7_75t_L g533 ( .A(n_501), .B(n_534), .Y(n_533) );
INVx3_ASAP7_75t_SL g544 ( .A(n_501), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_501), .B(n_573), .Y(n_605) );
OR2x2_ASAP7_75t_L g624 ( .A(n_501), .B(n_514), .Y(n_624) );
AND2x2_ASAP7_75t_L g629 ( .A(n_501), .B(n_581), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_501), .B(n_574), .Y(n_632) );
AND2x2_ASAP7_75t_L g644 ( .A(n_501), .B(n_525), .Y(n_644) );
AND2x2_ASAP7_75t_L g660 ( .A(n_501), .B(n_515), .Y(n_660) );
AND2x4_ASAP7_75t_L g663 ( .A(n_501), .B(n_535), .Y(n_663) );
OR2x2_ASAP7_75t_L g680 ( .A(n_501), .B(n_616), .Y(n_680) );
OR2x2_ASAP7_75t_L g711 ( .A(n_501), .B(n_557), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_501), .B(n_639), .Y(n_713) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_509), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g587 ( .A(n_513), .B(n_555), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_513), .B(n_574), .Y(n_706) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_525), .Y(n_513) );
AND2x2_ASAP7_75t_L g543 ( .A(n_514), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g573 ( .A(n_514), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g581 ( .A(n_514), .B(n_557), .Y(n_581) );
AND2x2_ASAP7_75t_L g599 ( .A(n_514), .B(n_535), .Y(n_599) );
OR2x2_ASAP7_75t_L g616 ( .A(n_514), .B(n_574), .Y(n_616) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g536 ( .A(n_515), .Y(n_536) );
AND2x2_ASAP7_75t_L g639 ( .A(n_515), .B(n_525), .Y(n_639) );
INVx2_ASAP7_75t_L g535 ( .A(n_525), .Y(n_535) );
INVx1_ASAP7_75t_L g651 ( .A(n_525), .Y(n_651) );
AND2x2_ASAP7_75t_L g701 ( .A(n_525), .B(n_544), .Y(n_701) );
AND2x2_ASAP7_75t_L g554 ( .A(n_534), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g585 ( .A(n_534), .B(n_544), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_534), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g572 ( .A(n_535), .B(n_544), .Y(n_572) );
OR2x2_ASAP7_75t_L g688 ( .A(n_536), .B(n_662), .Y(n_688) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_539), .B(n_668), .Y(n_674) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
OAI32xp33_ASAP7_75t_L g630 ( .A1(n_540), .A2(n_631), .A3(n_633), .B1(n_635), .B2(n_636), .Y(n_630) );
OR2x2_ASAP7_75t_L g647 ( .A(n_540), .B(n_589), .Y(n_647) );
OAI21xp33_ASAP7_75t_SL g672 ( .A1(n_540), .A2(n_550), .B(n_577), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .B1(n_550), .B2(n_553), .Y(n_541) );
INVxp33_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_543), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_544), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g598 ( .A(n_544), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g698 ( .A(n_544), .B(n_639), .Y(n_698) );
OR2x2_ASAP7_75t_L g722 ( .A(n_544), .B(n_616), .Y(n_722) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_545), .A2(n_604), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g582 ( .A(n_547), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_547), .B(n_552), .Y(n_600) );
AND2x2_ASAP7_75t_L g622 ( .A(n_548), .B(n_595), .Y(n_622) );
INVx1_ASAP7_75t_L g635 ( .A(n_548), .Y(n_635) );
OR2x2_ASAP7_75t_L g640 ( .A(n_548), .B(n_574), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_551), .B(n_589), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_552), .A2(n_571), .B1(n_576), .B2(n_580), .Y(n_570) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_555), .A2(n_613), .B1(n_620), .B2(n_621), .Y(n_619) );
AND2x2_ASAP7_75t_L g697 ( .A(n_555), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_557), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g716 ( .A(n_557), .B(n_599), .Y(n_716) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_559), .A2(n_567), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_582), .B1(n_583), .B2(n_588), .C(n_590), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_572), .B(n_574), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_572), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g591 ( .A(n_573), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_573), .A2(n_679), .B(n_680), .C(n_681), .Y(n_678) );
AND2x2_ASAP7_75t_L g683 ( .A(n_573), .B(n_663), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_SL g721 ( .A1(n_573), .A2(n_662), .B(n_722), .C(n_723), .Y(n_721) );
BUFx3_ASAP7_75t_L g613 ( .A(n_574), .Y(n_613) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_577), .B(n_634), .Y(n_677) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_577), .A2(n_697), .B(n_699), .C(n_705), .Y(n_696) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVxp67_ASAP7_75t_L g657 ( .A(n_579), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_581), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_585), .A2(n_602), .B(n_603), .C(n_611), .Y(n_601) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g686 ( .A(n_589), .Y(n_686) );
OR2x2_ASAP7_75t_L g703 ( .A(n_589), .B(n_633), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_597), .B2(n_600), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_592), .A2(n_604), .B1(n_605), .B2(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
OR2x2_ASAP7_75t_L g690 ( .A(n_594), .B(n_634), .Y(n_690) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g645 ( .A(n_595), .B(n_635), .Y(n_645) );
INVx1_ASAP7_75t_L g653 ( .A(n_596), .Y(n_653) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_599), .B(n_613), .Y(n_661) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_609), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g718 ( .A(n_610), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g648 ( .A(n_612), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_613), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_613), .B(n_644), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g664 ( .A(n_613), .B(n_639), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_613), .B(n_660), .Y(n_671) );
OAI211xp5_ASAP7_75t_L g675 ( .A1(n_613), .A2(n_623), .B(n_663), .C(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AOI221xp5_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_623), .B1(n_625), .B2(n_629), .C(n_630), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_627), .B(n_635), .Y(n_709) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_629), .A2(n_644), .B(n_646), .C(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_632), .B(n_639), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_633), .B(n_686), .Y(n_723) );
CKINVDCx16_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
INVxp33_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
AOI21xp33_ASAP7_75t_SL g649 ( .A1(n_638), .A2(n_650), .B(n_652), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_638), .B(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_639), .B(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_645), .B1(n_646), .B2(n_648), .C(n_649), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_645), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g679 ( .A(n_651), .Y(n_679) );
NAND5xp2_ASAP7_75t_L g654 ( .A(n_655), .B(n_682), .C(n_696), .D(n_707), .E(n_720), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B(n_665), .C(n_678), .Y(n_655) );
INVx2_ASAP7_75t_SL g702 ( .A(n_656), .Y(n_702) );
NAND4xp25_ASAP7_75t_SL g658 ( .A(n_659), .B(n_661), .C(n_662), .D(n_664), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g665 ( .A1(n_664), .A2(n_666), .B(n_669), .C(n_675), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_667), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_667), .A2(n_708), .B1(n_710), .B2(n_712), .C(n_714), .Y(n_707) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_684), .B1(n_687), .B2(n_689), .C(n_691), .Y(n_682) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_690), .A2(n_713), .B1(n_715), .B2(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_699) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
endmodule