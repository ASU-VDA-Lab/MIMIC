module fake_jpeg_30839_n_435 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_435);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_435;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_7),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_46),
.Y(n_144)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_52),
.Y(n_134)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_53),
.Y(n_143)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_14),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_61),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx10_ASAP7_75t_R g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_14),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_13),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_71),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_72),
.B(n_74),
.Y(n_129)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_75),
.B(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_11),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_76),
.B(n_79),
.Y(n_123)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_77),
.Y(n_133)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_11),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_23),
.B(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_10),
.C(n_1),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_29),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_84),
.B(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_35),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_31),
.A2(n_38),
.B1(n_28),
.B2(n_33),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_32),
.B1(n_26),
.B2(n_33),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_36),
.B(n_41),
.C(n_17),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_94),
.A2(n_107),
.B(n_6),
.C(n_8),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_38),
.B1(n_32),
.B2(n_35),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_98),
.B(n_111),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_102),
.B(n_142),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_37),
.B1(n_30),
.B2(n_44),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_110),
.B1(n_114),
.B2(n_126),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_33),
.B1(n_28),
.B2(n_44),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_104),
.A2(n_131),
.B1(n_137),
.B2(n_105),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_91),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_26),
.B(n_41),
.C(n_19),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_37),
.B1(n_30),
.B2(n_44),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_57),
.A2(n_33),
.B1(n_28),
.B2(n_40),
.Y(n_114)
);

AND2x4_ASAP7_75t_SL g117 ( 
.A(n_61),
.B(n_72),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_120),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_40),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_SL g184 ( 
.A(n_118),
.B(n_132),
.C(n_102),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_29),
.B1(n_42),
.B2(n_45),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_60),
.A2(n_42),
.B1(n_29),
.B2(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_R g132 ( 
.A(n_76),
.B(n_42),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_42),
.B1(n_1),
.B2(n_3),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_138),
.B1(n_140),
.B2(n_6),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_65),
.A2(n_42),
.B1(n_3),
.B2(n_4),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_68),
.A2(n_69),
.B1(n_90),
.B2(n_89),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_75),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_79),
.B(n_0),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_147),
.B(n_148),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g219 ( 
.A(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_151),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_152),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_80),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_159),
.B(n_185),
.CI(n_186),
.CON(n_204),
.SN(n_204)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_66),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_161),
.B(n_168),
.C(n_177),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_0),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_172),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_163),
.B(n_171),
.Y(n_228)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_91),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_111),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_95),
.B(n_8),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_8),
.B1(n_9),
.B2(n_121),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_121),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_178),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_101),
.B(n_9),
.C(n_107),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_106),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_182),
.Y(n_237)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_98),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_125),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_94),
.A2(n_141),
.B(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_104),
.A2(n_120),
.B1(n_139),
.B2(n_143),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_114),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_122),
.C(n_100),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_99),
.B1(n_108),
.B2(n_116),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_124),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_192),
.B(n_144),
.Y(n_227)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_108),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_144),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_183),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_108),
.B1(n_116),
.B2(n_97),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_231),
.B1(n_233),
.B2(n_187),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_200),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_126),
.B1(n_138),
.B2(n_145),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_159),
.B1(n_167),
.B2(n_166),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_171),
.A2(n_135),
.B(n_124),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_207),
.A2(n_232),
.B(n_209),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_162),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_224),
.B(n_227),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_172),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_168),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_116),
.B1(n_112),
.B2(n_115),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_182),
.A2(n_115),
.B1(n_122),
.B2(n_145),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_158),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_245),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_152),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_248),
.Y(n_282)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_202),
.A2(n_188),
.B1(n_149),
.B2(n_153),
.Y(n_245)
);

A2O1A1O1Ixp25_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_185),
.B(n_180),
.C(n_196),
.D(n_149),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_246),
.A2(n_278),
.B(n_220),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_177),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_247),
.B(n_255),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_202),
.A2(n_149),
.B1(n_159),
.B2(n_161),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_249),
.A2(n_252),
.B1(n_259),
.B2(n_208),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_254),
.B1(n_207),
.B2(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_160),
.B1(n_165),
.B2(n_155),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_257),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_229),
.B1(n_203),
.B2(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_226),
.B(n_148),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_146),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_210),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_179),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_262),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_175),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_197),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_195),
.C(n_193),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_275),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_201),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_150),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_211),
.Y(n_268)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_210),
.A2(n_100),
.B(n_156),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_234),
.B(n_220),
.Y(n_286)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_204),
.B(n_200),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_235),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_208),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_281),
.B(n_289),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_294),
.B1(n_304),
.B2(n_250),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

NAND2x1_ASAP7_75t_SL g291 ( 
.A(n_245),
.B(n_217),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_291),
.A2(n_300),
.B(n_275),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_292),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_243),
.A2(n_240),
.B1(n_234),
.B2(n_221),
.Y(n_294)
);

AOI22x1_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_219),
.B1(n_217),
.B2(n_230),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_298),
.A2(n_219),
.B(n_255),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_230),
.C(n_215),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_303),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_272),
.A2(n_221),
.B(n_223),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_223),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_245),
.A2(n_225),
.B1(n_219),
.B2(n_206),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_241),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_307),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_252),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_244),
.B(n_225),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_271),
.Y(n_334)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_259),
.B1(n_249),
.B2(n_257),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_313),
.A2(n_330),
.B1(n_331),
.B2(n_296),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_314),
.A2(n_310),
.B1(n_297),
.B2(n_293),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_300),
.A2(n_247),
.B(n_263),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_327),
.Y(n_352)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_307),
.B(n_254),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_322),
.Y(n_340)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_296),
.A2(n_284),
.B1(n_304),
.B2(n_294),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_323),
.A2(n_286),
.B1(n_299),
.B2(n_280),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_261),
.C(n_253),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_337),
.C(n_302),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_285),
.A2(n_303),
.B(n_296),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_242),
.C(n_266),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_329),
.B(n_285),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_281),
.A2(n_242),
.B1(n_246),
.B2(n_251),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_309),
.A2(n_258),
.B1(n_273),
.B2(n_277),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_333),
.Y(n_349)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_335),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_336),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_211),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_290),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_359),
.B1(n_314),
.B2(n_339),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_291),
.B1(n_298),
.B2(n_305),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_342),
.A2(n_344),
.B1(n_335),
.B2(n_321),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_343),
.B(n_351),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_317),
.A2(n_291),
.B1(n_298),
.B2(n_305),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_306),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_355),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_347),
.A2(n_353),
.B1(n_320),
.B2(n_338),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_293),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_327),
.Y(n_373)
);

NOR4xp25_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_280),
.C(n_302),
.D(n_297),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_362),
.C(n_363),
.Y(n_367)
);

OAI21xp33_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_317),
.B(n_326),
.Y(n_355)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_358),
.Y(n_371)
);

NOR4xp25_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_282),
.C(n_290),
.D(n_301),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_282),
.Y(n_361)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_361),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_311),
.C(n_283),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_311),
.C(n_283),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_350),
.Y(n_364)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_365),
.A2(n_368),
.B1(n_360),
.B2(n_340),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_350),
.Y(n_366)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_316),
.B1(n_323),
.B2(n_333),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_348),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_373),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_334),
.Y(n_372)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_349),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_382),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_375),
.A2(n_380),
.B1(n_345),
.B2(n_356),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_312),
.C(n_316),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_362),
.C(n_352),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_377),
.A2(n_335),
.B1(n_360),
.B2(n_340),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_331),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_342),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_343),
.A2(n_319),
.B1(n_332),
.B2(n_322),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_383),
.B(n_384),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_344),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_345),
.C(n_341),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_367),
.C(n_370),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_393),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_390),
.A2(n_392),
.B1(n_368),
.B2(n_365),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_391),
.A2(n_377),
.B1(n_379),
.B2(n_373),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_335),
.C(n_357),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_396),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_357),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_397),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_398),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_401),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_400),
.B(n_383),
.Y(n_411)
);

AO221x1_ASAP7_75t_L g401 ( 
.A1(n_385),
.A2(n_382),
.B1(n_301),
.B2(n_325),
.C(n_364),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_397),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_404),
.B(n_386),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_405),
.A2(n_389),
.B1(n_394),
.B2(n_392),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_369),
.C(n_372),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_395),
.C(n_396),
.Y(n_416)
);

OAI322xp33_ASAP7_75t_L g408 ( 
.A1(n_387),
.A2(n_366),
.A3(n_325),
.B1(n_308),
.B2(n_270),
.C1(n_268),
.C2(n_265),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g417 ( 
.A1(n_408),
.A2(n_325),
.B(n_214),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_414),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_412),
.A2(n_399),
.B1(n_402),
.B2(n_410),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_393),
.Y(n_415)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_415),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_416),
.B(n_400),
.C(n_406),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_405),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_403),
.A2(n_395),
.B1(n_325),
.B2(n_214),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_418),
.B(n_419),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_409),
.B(n_403),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_423),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_410),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_427),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_420),
.B(n_413),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_429),
.B(n_415),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_421),
.B(n_422),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_431),
.B(n_426),
.C(n_416),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_432),
.A2(n_423),
.B(n_430),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_425),
.C(n_412),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g435 ( 
.A(n_434),
.Y(n_435)
);


endmodule