module fake_jpeg_16946_n_215 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_38),
.Y(n_39)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_16),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_17),
.B1(n_26),
.B2(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_29),
.B1(n_26),
.B2(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_38),
.B1(n_29),
.B2(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_37),
.C(n_22),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_18),
.C(n_19),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_14),
.B1(n_23),
.B2(n_26),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_69),
.B1(n_29),
.B2(n_43),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_31),
.B1(n_35),
.B2(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_15),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_48),
.B1(n_59),
.B2(n_65),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_43),
.B(n_35),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_57),
.B(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_91),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_75),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_100),
.B(n_102),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_48),
.B1(n_66),
.B2(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_108),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_20),
.B(n_19),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_105),
.B(n_25),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_20),
.B(n_15),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_59),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_44),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_79),
.B1(n_36),
.B2(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_92),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_125),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_83),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_77),
.C(n_85),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_95),
.C(n_100),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_88),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_85),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_130),
.B(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_135),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_137),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_100),
.C(n_106),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_106),
.B1(n_127),
.B2(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_126),
.B1(n_112),
.B2(n_122),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_105),
.B(n_104),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_102),
.B1(n_105),
.B2(n_107),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_130),
.B1(n_109),
.B2(n_98),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_147),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_104),
.A3(n_112),
.B1(n_109),
.B2(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_112),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_119),
.B1(n_128),
.B2(n_126),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_155),
.B1(n_156),
.B2(n_161),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_98),
.B1(n_77),
.B2(n_81),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_86),
.B1(n_76),
.B2(n_49),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_135),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_138),
.B(n_137),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_76),
.B1(n_33),
.B2(n_28),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_76),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_134),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_158),
.B(n_154),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_171),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_157),
.C(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_172),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_132),
.C(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_34),
.C(n_33),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_131),
.B1(n_145),
.B2(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_175),
.B1(n_1),
.B2(n_2),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_178),
.C(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_181),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_49),
.C(n_36),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_36),
.C(n_34),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_52),
.C(n_5),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_34),
.C(n_33),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_28),
.C(n_52),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_1),
.B(n_4),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_1),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_176),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_192),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_166),
.B1(n_171),
.B2(n_164),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_4),
.Y(n_197)
);

NAND4xp25_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_176),
.C(n_169),
.D(n_5),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_44),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_7),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_196),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_197),
.A2(n_201),
.B(n_7),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_5),
.B(n_6),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_7),
.B(n_8),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_198),
.B(n_200),
.C(n_193),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_10),
.C(n_11),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_208),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_11),
.B(n_8),
.C(n_10),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_207),
.C(n_211),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_212),
.Y(n_215)
);


endmodule