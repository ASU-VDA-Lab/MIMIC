module fake_jpeg_11803_n_622 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_622);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_622;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

OR2x2_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_4),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_9),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_1),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_62),
.B(n_69),
.Y(n_145)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_74),
.Y(n_128)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_6),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_71),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_9),
.B(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_72),
.B(n_10),
.Y(n_163)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_18),
.B(n_5),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_5),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_76),
.B(n_123),
.Y(n_146)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_18),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_111),
.Y(n_156)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_18),
.A2(n_16),
.B1(n_13),
.B2(n_11),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_84),
.A2(n_54),
.B1(n_34),
.B2(n_43),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_85),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_28),
.B(n_13),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_105),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_13),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_89),
.B(n_126),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_22),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_22),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_31),
.B(n_13),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_43),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g148 ( 
.A(n_117),
.Y(n_148)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_29),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_43),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_121),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_48),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_54),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_31),
.B(n_45),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_137),
.B(n_200),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_68),
.A2(n_34),
.B1(n_54),
.B2(n_59),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_149),
.A2(n_155),
.B1(n_60),
.B2(n_36),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_151),
.B(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_45),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_153),
.B(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_76),
.A2(n_59),
.B1(n_52),
.B2(n_44),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g161 ( 
.A(n_71),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_161),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g247 ( 
.A1(n_163),
.A2(n_182),
.B(n_202),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_70),
.B(n_46),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_183),
.Y(n_222)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_75),
.A2(n_44),
.B1(n_59),
.B2(n_52),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g241 ( 
.A1(n_173),
.A2(n_56),
.B1(n_39),
.B2(n_35),
.Y(n_241)
);

INVx6_ASAP7_75t_SL g174 ( 
.A(n_91),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_78),
.B(n_46),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_107),
.A2(n_37),
.B(n_41),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_95),
.B(n_37),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_98),
.B(n_41),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_50),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_100),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_29),
.Y(n_225)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_102),
.A2(n_120),
.B1(n_36),
.B2(n_27),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_194),
.A2(n_36),
.B1(n_27),
.B2(n_44),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_80),
.B(n_48),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_88),
.B(n_51),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_199),
.B(n_50),
.Y(n_266)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_108),
.Y(n_200)
);

HAxp5_ASAP7_75t_SL g202 ( 
.A(n_112),
.B(n_55),
.CON(n_202),
.SN(n_202)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_211),
.A2(n_245),
.B1(n_271),
.B2(n_277),
.Y(n_294)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_212),
.Y(n_325)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_213),
.Y(n_302)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_216),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_217),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_220),
.Y(n_295)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_225),
.B(n_257),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_128),
.B(n_51),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_226),
.B(n_240),
.Y(n_297)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_139),
.Y(n_229)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_232),
.Y(n_334)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_149),
.A2(n_79),
.B1(n_61),
.B2(n_64),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_233),
.B(n_197),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_235),
.Y(n_317)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_237),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_156),
.B(n_24),
.C(n_39),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_253),
.C(n_172),
.Y(n_284)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_157),
.Y(n_239)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_239),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_241),
.A2(n_276),
.B1(n_160),
.B2(n_212),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_145),
.B(n_24),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_250),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_146),
.A2(n_115),
.B1(n_65),
.B2(n_106),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_243),
.A2(n_255),
.B1(n_280),
.B2(n_129),
.Y(n_339)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_244),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_194),
.A2(n_122),
.B1(n_99),
.B2(n_94),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_56),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_146),
.A2(n_85),
.B1(n_86),
.B2(n_90),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_251),
.A2(n_264),
.B1(n_180),
.B2(n_204),
.Y(n_313)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_141),
.B(n_59),
.C(n_35),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_138),
.A2(n_35),
.B1(n_58),
.B2(n_57),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_202),
.B(n_50),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_270),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_131),
.B(n_23),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_147),
.B(n_50),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_259),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_147),
.B(n_50),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_188),
.Y(n_260)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_261),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_162),
.B(n_23),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_262),
.B(n_266),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_263),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_164),
.A2(n_23),
.B1(n_58),
.B2(n_57),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_148),
.A2(n_39),
.B(n_58),
.C(n_57),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_256),
.Y(n_286)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_133),
.A2(n_56),
.B1(n_19),
.B2(n_60),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_167),
.B(n_19),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_272),
.B(n_274),
.Y(n_331)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_138),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_278),
.Y(n_318)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_143),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

BUFx4f_ASAP7_75t_SL g309 ( 
.A(n_275),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_181),
.A2(n_50),
.B1(n_19),
.B2(n_60),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_205),
.A2(n_55),
.B1(n_11),
.B2(n_2),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_132),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_152),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_281),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_142),
.A2(n_205),
.B1(n_169),
.B2(n_135),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_161),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_154),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_220),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_284),
.B(n_300),
.C(n_321),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_286),
.A2(n_340),
.B(n_277),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_226),
.A2(n_247),
.B1(n_234),
.B2(n_243),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_288),
.A2(n_313),
.B1(n_232),
.B2(n_268),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_254),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_305),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_222),
.B(n_180),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_314),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_172),
.C(n_195),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_252),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_255),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_245),
.A2(n_135),
.B1(n_133),
.B2(n_169),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_308),
.A2(n_329),
.B1(n_333),
.B2(n_261),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_269),
.B(n_142),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_209),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_4),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_238),
.B(n_177),
.C(n_130),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_241),
.A2(n_160),
.B1(n_158),
.B2(n_140),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_237),
.A2(n_158),
.B1(n_140),
.B2(n_136),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_219),
.A2(n_177),
.B1(n_134),
.B2(n_130),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_233),
.A2(n_134),
.B1(n_129),
.B2(n_55),
.Y(n_333)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_339),
.A2(n_233),
.B1(n_273),
.B2(n_275),
.Y(n_347)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_246),
.A2(n_175),
.A3(n_55),
.B1(n_2),
.B2(n_3),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_286),
.A2(n_276),
.B(n_246),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_345),
.A2(n_387),
.B(n_318),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_233),
.B1(n_253),
.B2(n_280),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_352),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_347),
.A2(n_367),
.B1(n_382),
.B2(n_385),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g351 ( 
.A(n_284),
.B(n_214),
.CI(n_218),
.CON(n_351),
.SN(n_351)
);

FAx1_ASAP7_75t_SL g426 ( 
.A(n_351),
.B(n_309),
.CI(n_295),
.CON(n_426),
.SN(n_426)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_294),
.A2(n_223),
.B1(n_213),
.B2(n_230),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_365),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_314),
.A2(n_301),
.B(n_300),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_354),
.A2(n_302),
.B(n_307),
.Y(n_425)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_299),
.A2(n_236),
.B1(n_278),
.B2(n_216),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_356),
.A2(n_360),
.B1(n_370),
.B2(n_374),
.Y(n_389)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

OA21x2_ASAP7_75t_R g359 ( 
.A1(n_304),
.A2(n_235),
.B(n_244),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_359),
.B(n_379),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_299),
.A2(n_229),
.B1(n_270),
.B2(n_239),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_364),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_332),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_337),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_380),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_249),
.B1(n_221),
.B2(n_260),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_305),
.A2(n_210),
.B1(n_215),
.B2(n_2),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_371),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_304),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_308),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_321),
.A2(n_0),
.B1(n_4),
.B2(n_322),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_376),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_373),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_304),
.A2(n_4),
.B1(n_319),
.B2(n_335),
.Y(n_374)
);

OAI22x1_ASAP7_75t_SL g376 ( 
.A1(n_301),
.A2(n_311),
.B1(n_290),
.B2(n_292),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_377),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_301),
.B(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_378),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_298),
.B(n_320),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_297),
.B(n_291),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_292),
.A2(n_283),
.B1(n_285),
.B2(n_287),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_291),
.B(n_283),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_303),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_285),
.B(n_287),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_384),
.B(n_386),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_293),
.A2(n_318),
.B1(n_336),
.B2(n_296),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_293),
.B(n_336),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_318),
.B(n_337),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_324),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_396),
.C(n_399),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_392),
.A2(n_420),
.B(n_363),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_357),
.A2(n_334),
.B1(n_319),
.B2(n_312),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_395),
.A2(n_414),
.B1(n_364),
.B2(n_352),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_296),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_384),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_418),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_310),
.C(n_324),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_303),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_409),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_369),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_348),
.A2(n_325),
.B1(n_330),
.B2(n_335),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_408),
.A2(n_422),
.B1(n_356),
.B2(n_349),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_317),
.C(n_341),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_357),
.A2(n_334),
.B1(n_312),
.B2(n_306),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_354),
.B(n_317),
.C(n_341),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_424),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_386),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_345),
.A2(n_306),
.B(n_338),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_350),
.A2(n_325),
.B1(n_330),
.B2(n_338),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_302),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_383),
.C(n_373),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_380),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_425),
.A2(n_426),
.B(n_345),
.Y(n_433)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_411),
.Y(n_427)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_427),
.Y(n_470)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_430),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_431),
.A2(n_434),
.B(n_458),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_433),
.A2(n_454),
.B(n_412),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_392),
.A2(n_344),
.B(n_369),
.Y(n_434)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_436),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_363),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_438),
.Y(n_488)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_439),
.Y(n_477)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_441),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_401),
.B(n_379),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_442),
.B(n_443),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_423),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_444),
.Y(n_487)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_405),
.Y(n_445)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_405),
.Y(n_446)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_446),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_449),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_413),
.A2(n_347),
.B1(n_361),
.B2(n_359),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_448),
.A2(n_453),
.B1(n_403),
.B2(n_406),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_401),
.B(n_382),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_424),
.B(n_372),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_459),
.Y(n_492)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_455),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_413),
.A2(n_374),
.B1(n_346),
.B2(n_367),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_393),
.A2(n_426),
.B(n_425),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_396),
.B(n_378),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_409),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_403),
.A2(n_378),
.B1(n_363),
.B2(n_353),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_402),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_412),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_366),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_388),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_475),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_432),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_464),
.B(n_479),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_465),
.A2(n_434),
.B1(n_461),
.B2(n_416),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_453),
.A2(n_406),
.B1(n_403),
.B2(n_390),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_468),
.A2(n_482),
.B1(n_465),
.B2(n_466),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_458),
.A2(n_393),
.B1(n_410),
.B2(n_417),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_469),
.A2(n_478),
.B1(n_489),
.B2(n_438),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_473),
.A2(n_351),
.B(n_445),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_474),
.B(n_415),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_437),
.B(n_399),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_431),
.A2(n_410),
.B1(n_417),
.B2(n_407),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_435),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_448),
.A2(n_390),
.B1(n_400),
.B2(n_418),
.Y(n_482)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_455),
.A2(n_407),
.B1(n_389),
.B2(n_398),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_495),
.A2(n_502),
.B1(n_512),
.B2(n_490),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_476),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_496),
.B(n_501),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_460),
.C(n_451),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_504),
.C(n_519),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_462),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_499),
.B(n_506),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_460),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_520),
.Y(n_524)
);

NAND4xp25_ASAP7_75t_SL g501 ( 
.A(n_483),
.B(n_295),
.C(n_454),
.D(n_397),
.Y(n_501)
);

FAx1_ASAP7_75t_L g503 ( 
.A(n_469),
.B(n_433),
.CI(n_426),
.CON(n_503),
.SN(n_503)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_503),
.B(n_510),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_451),
.C(n_457),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_480),
.Y(n_505)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_505),
.Y(n_545)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_467),
.Y(n_506)
);

CKINVDCx14_ASAP7_75t_R g507 ( 
.A(n_492),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_507),
.A2(n_518),
.B1(n_429),
.B2(n_440),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_509),
.Y(n_546)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_480),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_511),
.A2(n_515),
.B1(n_491),
.B2(n_487),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_482),
.A2(n_370),
.B1(n_438),
.B2(n_452),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_486),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_513),
.B(n_517),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_478),
.B(n_415),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_484),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_489),
.A2(n_395),
.B1(n_414),
.B2(n_419),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_516),
.A2(n_351),
.B(n_485),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_427),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_484),
.C(n_473),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_481),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_521),
.B(n_508),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_488),
.B(n_351),
.C(n_444),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_522),
.B(n_342),
.C(n_470),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_523),
.B(n_527),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_468),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_525),
.B(n_526),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_494),
.B(n_466),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_529),
.A2(n_530),
.B(n_503),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_522),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_502),
.A2(n_493),
.B1(n_491),
.B2(n_487),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_539),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_494),
.B(n_477),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_534),
.B(n_535),
.C(n_519),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_498),
.B(n_477),
.Y(n_535)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_536),
.Y(n_549)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_537),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_511),
.A2(n_472),
.B1(n_441),
.B2(n_471),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_504),
.B(n_472),
.C(n_471),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_540),
.B(n_544),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_515),
.A2(n_446),
.B1(n_439),
.B2(n_436),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_501),
.Y(n_552)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_543),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_520),
.B(n_428),
.C(n_421),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_547),
.B(n_556),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_548),
.B(n_525),
.Y(n_574)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_552),
.Y(n_583)
);

FAx1_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_503),
.CI(n_536),
.CON(n_554),
.SN(n_554)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_565),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_514),
.C(n_517),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_516),
.C(n_497),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_557),
.B(n_563),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_538),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_558),
.B(n_560),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_499),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_542),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_562),
.B(n_532),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_528),
.B(n_512),
.C(n_513),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_518),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_564),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_542),
.B(n_510),
.Y(n_566)
);

INVxp33_ASAP7_75t_SL g575 ( 
.A(n_566),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_563),
.B(n_528),
.C(n_534),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_570),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_559),
.A2(n_539),
.B1(n_541),
.B2(n_531),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_571),
.B(n_572),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_549),
.A2(n_544),
.B1(n_527),
.B2(n_529),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_574),
.B(n_576),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_526),
.C(n_524),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_565),
.A2(n_523),
.B(n_524),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_578),
.A2(n_579),
.B(n_548),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_557),
.A2(n_397),
.B(n_358),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_555),
.B(n_385),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_580),
.B(n_581),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_561),
.B(n_355),
.Y(n_581)
);

AOI21x1_ASAP7_75t_L g598 ( 
.A1(n_586),
.A2(n_574),
.B(n_575),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_556),
.C(n_551),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_587),
.B(n_592),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g588 ( 
.A1(n_577),
.A2(n_582),
.B(n_583),
.Y(n_588)
);

NOR2x1_ASAP7_75t_SL g597 ( 
.A(n_588),
.B(n_576),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_577),
.A2(n_554),
.B(n_550),
.Y(n_590)
);

AOI21xp33_ASAP7_75t_L g601 ( 
.A1(n_590),
.A2(n_594),
.B(n_368),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_569),
.B(n_550),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_567),
.B(n_566),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_593),
.B(n_570),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_572),
.A2(n_554),
.B(n_552),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_575),
.A2(n_566),
.B1(n_555),
.B2(n_551),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_595),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_573),
.B(n_349),
.C(n_381),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_362),
.C(n_377),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_597),
.B(n_598),
.C(n_599),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_580),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_600),
.B(n_602),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_601),
.B(n_603),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_589),
.B(n_343),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_584),
.B(n_430),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_604),
.B(n_591),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_605),
.A2(n_594),
.B(n_590),
.Y(n_607)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_607),
.Y(n_616)
);

AO21x1_ASAP7_75t_L g613 ( 
.A1(n_608),
.A2(n_606),
.B(n_595),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_SL g612 ( 
.A1(n_606),
.A2(n_587),
.B(n_585),
.Y(n_612)
);

AOI21xp33_ASAP7_75t_L g615 ( 
.A1(n_612),
.A2(n_309),
.B(n_387),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_613),
.A2(n_615),
.B(n_616),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_609),
.A2(n_610),
.B1(n_611),
.B2(n_602),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_614),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_618),
.A2(n_342),
.B(n_387),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_619),
.B(n_617),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_620),
.A2(n_387),
.B(n_307),
.Y(n_621)
);

FAx1_ASAP7_75t_SL g622 ( 
.A(n_621),
.B(n_371),
.CI(n_614),
.CON(n_622),
.SN(n_622)
);


endmodule