module fake_jpeg_17844_n_347 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_23),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_0),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_26),
.Y(n_68)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_24),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_49),
.B1(n_40),
.B2(n_20),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_23),
.B1(n_19),
.B2(n_35),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_62),
.B1(n_49),
.B2(n_48),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_23),
.B1(n_19),
.B2(n_35),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_34),
.C(n_36),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_34),
.C(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_64),
.B(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_23),
.B1(n_19),
.B2(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_44),
.B1(n_22),
.B2(n_33),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_51),
.B(n_45),
.C(n_42),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_32),
.B(n_29),
.C(n_27),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_92),
.B1(n_58),
.B2(n_34),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_98),
.B1(n_102),
.B2(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_20),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_100),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_101),
.C(n_52),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_33),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_18),
.B(n_25),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_37),
.B1(n_32),
.B2(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_99),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_50),
.B1(n_43),
.B2(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_33),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_50),
.C(n_43),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_50),
.B1(n_43),
.B2(n_22),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_32),
.B1(n_37),
.B2(n_18),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_72),
.B1(n_66),
.B2(n_70),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_133),
.B1(n_134),
.B2(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_25),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_121),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_52),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_69),
.B1(n_60),
.B2(n_50),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_128),
.B1(n_132),
.B2(n_34),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_120),
.A2(n_127),
.B(n_34),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_18),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_27),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_86),
.B(n_65),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_60),
.B1(n_65),
.B2(n_52),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_98),
.B1(n_102),
.B2(n_93),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_129),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_1),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_79),
.B(n_82),
.C(n_29),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_58),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_93),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_78),
.B1(n_92),
.B2(n_103),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_36),
.B1(n_30),
.B2(n_29),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_82),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_142),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_148),
.B1(n_151),
.B2(n_157),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_94),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_117),
.B(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_156),
.Y(n_177)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_79),
.B1(n_88),
.B2(n_93),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_160),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_88),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_71),
.B1(n_36),
.B2(n_30),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_71),
.B1(n_36),
.B2(n_30),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_127),
.B1(n_134),
.B2(n_133),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_2),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_74),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_124),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_31),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_165),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_131),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_117),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_151),
.C(n_162),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_107),
.A3(n_122),
.B1(n_117),
.B2(n_118),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_185),
.Y(n_219)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_189),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_31),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_109),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_186),
.B1(n_194),
.B2(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_118),
.B1(n_127),
.B2(n_112),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_144),
.B(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_121),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_140),
.B(n_119),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_130),
.B(n_120),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_195),
.B(n_2),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_164),
.A2(n_125),
.B1(n_130),
.B2(n_128),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_143),
.A2(n_34),
.B(n_31),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_139),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

AOI22x1_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_153),
.B1(n_141),
.B2(n_145),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_198),
.A2(n_203),
.B1(n_192),
.B2(n_181),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_211),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_150),
.B1(n_147),
.B2(n_140),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_215),
.B1(n_218),
.B2(n_196),
.Y(n_240)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_206),
.C(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_186),
.C(n_175),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_163),
.C(n_160),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_207),
.B(n_223),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_147),
.A3(n_144),
.B1(n_139),
.B2(n_161),
.C1(n_157),
.C2(n_158),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_176),
.B(n_168),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_155),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_217),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_142),
.C(n_137),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_146),
.B1(n_154),
.B2(n_2),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_154),
.B1(n_3),
.B2(n_2),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_105),
.C(n_31),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_194),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_224),
.A2(n_3),
.B(n_4),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_189),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_174),
.Y(n_228)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_205),
.C(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_202),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_233),
.A2(n_238),
.B(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

XNOR2x2_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_177),
.Y(n_238)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_182),
.B1(n_183),
.B2(n_170),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_177),
.B(n_191),
.C(n_180),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_246),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_172),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_252),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_201),
.A2(n_195),
.B1(n_170),
.B2(n_187),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_253),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_220),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_105),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_105),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_248),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_274),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_223),
.C(n_200),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_268),
.C(n_273),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_210),
.B1(n_218),
.B2(n_207),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_247),
.B1(n_240),
.B2(n_231),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_221),
.C(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_3),
.C(n_4),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_10),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_230),
.B(n_10),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_277),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_237),
.B(n_246),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_256),
.B(n_267),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_234),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_289),
.C(n_295),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_235),
.B1(n_250),
.B2(n_245),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_286),
.B1(n_265),
.B2(n_259),
.Y(n_308)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_233),
.B1(n_236),
.B2(n_242),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_288),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_234),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_255),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_243),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_266),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_231),
.C(n_249),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_SL g299 ( 
.A(n_294),
.B(n_270),
.C(n_263),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_9),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_272),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_299),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_305),
.B1(n_278),
.B2(n_304),
.Y(n_312)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_268),
.C(n_262),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_274),
.C(n_254),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_254),
.C(n_267),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_284),
.A2(n_276),
.B1(n_256),
.B2(n_265),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_260),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_310),
.C(n_295),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_273),
.C(n_3),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_286),
.A2(n_5),
.B(n_6),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_5),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_312),
.B(n_313),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_302),
.B1(n_279),
.B2(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_315),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_301),
.B(n_281),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_316),
.B(n_318),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_319),
.B(n_320),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_296),
.B(n_6),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_7),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_297),
.Y(n_325)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_323),
.B(n_322),
.Y(n_328)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_7),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_9),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_323),
.C(n_14),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_332),
.C(n_12),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

AOI21xp33_ASAP7_75t_L g342 ( 
.A1(n_335),
.A2(n_333),
.B(n_301),
.Y(n_342)
);

AOI31xp67_ASAP7_75t_L g338 ( 
.A1(n_327),
.A2(n_17),
.A3(n_12),
.B(n_16),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_17),
.B(n_337),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_325),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_340),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_342),
.B(n_336),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_343),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_344),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_346),
.Y(n_347)
);


endmodule