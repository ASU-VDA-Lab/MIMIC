module fake_jpeg_30477_n_103 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_18),
.B(n_25),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_46),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_0),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_1),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_36),
.B1(n_39),
.B2(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_59),
.B1(n_7),
.B2(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_2),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_36),
.B(n_39),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_10),
.B(n_11),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_40),
.B1(n_31),
.B2(n_16),
.Y(n_59)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_15),
.C(n_30),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_54),
.C(n_17),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_71)
);

NAND2x1_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_4),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_6),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_9),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_13),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_14),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_74),
.C(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_71),
.B1(n_63),
.B2(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_84),
.B1(n_90),
.B2(n_82),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_78),
.B1(n_81),
.B2(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_92),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_88),
.B1(n_80),
.B2(n_86),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_80),
.B1(n_26),
.B2(n_27),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_21),
.Y(n_103)
);


endmodule