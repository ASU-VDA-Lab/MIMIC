module real_aes_5884_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_904;
wire n_683;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_298;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_266;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_0), .A2(n_97), .B1(n_521), .B2(n_523), .Y(n_520) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_1), .Y(n_649) );
AND2x4_ASAP7_75t_L g663 ( .A(n_1), .B(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g672 ( .A(n_1), .B(n_239), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_2), .A2(n_202), .B1(n_419), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_3), .A2(n_108), .B1(n_675), .B2(n_688), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_4), .A2(n_143), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g625 ( .A(n_5), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_6), .A2(n_46), .B1(n_533), .B2(n_534), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_7), .A2(n_15), .B1(n_360), .B2(n_362), .Y(n_359) );
AOI21xp33_ASAP7_75t_L g309 ( .A1(n_8), .A2(n_310), .B(n_311), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_9), .A2(n_94), .B1(n_384), .B2(n_386), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_10), .A2(n_158), .B1(n_336), .B2(n_337), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_11), .A2(n_102), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_12), .A2(n_368), .B(n_370), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_13), .A2(n_245), .B1(n_325), .B2(n_333), .Y(n_397) );
XNOR2x2_ASAP7_75t_L g619 ( .A(n_14), .B(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_16), .Y(n_673) );
AO22x2_ASAP7_75t_L g687 ( .A1(n_17), .A2(n_59), .B1(n_675), .B2(n_688), .Y(n_687) );
AO22x1_ASAP7_75t_L g689 ( .A1(n_18), .A2(n_248), .B1(n_690), .B2(n_692), .Y(n_689) );
INVxp33_ASAP7_75t_SL g724 ( .A(n_19), .Y(n_724) );
INVx1_ASAP7_75t_L g928 ( .A(n_20), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_21), .A2(n_72), .B1(n_362), .B2(n_415), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_22), .A2(n_68), .B1(n_332), .B2(n_336), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_23), .A2(n_57), .B1(n_360), .B2(n_523), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_24), .A2(n_187), .B1(n_373), .B2(n_375), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_25), .A2(n_39), .B1(n_445), .B2(n_526), .C(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g410 ( .A(n_26), .Y(n_410) );
INVx1_ASAP7_75t_L g529 ( .A(n_27), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_28), .A2(n_155), .B1(n_362), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_29), .A2(n_104), .B1(n_671), .B2(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g279 ( .A(n_30), .Y(n_279) );
INVxp67_ASAP7_75t_L g289 ( .A(n_30), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_30), .B(n_183), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_31), .A2(n_192), .B1(n_665), .B2(n_675), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_32), .A2(n_106), .B1(n_690), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_33), .A2(n_42), .B1(n_329), .B2(n_330), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_34), .A2(n_122), .B1(n_296), .B2(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g500 ( .A(n_35), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_36), .A2(n_87), .B1(n_344), .B2(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_37), .B(n_263), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_38), .A2(n_213), .B1(n_360), .B2(n_362), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_40), .A2(n_85), .B1(n_533), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_41), .A2(n_238), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_43), .A2(n_190), .B1(n_282), .B2(n_324), .Y(n_497) );
INVx1_ASAP7_75t_L g886 ( .A(n_44), .Y(n_886) );
AOI21xp33_ASAP7_75t_L g498 ( .A1(n_45), .A2(n_409), .B(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_47), .A2(n_229), .B1(n_415), .B2(n_523), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_48), .A2(n_211), .B1(n_688), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_49), .A2(n_124), .B1(n_360), .B2(n_362), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_50), .A2(n_147), .B1(n_292), .B2(n_296), .Y(n_496) );
INVx2_ASAP7_75t_L g647 ( .A(n_51), .Y(n_647) );
INVx1_ASAP7_75t_L g882 ( .A(n_52), .Y(n_882) );
INVxp33_ASAP7_75t_SL g676 ( .A(n_53), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_54), .A2(n_114), .B1(n_344), .B2(n_481), .Y(n_623) );
INVx1_ASAP7_75t_L g662 ( .A(n_55), .Y(n_662) );
AND2x4_ASAP7_75t_L g668 ( .A(n_55), .B(n_647), .Y(n_668) );
INVx1_ASAP7_75t_SL g691 ( .A(n_55), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_56), .A2(n_88), .B1(n_344), .B2(n_900), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_58), .A2(n_180), .B1(n_428), .B2(n_917), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_60), .A2(n_84), .B1(n_282), .B2(n_292), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_61), .A2(n_173), .B1(n_351), .B2(n_583), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_62), .A2(n_210), .B1(n_344), .B2(n_423), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_63), .A2(n_148), .B1(n_422), .B2(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g476 ( .A(n_64), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_65), .A2(n_156), .B1(n_598), .B2(n_601), .Y(n_597) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_66), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_67), .A2(n_71), .B1(n_419), .B2(n_518), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_69), .A2(n_243), .B1(n_430), .B2(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g594 ( .A(n_70), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_73), .A2(n_118), .B1(n_355), .B2(n_357), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_74), .A2(n_236), .B1(n_344), .B2(n_346), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_75), .A2(n_100), .B1(n_332), .B2(n_336), .Y(n_398) );
INVx1_ASAP7_75t_L g264 ( .A(n_76), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_76), .B(n_182), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_77), .A2(n_159), .B1(n_930), .B2(n_931), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_78), .A2(n_152), .B1(n_444), .B2(n_446), .Y(n_443) );
OAI22x1_ASAP7_75t_L g341 ( .A1(n_79), .A2(n_342), .B1(n_364), .B2(n_388), .Y(n_341) );
NAND5xp2_ASAP7_75t_SL g342 ( .A(n_79), .B(n_343), .C(n_348), .D(n_354), .E(n_359), .Y(n_342) );
INVx1_ASAP7_75t_L g630 ( .A(n_80), .Y(n_630) );
AO22x1_ASAP7_75t_L g572 ( .A1(n_81), .A2(n_98), .B1(n_471), .B2(n_573), .Y(n_572) );
AOI21xp5_ASAP7_75t_SL g924 ( .A1(n_82), .A2(n_925), .B(n_927), .Y(n_924) );
XNOR2x1_ASAP7_75t_L g254 ( .A(n_83), .B(n_255), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_83), .A2(n_131), .B1(n_675), .B2(n_688), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_86), .B(n_445), .Y(n_468) );
AO221x2_ASAP7_75t_L g657 ( .A1(n_89), .A2(n_90), .B1(n_658), .B2(n_665), .C(n_669), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_89), .A2(n_911), .B1(n_934), .B2(n_937), .Y(n_910) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_89), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_91), .B(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_92), .A2(n_113), .B1(n_449), .B2(n_473), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_93), .A2(n_246), .B1(n_660), .B2(n_688), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_95), .A2(n_212), .B1(n_351), .B2(n_428), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_96), .A2(n_161), .B1(n_349), .B2(n_351), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_99), .A2(n_216), .B1(n_332), .B2(n_333), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_101), .A2(n_402), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_103), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_105), .B(n_306), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_107), .A2(n_127), .B1(n_415), .B2(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g542 ( .A(n_108), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_109), .A2(n_140), .B1(n_357), .B2(n_428), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_110), .A2(n_166), .B1(n_329), .B2(n_330), .Y(n_505) );
INVx1_ASAP7_75t_L g312 ( .A(n_111), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_112), .A2(n_223), .B1(n_344), .B2(n_346), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_115), .A2(n_203), .B1(n_355), .B2(n_357), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_116), .A2(n_128), .B1(n_423), .B2(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_117), .A2(n_172), .B1(n_536), .B2(n_539), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_119), .A2(n_186), .B1(n_690), .B2(n_697), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_120), .A2(n_228), .B1(n_324), .B2(n_325), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_121), .A2(n_150), .B1(n_425), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_123), .A2(n_146), .B1(n_449), .B2(n_534), .Y(n_636) );
INVx1_ASAP7_75t_L g371 ( .A(n_125), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_126), .A2(n_193), .B1(n_292), .B2(n_296), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_129), .A2(n_184), .B1(n_325), .B2(n_333), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_130), .A2(n_132), .B1(n_346), .B2(n_357), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_133), .A2(n_178), .B1(n_355), .B2(n_430), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_134), .A2(n_160), .B1(n_448), .B2(n_450), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_135), .A2(n_234), .B1(n_415), .B2(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_136), .A2(n_244), .B1(n_346), .B2(n_430), .Y(n_918) );
INVx1_ASAP7_75t_L g880 ( .A(n_137), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_138), .A2(n_214), .B1(n_258), .B2(n_337), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_139), .A2(n_220), .B1(n_258), .B2(n_337), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_141), .A2(n_235), .B1(n_423), .B2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_142), .A2(n_174), .B1(n_418), .B2(n_420), .Y(n_417) );
XNOR2x1_ASAP7_75t_L g465 ( .A(n_144), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g887 ( .A(n_145), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_149), .A2(n_176), .B1(n_660), .B2(n_671), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_151), .A2(n_196), .B1(n_258), .B2(n_282), .Y(n_257) );
INVx1_ASAP7_75t_L g555 ( .A(n_153), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_154), .A2(n_217), .B1(n_533), .B2(n_575), .Y(n_574) );
OA22x2_ASAP7_75t_L g269 ( .A1(n_157), .A2(n_183), .B1(n_263), .B2(n_267), .Y(n_269) );
INVx1_ASAP7_75t_L g301 ( .A(n_157), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_162), .A2(n_197), .B1(n_470), .B2(n_638), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_163), .A2(n_204), .B1(n_551), .B2(n_553), .C(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g406 ( .A(n_164), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_165), .A2(n_433), .B(n_436), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_167), .A2(n_225), .B1(n_357), .B2(n_428), .Y(n_516) );
AOI221x1_ASAP7_75t_L g592 ( .A1(n_168), .A2(n_207), .B1(n_384), .B2(n_435), .C(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_169), .A2(n_175), .B1(n_349), .B2(n_351), .Y(n_606) );
INVx1_ASAP7_75t_L g442 ( .A(n_170), .Y(n_442) );
INVx1_ASAP7_75t_L g439 ( .A(n_171), .Y(n_439) );
INVx1_ASAP7_75t_L g719 ( .A(n_177), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_179), .A2(n_191), .B1(n_660), .B2(n_692), .Y(n_705) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_181), .A2(n_412), .B1(n_452), .B2(n_453), .Y(n_411) );
INVx1_ASAP7_75t_L g453 ( .A(n_181), .Y(n_453) );
INVx1_ASAP7_75t_L g281 ( .A(n_182), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_182), .B(n_299), .Y(n_321) );
OAI21xp33_ASAP7_75t_L g302 ( .A1(n_183), .A2(n_198), .B(n_290), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_185), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_188), .A2(n_205), .B1(n_386), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_189), .A2(n_222), .B1(n_349), .B2(n_351), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_194), .A2(n_209), .B1(n_375), .B2(n_559), .Y(n_558) );
INVx1_ASAP7_75t_SL g720 ( .A(n_195), .Y(n_720) );
INVx1_ASAP7_75t_L g266 ( .A(n_198), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_198), .B(n_231), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_199), .A2(n_227), .B1(n_329), .B2(n_330), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g875 ( .A1(n_200), .A2(n_876), .B1(n_904), .B2(n_905), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_200), .Y(n_904) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_201), .A2(n_306), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g491 ( .A(n_206), .Y(n_491) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_208), .A2(n_590), .B(n_612), .Y(n_589) );
INVx1_ASAP7_75t_L g615 ( .A(n_208), .Y(n_615) );
INVx1_ASAP7_75t_L g890 ( .A(n_215), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g722 ( .A(n_218), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_219), .B(n_553), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_221), .A2(n_224), .B1(n_427), .B2(n_429), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_226), .A2(n_242), .B1(n_386), .B2(n_533), .Y(n_560) );
AOI22x1_ASAP7_75t_L g932 ( .A1(n_230), .A2(n_237), .B1(n_470), .B2(n_534), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_231), .B(n_274), .Y(n_273) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_232), .A2(n_324), .B(n_405), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_233), .A2(n_240), .B1(n_428), .B2(n_430), .Y(n_622) );
INVx1_ASAP7_75t_L g664 ( .A(n_239), .Y(n_664) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_239), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_241), .B(n_379), .Y(n_378) );
XNOR2x1_ASAP7_75t_L g511 ( .A(n_246), .B(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_247), .A2(n_570), .B(n_572), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_650), .B(n_653), .Y(n_249) );
AOI21xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_459), .B(n_642), .Y(n_250) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_251), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_338), .B1(n_455), .B2(n_456), .Y(n_251) );
INVx2_ASAP7_75t_L g455 ( .A(n_252), .Y(n_455) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2x1_ASAP7_75t_L g255 ( .A(n_256), .B(n_322), .Y(n_255) );
NAND4xp25_ASAP7_75t_L g256 ( .A(n_257), .B(n_291), .C(n_305), .D(n_309), .Y(n_256) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_270), .Y(n_258) );
AND2x4_ASAP7_75t_L g329 ( .A(n_259), .B(n_294), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_259), .B(n_303), .Y(n_330) );
AND2x4_ASAP7_75t_L g332 ( .A(n_259), .B(n_326), .Y(n_332) );
AND2x4_ASAP7_75t_L g345 ( .A(n_259), .B(n_334), .Y(n_345) );
AND2x4_ASAP7_75t_L g350 ( .A(n_259), .B(n_326), .Y(n_350) );
AND2x4_ASAP7_75t_L g361 ( .A(n_259), .B(n_294), .Y(n_361) );
AND2x2_ASAP7_75t_L g363 ( .A(n_259), .B(n_303), .Y(n_363) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_268), .Y(n_259) );
AND2x2_ASAP7_75t_L g308 ( .A(n_260), .B(n_269), .Y(n_308) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g293 ( .A(n_261), .B(n_269), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
NAND2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g267 ( .A(n_263), .Y(n_267) );
INVx3_ASAP7_75t_L g274 ( .A(n_263), .Y(n_274) );
NAND2xp33_ASAP7_75t_L g280 ( .A(n_263), .B(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
INVx1_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_264), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_266), .A2(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g287 ( .A(n_269), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g358 ( .A(n_270), .B(n_293), .Y(n_358) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g334 ( .A(n_271), .Y(n_334) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
AND2x2_ASAP7_75t_L g283 ( .A(n_272), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g294 ( .A(n_272), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g304 ( .A(n_272), .Y(n_304) );
AND2x4_ASAP7_75t_L g326 ( .A(n_272), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_274), .B(n_279), .Y(n_278) );
INVxp67_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_275), .B(n_298), .C(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_287), .Y(n_282) );
AND2x4_ASAP7_75t_L g377 ( .A(n_283), .B(n_287), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g316 ( .A(n_285), .Y(n_316) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g310 ( .A(n_293), .B(n_303), .Y(n_310) );
AND2x4_ASAP7_75t_L g325 ( .A(n_293), .B(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g333 ( .A(n_293), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g356 ( .A(n_293), .B(n_326), .Y(n_356) );
AND2x2_ASAP7_75t_L g374 ( .A(n_293), .B(n_294), .Y(n_374) );
AND2x2_ASAP7_75t_L g382 ( .A(n_293), .B(n_303), .Y(n_382) );
AND2x2_ASAP7_75t_L g485 ( .A(n_293), .B(n_326), .Y(n_485) );
AND2x4_ASAP7_75t_L g324 ( .A(n_294), .B(n_308), .Y(n_324) );
AND2x4_ASAP7_75t_L g369 ( .A(n_294), .B(n_308), .Y(n_369) );
AND2x4_ASAP7_75t_L g303 ( .A(n_295), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_303), .Y(n_296) );
AND2x4_ASAP7_75t_L g336 ( .A(n_297), .B(n_326), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_297), .B(n_334), .Y(n_337) );
AND2x4_ASAP7_75t_L g347 ( .A(n_297), .B(n_334), .Y(n_347) );
AND2x4_ASAP7_75t_L g353 ( .A(n_297), .B(n_326), .Y(n_353) );
AND2x4_ASAP7_75t_L g387 ( .A(n_297), .B(n_303), .Y(n_387) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x4_ASAP7_75t_L g307 ( .A(n_303), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g409 ( .A(n_303), .B(n_308), .Y(n_409) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g385 ( .A(n_307), .Y(n_385) );
BUFx8_ASAP7_75t_SL g445 ( .A(n_307), .Y(n_445) );
INVx2_ASAP7_75t_L g552 ( .A(n_307), .Y(n_552) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_307), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_313), .B(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_313), .B(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g557 ( .A(n_313), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_313), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g895 ( .A(n_313), .Y(n_895) );
INVx4_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g407 ( .A(n_314), .Y(n_407) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_315), .Y(n_478) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B(n_320), .Y(n_315) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_317), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND4xp25_ASAP7_75t_L g322 ( .A(n_323), .B(n_328), .C(n_331), .D(n_335), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_411), .B2(n_454), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_339), .A2(n_454), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_339), .Y(n_457) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
XNOR2x1_ASAP7_75t_L g340 ( .A(n_341), .B(n_392), .Y(n_340) );
NAND4xp25_ASAP7_75t_L g389 ( .A(n_343), .B(n_348), .C(n_359), .D(n_378), .Y(n_389) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_345), .Y(n_419) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_345), .Y(n_487) );
BUFx3_ASAP7_75t_L g420 ( .A(n_346), .Y(n_420) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx6_ASAP7_75t_L g482 ( .A(n_347), .Y(n_482) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_350), .Y(n_423) );
BUFx12f_ASAP7_75t_L g518 ( .A(n_350), .Y(n_518) );
INVx4_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g425 ( .A(n_352), .Y(n_425) );
INVx2_ASAP7_75t_SL g519 ( .A(n_352), .Y(n_519) );
INVx4_ASAP7_75t_L g634 ( .A(n_352), .Y(n_634) );
INVx4_ASAP7_75t_L g917 ( .A(n_352), .Y(n_917) );
INVx8_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_354), .B(n_383), .Y(n_391) );
BUFx8_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_356), .Y(n_428) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx12f_ASAP7_75t_L g430 ( .A(n_358), .Y(n_430) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx12f_ASAP7_75t_L g415 ( .A(n_361), .Y(n_415) );
INVx3_ASAP7_75t_L g522 ( .A(n_361), .Y(n_522) );
BUFx3_ASAP7_75t_L g416 ( .A(n_362), .Y(n_416) );
BUFx5_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx3_ASAP7_75t_L g489 ( .A(n_363), .Y(n_489) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_363), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_378), .C(n_383), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g390 ( .A(n_366), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_372), .Y(n_366) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g449 ( .A(n_369), .Y(n_449) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_369), .Y(n_533) );
INVx1_ASAP7_75t_L g926 ( .A(n_369), .Y(n_926) );
INVx2_ASAP7_75t_L g451 ( .A(n_373), .Y(n_451) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_374), .Y(n_470) );
INVx2_ASAP7_75t_L g538 ( .A(n_374), .Y(n_538) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g438 ( .A(n_376), .Y(n_438) );
INVx4_ASAP7_75t_L g534 ( .A(n_376), .Y(n_534) );
INVx3_ASAP7_75t_L g601 ( .A(n_376), .Y(n_601) );
INVx5_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx2_ASAP7_75t_L g471 ( .A(n_377), .Y(n_471) );
BUFx4f_ASAP7_75t_L g894 ( .A(n_377), .Y(n_894) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g435 ( .A(n_380), .Y(n_435) );
INVx2_ASAP7_75t_L g627 ( .A(n_380), .Y(n_627) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g495 ( .A(n_381), .Y(n_495) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g402 ( .A(n_382), .Y(n_402) );
INVx3_ASAP7_75t_L g527 ( .A(n_382), .Y(n_527) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g446 ( .A(n_386), .Y(n_446) );
INVx4_ASAP7_75t_L g888 ( .A(n_386), .Y(n_888) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_387), .Y(n_473) );
INVx3_ASAP7_75t_L g540 ( .A(n_387), .Y(n_540) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
XOR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_410), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_395), .B(n_400), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .C(n_398), .D(n_399), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .C(n_404), .D(n_408), .Y(n_400) );
INVx1_ASAP7_75t_L g571 ( .A(n_402), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx4_ASAP7_75t_L g441 ( .A(n_407), .Y(n_441) );
INVx4_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
INVx1_ASAP7_75t_L g452 ( .A(n_412), .Y(n_452) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_431), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_417), .C(n_421), .D(n_426), .Y(n_413) );
BUFx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_443), .C(n_447), .Y(n_431) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_440), .B2(n_442), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g458 ( .A(n_454), .Y(n_458) );
INVx1_ASAP7_75t_L g652 ( .A(n_459), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_562), .B2(n_641), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_508), .B2(n_561), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OA22x2_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_490), .B2(n_507), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_479), .Y(n_466) );
NAND4xp25_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .C(n_472), .D(n_474), .Y(n_467) );
BUFx3_ASAP7_75t_L g596 ( .A(n_473), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_477), .B(n_928), .Y(n_927) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g531 ( .A(n_478), .Y(n_531) );
INVx1_ASAP7_75t_L g573 ( .A(n_478), .Y(n_573) );
NAND4xp25_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .C(n_486), .D(n_488), .Y(n_479) );
INVx5_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g515 ( .A(n_482), .Y(n_515) );
INVx1_ASAP7_75t_L g611 ( .A(n_482), .Y(n_611) );
INVx1_ASAP7_75t_L g900 ( .A(n_482), .Y(n_900) );
BUFx4f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g507 ( .A(n_490), .Y(n_507) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_506), .Y(n_490) );
NOR3xp33_ASAP7_75t_SL g506 ( .A(n_491), .B(n_493), .C(n_501), .Y(n_506) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
NAND4xp75_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .C(n_497), .D(n_498), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .C(n_504), .D(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g561 ( .A(n_508), .Y(n_561) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
XNOR2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_541), .Y(n_510) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
NAND4xp25_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .C(n_517), .D(n_520), .Y(n_513) );
BUFx12f_ASAP7_75t_L g583 ( .A(n_518), .Y(n_583) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g581 ( .A(n_522), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_532), .C(n_535), .Y(n_524) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_SL g553 ( .A(n_527), .Y(n_553) );
INVx2_ASAP7_75t_L g892 ( .A(n_527), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_530), .B(n_630), .Y(n_629) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g881 ( .A(n_533), .Y(n_881) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g575 ( .A(n_537), .Y(n_575) );
INVx2_ASAP7_75t_L g884 ( .A(n_537), .Y(n_884) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g559 ( .A(n_538), .Y(n_559) );
INVx2_ASAP7_75t_L g600 ( .A(n_538), .Y(n_600) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g638 ( .A(n_540), .Y(n_638) );
INVx2_ASAP7_75t_L g931 ( .A(n_540), .Y(n_931) );
XNOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_549), .Y(n_543) );
NAND4xp25_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .C(n_547), .D(n_548), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_558), .C(n_560), .Y(n_549) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g577 ( .A(n_552), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_552), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g641 ( .A(n_562), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_586), .B1(n_639), .B2(n_640), .Y(n_562) );
INVx1_ASAP7_75t_L g639 ( .A(n_563), .Y(n_639) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
XNOR2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NOR2xp67_ASAP7_75t_L g567 ( .A(n_568), .B(n_578), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_574), .C(n_576), .Y(n_568) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .C(n_584), .D(n_585), .Y(n_578) );
BUFx4f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
XOR2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_619), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_591), .B(n_602), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .C(n_597), .Y(n_591) );
INVx1_ASAP7_75t_L g617 ( .A(n_592), .Y(n_617) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_595), .Y(n_618) );
INVx1_ASAP7_75t_L g614 ( .A(n_597), .Y(n_614) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_607), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g613 ( .A(n_604), .B(n_614), .C(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_608), .B(n_617), .C(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .C(n_631), .D(n_635), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
OA21x2_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_628), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
BUFx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .C(n_649), .Y(n_644) );
AND2x2_ASAP7_75t_L g908 ( .A(n_645), .B(n_909), .Y(n_908) );
AND2x2_ASAP7_75t_L g935 ( .A(n_645), .B(n_936), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_645), .A2(n_649), .B(n_691), .Y(n_940) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AO21x1_ASAP7_75t_L g938 ( .A1(n_646), .A2(n_939), .B(n_940), .Y(n_938) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g661 ( .A(n_647), .B(n_662), .Y(n_661) );
AND3x4_ASAP7_75t_L g690 ( .A(n_647), .B(n_663), .C(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_648), .B(n_909), .Y(n_936) );
INVx1_ASAP7_75t_L g909 ( .A(n_649), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_873), .B1(n_875), .B2(n_906), .C(n_910), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_833), .C(n_849), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_677), .B(n_780), .C(n_806), .Y(n_655) );
HB1xp67_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_657), .B(n_790), .Y(n_789) );
AOI211xp5_ASAP7_75t_L g806 ( .A1(n_657), .A2(n_807), .B(n_811), .C(n_823), .Y(n_806) );
INVx2_ASAP7_75t_L g834 ( .A(n_657), .Y(n_834) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_658), .Y(n_874) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_659), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
AND2x4_ASAP7_75t_L g671 ( .A(n_661), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g692 ( .A(n_661), .B(n_672), .Y(n_692) );
AND2x2_ASAP7_75t_L g697 ( .A(n_661), .B(n_672), .Y(n_697) );
AND2x4_ASAP7_75t_L g667 ( .A(n_663), .B(n_668), .Y(n_667) );
AND2x4_ASAP7_75t_L g688 ( .A(n_663), .B(n_668), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_663), .B(n_668), .Y(n_723) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g675 ( .A(n_668), .B(n_672), .Y(n_675) );
AND2x2_ASAP7_75t_L g695 ( .A(n_668), .B(n_672), .Y(n_695) );
AND2x2_ASAP7_75t_L g712 ( .A(n_668), .B(n_672), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_673), .B1(n_674), .B2(n_676), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_670), .A2(n_674), .B1(n_719), .B2(n_720), .Y(n_718) );
INVx3_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR4xp25_ASAP7_75t_SL g677 ( .A(n_678), .B(n_734), .C(n_742), .D(n_760), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_698), .A3(n_708), .B1(n_714), .B2(n_727), .C1(n_728), .C2(n_730), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_685), .Y(n_679) );
INVx5_ASAP7_75t_L g735 ( .A(n_680), .Y(n_735) );
INVx3_ASAP7_75t_L g745 ( .A(n_680), .Y(n_745) );
AOI32xp33_ASAP7_75t_L g771 ( .A1(n_680), .A2(n_772), .A3(n_774), .B1(n_776), .B2(n_778), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_680), .B(n_716), .Y(n_822) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g763 ( .A(n_681), .B(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g779 ( .A(n_681), .B(n_686), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_681), .B(n_727), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_681), .B(n_761), .Y(n_840) );
AND2x2_ASAP7_75t_L g867 ( .A(n_681), .B(n_732), .Y(n_867) );
INVx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g731 ( .A(n_682), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g759 ( .A(n_682), .B(n_752), .Y(n_759) );
OR2x2_ASAP7_75t_L g801 ( .A(n_682), .B(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx2_ASAP7_75t_L g802 ( .A(n_685), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_685), .B(n_717), .Y(n_872) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_693), .Y(n_685) );
CKINVDCx6p67_ASAP7_75t_R g727 ( .A(n_686), .Y(n_727) );
INVx1_ASAP7_75t_L g733 ( .A(n_686), .Y(n_733) );
OR2x2_ASAP7_75t_L g752 ( .A(n_686), .B(n_693), .Y(n_752) );
AND2x2_ASAP7_75t_L g815 ( .A(n_686), .B(n_748), .Y(n_815) );
OR2x6_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g748 ( .A(n_693), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_693), .B(n_738), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_693), .B(n_717), .Y(n_777) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_693), .Y(n_785) );
BUFx2_ASAP7_75t_L g791 ( .A(n_693), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_693), .B(n_717), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_693), .B(n_779), .Y(n_843) );
AND2x4_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_707), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_699), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g729 ( .A(n_700), .B(n_708), .Y(n_729) );
AND2x2_ASAP7_75t_L g861 ( .A(n_700), .B(n_740), .Y(n_861) );
AND2x2_ASAP7_75t_L g863 ( .A(n_700), .B(n_864), .Y(n_863) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
OR2x2_ASAP7_75t_L g707 ( .A(n_701), .B(n_704), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_701), .Y(n_726) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
OR2x2_ASAP7_75t_L g725 ( .A(n_704), .B(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_704), .B(n_708), .Y(n_753) );
OR2x2_ASAP7_75t_L g775 ( .A(n_704), .B(n_710), .Y(n_775) );
AND2x2_ASAP7_75t_L g795 ( .A(n_704), .B(n_726), .Y(n_795) );
INVx1_ASAP7_75t_L g810 ( .A(n_704), .Y(n_810) );
AND2x2_ASAP7_75t_L g820 ( .A(n_704), .B(n_794), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_704), .B(n_740), .Y(n_870) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g741 ( .A(n_707), .Y(n_741) );
OR2x2_ASAP7_75t_L g761 ( .A(n_707), .B(n_740), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_707), .B(n_787), .Y(n_786) );
OAI322xp33_ASAP7_75t_L g838 ( .A1(n_707), .A2(n_716), .A3(n_730), .B1(n_747), .B2(n_756), .C1(n_779), .C2(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_707), .B(n_738), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_708), .B(n_715), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_708), .B(n_726), .Y(n_770) );
AND2x2_ASAP7_75t_L g799 ( .A(n_708), .B(n_795), .Y(n_799) );
INVx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g740 ( .A(n_710), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_710), .B(n_738), .Y(n_787) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_725), .Y(n_715) );
INVx1_ASAP7_75t_L g797 ( .A(n_716), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_716), .B(n_790), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_716), .B(n_775), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_716), .B(n_861), .Y(n_860) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_L g738 ( .A(n_717), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_717), .B(n_748), .Y(n_747) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_717), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_717), .B(n_740), .Y(n_826) );
OR2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g757 ( .A(n_725), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_725), .B(n_740), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_725), .B(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_726), .B(n_832), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_726), .A2(n_746), .B1(n_757), .B2(n_815), .C(n_858), .Y(n_857) );
AND2x2_ASAP7_75t_L g790 ( .A(n_727), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g856 ( .A(n_727), .Y(n_856) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_729), .B(n_731), .C(n_797), .Y(n_796) );
OAI21xp5_ASAP7_75t_SL g829 ( .A1(n_729), .A2(n_739), .B(n_830), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_729), .A2(n_739), .B1(n_846), .B2(n_851), .C(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_731), .B(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_732), .B(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
CKINVDCx14_ASAP7_75t_R g859 ( .A(n_735), .Y(n_859) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_L g750 ( .A(n_738), .B(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g805 ( .A(n_738), .B(n_795), .Y(n_805) );
INVx1_ASAP7_75t_SL g854 ( .A(n_738), .Y(n_854) );
AND2x2_ASAP7_75t_L g813 ( .A(n_739), .B(n_797), .Y(n_813) );
AOI211xp5_ASAP7_75t_L g844 ( .A1(n_739), .A2(n_772), .B(n_845), .C(n_848), .Y(n_844) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_740), .B(n_757), .Y(n_756) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_740), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_740), .B(n_805), .Y(n_804) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_749), .B(n_753), .C(n_754), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI311xp33_ASAP7_75t_L g788 ( .A1(n_745), .A2(n_789), .A3(n_792), .B1(n_796), .C1(n_798), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_745), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AOI21xp33_ASAP7_75t_L g841 ( .A1(n_747), .A2(n_769), .B(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g765 ( .A(n_748), .Y(n_765) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_752), .A2(n_753), .B1(n_808), .B2(n_809), .Y(n_807) );
OAI221xp5_ASAP7_75t_L g823 ( .A1(n_752), .A2(n_762), .B1(n_824), .B2(n_827), .C(n_829), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_753), .B(n_872), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_766), .B2(n_769), .C(n_771), .Y(n_760) );
INVx1_ASAP7_75t_L g819 ( .A(n_761), .Y(n_819) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g846 ( .A(n_765), .Y(n_846) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_770), .B(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g848 ( .A(n_772), .B(n_799), .Y(n_848) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g851 ( .A(n_777), .Y(n_851) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_779), .A2(n_834), .B1(n_835), .B2(n_844), .Y(n_833) );
AOI211xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_783), .B(n_788), .C(n_803), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI21xp33_ASAP7_75t_L g803 ( .A1(n_782), .A2(n_802), .B(n_804), .Y(n_803) );
OAI221xp5_ASAP7_75t_L g811 ( .A1(n_782), .A2(n_812), .B1(n_814), .B2(n_816), .C(n_818), .Y(n_811) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_785), .B(n_819), .Y(n_837) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_797), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_797), .B(n_819), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_802), .B(n_822), .Y(n_821) );
OAI221xp5_ASAP7_75t_L g852 ( .A1(n_808), .A2(n_810), .B1(n_853), .B2(n_855), .C(n_857), .Y(n_852) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
AOI211xp5_ASAP7_75t_L g862 ( .A1(n_815), .A2(n_863), .B(n_865), .C(n_871), .Y(n_862) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OAI21xp33_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B(n_821), .Y(n_818) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g864 ( .A(n_826), .Y(n_864) );
INVx1_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
OAI321xp33_ASAP7_75t_L g849 ( .A1(n_834), .A2(n_842), .A3(n_850), .B1(n_859), .B2(n_860), .C(n_862), .Y(n_849) );
NOR4xp25_ASAP7_75t_SL g835 ( .A(n_836), .B(n_838), .C(n_840), .D(n_841), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_854), .B(n_870), .Y(n_869) );
CKINVDCx14_ASAP7_75t_R g855 ( .A(n_856), .Y(n_855) );
INVxp67_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_876), .Y(n_905) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_878), .B(n_896), .Y(n_877) );
NOR3xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_885), .C(n_889), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_879) );
INVxp67_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
OAI21xp33_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_891), .B(n_893), .Y(n_889) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_901), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
NAND2xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx1_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
XNOR2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_933), .Y(n_913) );
NOR3xp33_ASAP7_75t_SL g914 ( .A(n_915), .B(n_919), .C(n_922), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_918), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
NAND4xp25_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .C(n_929), .D(n_932), .Y(n_922) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
endmodule