module fake_jpeg_409_n_39 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_5),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_18),
.B1(n_9),
.B2(n_8),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_10),
.B1(n_9),
.B2(n_7),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_0),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_14),
.C(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_22),
.B(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_13),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_6),
.B1(n_8),
.B2(n_29),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_16),
.Y(n_26)
);

AO221x1_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_8),
.B1(n_21),
.B2(n_0),
.C(n_6),
.Y(n_31)
);

NAND4xp25_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_24),
.C(n_28),
.D(n_33),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_23),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_30),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_30),
.B1(n_32),
.B2(n_25),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_37),
.B(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_36),
.Y(n_39)
);


endmodule