module fake_jpeg_4491_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_66),
.Y(n_94)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_28),
.B1(n_29),
.B2(n_20),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_18),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_73),
.Y(n_117)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_92),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_75),
.A2(n_77),
.B1(n_80),
.B2(n_84),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_28),
.B1(n_33),
.B2(n_19),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_29),
.B1(n_18),
.B2(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_49),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_32),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_18),
.B1(n_25),
.B2(n_34),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_25),
.B1(n_26),
.B2(n_22),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_88),
.B1(n_91),
.B2(n_97),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_49),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_17),
.B(n_32),
.C(n_24),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_33),
.B1(n_21),
.B2(n_23),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_23),
.B1(n_17),
.B2(n_24),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_98),
.B(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_66),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_91)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_55),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_23),
.B1(n_30),
.B2(n_35),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_54),
.B(n_44),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_63),
.A3(n_54),
.B1(n_64),
.B2(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_114),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_64),
.B1(n_63),
.B2(n_35),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_61),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_98),
.C(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_108),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_112),
.B(n_114),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_86),
.Y(n_137)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_115),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_91),
.C(n_95),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_59),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_119),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_31),
.B1(n_35),
.B2(n_17),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_59),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_17),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_99),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_100),
.B(n_119),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_142),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_98),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_17),
.B(n_74),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_136),
.B(n_17),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_137),
.B(n_24),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_123),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_94),
.B1(n_92),
.B2(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_87),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_150),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_39),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_97),
.B1(n_82),
.B2(n_81),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_117),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_107),
.B1(n_116),
.B2(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_155),
.B1(n_156),
.B2(n_73),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_145),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_154),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_104),
.B1(n_108),
.B2(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_104),
.A2(n_74),
.B1(n_82),
.B2(n_81),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_169),
.B(n_185),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_160),
.B(n_165),
.Y(n_199)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_164),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_170),
.B1(n_190),
.B2(n_138),
.Y(n_193)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_101),
.C(n_71),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_171),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_130),
.A2(n_121),
.B(n_111),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_74),
.B1(n_106),
.B2(n_71),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_132),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_177),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_150),
.B(n_152),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_44),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_136),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_178),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_73),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_13),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_13),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_70),
.B(n_106),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_135),
.B(n_96),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_187),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_70),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_138),
.B1(n_135),
.B2(n_151),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_209),
.B1(n_181),
.B2(n_164),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_204),
.B1(n_210),
.B2(n_219),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_203),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_202),
.B(n_32),
.CI(n_35),
.CON(n_237),
.SN(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_180),
.B1(n_173),
.B2(n_160),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_128),
.B1(n_149),
.B2(n_137),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_142),
.B1(n_128),
.B2(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_157),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_134),
.B(n_131),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_32),
.B(n_30),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_158),
.A2(n_143),
.B1(n_157),
.B2(n_129),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_189),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_234),
.B1(n_205),
.B2(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_231),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_188),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_227),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_165),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_208),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_177),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_166),
.B(n_162),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_240),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_168),
.C(n_178),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_243),
.C(n_215),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_235),
.B(n_32),
.Y(n_264)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_167),
.B1(n_157),
.B2(n_96),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_70),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_238),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_237),
.B(n_239),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_129),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_32),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_207),
.C(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_250),
.C(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_207),
.C(n_197),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_216),
.C(n_206),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_236),
.B(n_225),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_193),
.B1(n_204),
.B2(n_199),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_228),
.B1(n_220),
.B2(n_242),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_202),
.C(n_191),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_260),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_201),
.C(n_217),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_221),
.A2(n_195),
.B1(n_31),
.B2(n_30),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_32),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_265),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_235),
.B1(n_237),
.B2(n_229),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_31),
.C(n_1),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_244),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_258),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_272),
.A2(n_275),
.B1(n_279),
.B2(n_281),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_246),
.B(n_226),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_251),
.B1(n_265),
.B2(n_257),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_31),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_282),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_255),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_248),
.A2(n_7),
.B1(n_15),
.B2(n_13),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_267),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_259),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_260),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_288),
.B1(n_294),
.B2(n_282),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_250),
.B1(n_247),
.B2(n_256),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_267),
.C(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_296),
.C(n_9),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_6),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_292),
.C(n_295),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_6),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_0),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_2),
.C(n_3),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_8),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_5),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_281),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_301),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_283),
.B1(n_279),
.B2(n_274),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_303),
.B(n_10),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_8),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_2),
.C(n_3),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_5),
.B(n_10),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_311),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_294),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_SL g321 ( 
.A(n_309),
.B(n_4),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_3),
.C(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_290),
.C(n_10),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_4),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_300),
.B(n_297),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_292),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_320),
.B(n_16),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_309),
.B1(n_306),
.B2(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_325),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_15),
.B(n_16),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_321),
.B(n_316),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_16),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_332),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_R g335 ( 
.A1(n_331),
.A2(n_323),
.B(n_330),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_326),
.Y(n_338)
);


endmodule