module fake_jpeg_27647_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_56),
.B(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_19),
.B1(n_15),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_15),
.B1(n_19),
.B2(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_27),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_20),
.B1(n_16),
.B2(n_32),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_30),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_29),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_22),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_29),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_86),
.B(n_24),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_15),
.B1(n_55),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_100),
.B1(n_70),
.B2(n_68),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_65),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_101),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_59),
.A2(n_25),
.B(n_23),
.C(n_22),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_25),
.B1(n_16),
.B2(n_23),
.Y(n_100)
);

AND2x4_ASAP7_75t_SL g101 ( 
.A(n_61),
.B(n_38),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_39),
.C(n_38),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_58),
.C(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_25),
.B1(n_31),
.B2(n_26),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_23),
.C(n_28),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_110),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_124),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_79),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_109),
.B(n_18),
.Y(n_143)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_114),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_71),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_24),
.C(n_26),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_120),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_21),
.A3(n_22),
.B1(n_10),
.B2(n_11),
.C1(n_14),
.C2(n_12),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_100),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_63),
.C(n_65),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_102),
.C(n_101),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_102),
.B(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_127),
.B(n_137),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_129),
.C(n_130),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_101),
.B(n_92),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_96),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_98),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_141),
.C(n_143),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_94),
.B1(n_90),
.B2(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_118),
.B1(n_105),
.B2(n_113),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_94),
.B(n_84),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_112),
.B(n_85),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_10),
.C(n_2),
.Y(n_156)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_110),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_111),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_116),
.B1(n_88),
.B2(n_16),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_152),
.B1(n_154),
.B2(n_156),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_88),
.C(n_85),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_146),
.C(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_127),
.B1(n_141),
.B2(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_164),
.C(n_167),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_149),
.B1(n_155),
.B2(n_146),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_169),
.B1(n_150),
.B2(n_157),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_130),
.C(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_37),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_133),
.C(n_128),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_125),
.A3(n_91),
.B1(n_74),
.B2(n_78),
.C1(n_77),
.C2(n_18),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_164),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_174),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_0),
.B(n_3),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_172),
.A2(n_173),
.B(n_176),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_156),
.B(n_3),
.Y(n_173)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_0),
.B(n_3),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_168),
.B(n_5),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_6),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_163),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_185),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_162),
.C(n_167),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_173),
.B(n_7),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_7),
.B(n_8),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_17),
.C(n_69),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_189),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_6),
.C(n_7),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_181),
.C(n_182),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_194),
.C(n_9),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_8),
.B(n_9),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_193),
.B(n_38),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_195),
.Y(n_198)
);


endmodule