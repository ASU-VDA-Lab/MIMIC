module real_aes_8667_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g510 ( .A1(n_0), .A2(n_153), .B(n_511), .C(n_512), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_1), .B(n_172), .Y(n_514) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_90), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_3), .A2(n_139), .B(n_144), .C(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_4), .A2(n_134), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_5), .B(n_209), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_6), .A2(n_134), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_7), .B(n_172), .Y(n_238) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_8), .A2(n_157), .B(n_465), .Y(n_464) );
AND2x6_ASAP7_75t_L g139 ( .A(n_9), .B(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_10), .A2(n_139), .B(n_144), .C(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g151 ( .A(n_11), .Y(n_151) );
INVx1_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_12), .B(n_42), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_13), .B(n_149), .Y(n_186) );
INVx1_ASAP7_75t_L g132 ( .A(n_14), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_15), .B(n_209), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_16), .A2(n_152), .B(n_166), .C(n_170), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_17), .B(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_18), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_19), .B(n_278), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_20), .A2(n_196), .B(n_197), .C(n_199), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_21), .A2(n_144), .B(n_213), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_22), .B(n_149), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_23), .B(n_149), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_24), .Y(n_220) );
INVx1_ASAP7_75t_L g208 ( .A(n_25), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_26), .A2(n_144), .B(n_213), .C(n_468), .Y(n_467) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_27), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_28), .Y(n_179) );
INVx1_ASAP7_75t_L g274 ( .A(n_29), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_30), .A2(n_134), .B(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_31), .A2(n_102), .B1(n_111), .B2(n_751), .Y(n_101) );
INVx2_ASAP7_75t_L g137 ( .A(n_32), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_33), .A2(n_225), .B(n_446), .C(n_480), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_34), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_35), .A2(n_196), .B(n_234), .C(n_236), .Y(n_233) );
INVxp67_ASAP7_75t_L g275 ( .A(n_36), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_37), .B(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_38), .A2(n_144), .B(n_207), .C(n_213), .Y(n_206) );
CKINVDCx14_ASAP7_75t_R g232 ( .A(n_39), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_40), .A2(n_47), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_40), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_41), .A2(n_46), .B1(n_725), .B2(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_41), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_42), .B(n_106), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_43), .A2(n_148), .B(n_150), .C(n_153), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_44), .B(n_269), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_45), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_46), .Y(n_725) );
INVx1_ASAP7_75t_L g742 ( .A(n_47), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_48), .B(n_209), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_49), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_50), .B(n_134), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_51), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_52), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_53), .A2(n_225), .B(n_446), .C(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g513 ( .A(n_54), .Y(n_513) );
INVx1_ASAP7_75t_L g448 ( .A(n_55), .Y(n_448) );
INVx1_ASAP7_75t_L g194 ( .A(n_56), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_57), .B(n_134), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_58), .Y(n_494) );
CKINVDCx14_ASAP7_75t_R g142 ( .A(n_59), .Y(n_142) );
INVx1_ASAP7_75t_L g140 ( .A(n_60), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_61), .B(n_134), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_62), .B(n_172), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_63), .A2(n_212), .B(n_459), .C(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g131 ( .A(n_64), .Y(n_131) );
INVx1_ASAP7_75t_SL g235 ( .A(n_65), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_66), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_67), .B(n_209), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_68), .B(n_172), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_69), .B(n_152), .Y(n_523) );
INVx1_ASAP7_75t_L g223 ( .A(n_70), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_71), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_72), .B(n_185), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_73), .A2(n_144), .B(n_225), .C(n_499), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_74), .Y(n_457) );
INVx1_ASAP7_75t_L g110 ( .A(n_75), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_76), .A2(n_134), .B(n_141), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_77), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_78), .A2(n_134), .B(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_79), .A2(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g164 ( .A(n_80), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_81), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_82), .B(n_184), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_83), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_84), .A2(n_134), .B(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g167 ( .A(n_85), .Y(n_167) );
INVx2_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx1_ASAP7_75t_L g183 ( .A(n_87), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_88), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_89), .B(n_149), .Y(n_524) );
INVx2_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
OR2x2_ASAP7_75t_L g437 ( .A(n_90), .B(n_119), .Y(n_437) );
OR2x2_ASAP7_75t_L g744 ( .A(n_90), .B(n_732), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_91), .A2(n_144), .B(n_222), .C(n_225), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_92), .B(n_134), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_93), .Y(n_481) );
INVxp67_ASAP7_75t_L g461 ( .A(n_94), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_95), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g198 ( .A(n_97), .Y(n_198) );
INVx1_ASAP7_75t_L g500 ( .A(n_98), .Y(n_500) );
INVx1_ASAP7_75t_L g520 ( .A(n_99), .Y(n_520) );
AND2x2_ASAP7_75t_L g451 ( .A(n_100), .B(n_128), .Y(n_451) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_103), .Y(n_752) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO221x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_734), .B1(n_737), .B2(n_745), .C(n_747), .Y(n_111) );
OAI222xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_723), .B1(n_724), .B2(n_727), .C1(n_730), .C2(n_733), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_122), .B1(n_434), .B2(n_438), .Y(n_113) );
AOI22x1_ASAP7_75t_SL g727 ( .A1(n_114), .A2(n_434), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_118), .B(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_119), .Y(n_732) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
INVx2_ASAP7_75t_L g728 ( .A(n_122), .Y(n_728) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_364), .Y(n_122) );
NAND5xp2_ASAP7_75t_L g123 ( .A(n_124), .B(n_279), .C(n_311), .D(n_328), .E(n_351), .Y(n_123) );
AOI221xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_202), .B1(n_239), .B2(n_243), .C(n_247), .Y(n_124) );
INVx1_ASAP7_75t_L g391 ( .A(n_125), .Y(n_391) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_174), .Y(n_125) );
AND3x2_ASAP7_75t_L g366 ( .A(n_126), .B(n_176), .C(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_159), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_127), .B(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g254 ( .A(n_127), .Y(n_254) );
AND2x2_ASAP7_75t_L g258 ( .A(n_127), .B(n_190), .Y(n_258) );
INVx2_ASAP7_75t_L g288 ( .A(n_127), .Y(n_288) );
OR2x2_ASAP7_75t_L g299 ( .A(n_127), .B(n_191), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_127), .B(n_175), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_127), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g378 ( .A(n_127), .B(n_191), .Y(n_378) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_133), .B(n_156), .Y(n_127) );
INVx1_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_128), .A2(n_180), .B(n_205), .C(n_206), .Y(n_204) );
INVx2_ASAP7_75t_L g228 ( .A(n_128), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_128), .A2(n_444), .B(n_445), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_128), .A2(n_478), .B(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_L g158 ( .A(n_129), .B(n_130), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
BUFx2_ASAP7_75t_L g269 ( .A(n_134), .Y(n_269) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_139), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_135), .B(n_139), .Y(n_180) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g212 ( .A(n_136), .Y(n_212) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
INVx1_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
INVx1_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_138), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_138), .Y(n_152) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
INVx1_ASAP7_75t_L g470 ( .A(n_138), .Y(n_470) );
INVx4_ASAP7_75t_SL g155 ( .A(n_139), .Y(n_155) );
BUFx3_ASAP7_75t_L g213 ( .A(n_139), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_SL g141 ( .A1(n_142), .A2(n_143), .B(n_147), .C(n_155), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_SL g163 ( .A1(n_143), .A2(n_155), .B(n_164), .C(n_165), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_SL g193 ( .A1(n_143), .A2(n_155), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_143), .A2(n_155), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_143), .A2(n_155), .B(n_271), .C(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g446 ( .A(n_143), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_143), .A2(n_155), .B(n_457), .C(n_458), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_SL g508 ( .A1(n_143), .A2(n_155), .B(n_509), .C(n_510), .Y(n_508) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx3_ASAP7_75t_L g154 ( .A(n_145), .Y(n_154) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_145), .Y(n_237) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g196 ( .A(n_149), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx5_ASAP7_75t_L g209 ( .A(n_152), .Y(n_209) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_154), .Y(n_450) );
INVx1_ASAP7_75t_L g225 ( .A(n_155), .Y(n_225) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_157), .Y(n_161) );
INVx4_ASAP7_75t_L g173 ( .A(n_157), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_157), .A2(n_466), .B(n_467), .Y(n_465) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g266 ( .A(n_158), .Y(n_266) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_159), .Y(n_257) );
AND2x2_ASAP7_75t_L g319 ( .A(n_159), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_159), .B(n_175), .Y(n_338) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g246 ( .A(n_160), .B(n_175), .Y(n_246) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_160), .Y(n_253) );
AND2x2_ASAP7_75t_L g305 ( .A(n_160), .B(n_191), .Y(n_305) );
NAND3xp33_ASAP7_75t_L g330 ( .A(n_160), .B(n_174), .C(n_288), .Y(n_330) );
AND2x2_ASAP7_75t_L g395 ( .A(n_160), .B(n_176), .Y(n_395) );
AND2x2_ASAP7_75t_L g429 ( .A(n_160), .B(n_175), .Y(n_429) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_171), .Y(n_160) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_161), .A2(n_192), .B(n_201), .Y(n_191) );
OA21x2_ASAP7_75t_L g229 ( .A1(n_161), .A2(n_230), .B(n_238), .Y(n_229) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_161), .A2(n_455), .B(n_462), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_168), .B(n_198), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_168), .A2(n_209), .B1(n_274), .B2(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g459 ( .A(n_168), .Y(n_459) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_172), .A2(n_507), .B(n_514), .Y(n_506) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_173), .B(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_173), .B(n_215), .Y(n_214) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_173), .A2(n_219), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_173), .B(n_484), .Y(n_483) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_173), .A2(n_497), .B(n_504), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_173), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_173), .A2(n_519), .B(n_525), .Y(n_518) );
INVxp67_ASAP7_75t_L g255 ( .A(n_174), .Y(n_255) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_190), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_175), .B(n_288), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_175), .B(n_319), .Y(n_327) );
AND2x2_ASAP7_75t_L g377 ( .A(n_175), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g405 ( .A(n_175), .Y(n_405) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g312 ( .A(n_176), .B(n_305), .Y(n_312) );
BUFx3_ASAP7_75t_L g344 ( .A(n_176), .Y(n_344) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_188), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_177), .B(n_494), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_180), .A2(n_220), .B(n_221), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_180), .A2(n_520), .B(n_521), .Y(n_519) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_187), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_184), .A2(n_187), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_184), .A2(n_448), .B(n_449), .C(n_450), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_184), .A2(n_450), .B(n_481), .C(n_482), .Y(n_480) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g320 ( .A(n_190), .Y(n_320) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_191), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_196), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_196), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g472 ( .A(n_199), .Y(n_472) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_202), .A2(n_380), .B1(n_382), .B2(n_383), .Y(n_379) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_216), .Y(n_202) );
AND2x2_ASAP7_75t_L g239 ( .A(n_203), .B(n_240), .Y(n_239) );
INVx3_ASAP7_75t_SL g250 ( .A(n_203), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_203), .B(n_283), .Y(n_315) );
OR2x2_ASAP7_75t_L g334 ( .A(n_203), .B(n_217), .Y(n_334) );
AND2x2_ASAP7_75t_L g339 ( .A(n_203), .B(n_291), .Y(n_339) );
AND2x2_ASAP7_75t_L g342 ( .A(n_203), .B(n_284), .Y(n_342) );
AND2x2_ASAP7_75t_L g354 ( .A(n_203), .B(n_229), .Y(n_354) );
AND2x2_ASAP7_75t_L g370 ( .A(n_203), .B(n_218), .Y(n_370) );
AND2x4_ASAP7_75t_L g373 ( .A(n_203), .B(n_241), .Y(n_373) );
OR2x2_ASAP7_75t_L g390 ( .A(n_203), .B(n_326), .Y(n_390) );
OR2x2_ASAP7_75t_L g421 ( .A(n_203), .B(n_263), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_203), .B(n_349), .Y(n_423) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .C(n_211), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_209), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g511 ( .A(n_209), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_211), .A2(n_491), .B(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_212), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g297 ( .A(n_216), .B(n_261), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_216), .B(n_284), .Y(n_416) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_229), .Y(n_216) );
AND2x2_ASAP7_75t_L g249 ( .A(n_217), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g283 ( .A(n_217), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g291 ( .A(n_217), .B(n_263), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_217), .B(n_241), .Y(n_309) );
OR2x2_ASAP7_75t_L g326 ( .A(n_217), .B(n_284), .Y(n_326) );
INVx2_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g242 ( .A(n_218), .Y(n_242) );
AND2x2_ASAP7_75t_L g349 ( .A(n_218), .B(n_229), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
INVx2_ASAP7_75t_L g241 ( .A(n_229), .Y(n_241) );
INVx1_ASAP7_75t_L g361 ( .A(n_229), .Y(n_361) );
AND2x2_ASAP7_75t_L g411 ( .A(n_229), .B(n_250), .Y(n_411) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_237), .Y(n_502) );
AND2x2_ASAP7_75t_L g260 ( .A(n_240), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g295 ( .A(n_240), .B(n_250), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_240), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
AND2x2_ASAP7_75t_L g282 ( .A(n_241), .B(n_250), .Y(n_282) );
OR2x2_ASAP7_75t_L g398 ( .A(n_242), .B(n_372), .Y(n_398) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_245), .B(n_378), .Y(n_384) );
INVx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OAI32xp33_ASAP7_75t_L g340 ( .A1(n_246), .A2(n_341), .A3(n_343), .B1(n_345), .B2(n_346), .Y(n_340) );
OR2x2_ASAP7_75t_L g357 ( .A(n_246), .B(n_299), .Y(n_357) );
OAI21xp33_ASAP7_75t_SL g382 ( .A1(n_246), .A2(n_256), .B(n_287), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_251), .B1(n_256), .B2(n_259), .Y(n_247) );
INVxp33_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_249), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_250), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g308 ( .A(n_250), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g408 ( .A(n_250), .B(n_349), .Y(n_408) );
OR2x2_ASAP7_75t_L g432 ( .A(n_250), .B(n_326), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g415 ( .A1(n_251), .A2(n_314), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g292 ( .A(n_253), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_253), .B(n_258), .Y(n_310) );
AND2x2_ASAP7_75t_L g332 ( .A(n_254), .B(n_305), .Y(n_332) );
INVx1_ASAP7_75t_L g345 ( .A(n_254), .Y(n_345) );
OR2x2_ASAP7_75t_L g350 ( .A(n_254), .B(n_284), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_257), .B(n_299), .Y(n_298) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_258), .A2(n_281), .B1(n_286), .B2(n_290), .Y(n_280) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_261), .A2(n_323), .B1(n_330), .B2(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g407 ( .A(n_261), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_263), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g426 ( .A(n_263), .B(n_309), .Y(n_426) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .B(n_276), .Y(n_263) );
INVx1_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_266), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_268), .A2(n_277), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI21xp5_ASAP7_75t_SL g487 ( .A1(n_278), .A2(n_488), .B(n_489), .Y(n_487) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_292), .B1(n_293), .B2(n_298), .C(n_300), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_282), .B(n_284), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_282), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g301 ( .A(n_283), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_283), .A2(n_389), .B(n_390), .C(n_391), .Y(n_388) );
AND2x2_ASAP7_75t_L g393 ( .A(n_283), .B(n_373), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_SL g431 ( .A1(n_283), .A2(n_372), .B(n_432), .C(n_433), .Y(n_431) );
BUFx3_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_287), .B(n_344), .Y(n_387) );
AOI211xp5_ASAP7_75t_L g406 ( .A1(n_287), .A2(n_407), .B(n_409), .C(n_415), .Y(n_406) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVxp67_ASAP7_75t_L g367 ( .A(n_289), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_291), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AOI211xp5_ASAP7_75t_L g311 ( .A1(n_295), .A2(n_312), .B(n_313), .C(n_321), .Y(n_311) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g396 ( .A(n_299), .Y(n_396) );
OR2x2_ASAP7_75t_L g413 ( .A(n_299), .B(n_343), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_302), .B1(n_307), .B2(n_310), .Y(n_300) );
OAI22xp33_ASAP7_75t_L g313 ( .A1(n_302), .A2(n_314), .B1(n_315), .B2(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
OR2x2_ASAP7_75t_L g400 ( .A(n_304), .B(n_344), .Y(n_400) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g355 ( .A(n_305), .B(n_345), .Y(n_355) );
INVx1_ASAP7_75t_L g363 ( .A(n_306), .Y(n_363) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_309), .B(n_323), .Y(n_371) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_319), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g428 ( .A(n_320), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B(n_327), .Y(n_321) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_323), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_323), .B(n_354), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_323), .B(n_349), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_323), .B(n_370), .Y(n_381) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_323), .A2(n_333), .B(n_373), .C(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AOI221xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_333), .B1(n_335), .B2(n_339), .C(n_340), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_337), .B(n_345), .Y(n_419) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g430 ( .A1(n_339), .A2(n_354), .B(n_356), .C(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_342), .B(n_349), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_343), .B(n_396), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_344), .Y(n_343) );
INVxp33_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AOI21xp33_ASAP7_75t_SL g359 ( .A1(n_348), .A2(n_360), .B(n_362), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_348), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_349), .B(n_403), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_356), .B2(n_358), .C(n_359), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_355), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g389 ( .A(n_361), .Y(n_389) );
NAND5xp2_ASAP7_75t_L g364 ( .A(n_365), .B(n_392), .C(n_406), .D(n_417), .E(n_430), .Y(n_364) );
AOI211xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B(n_375), .C(n_388), .Y(n_365) );
INVx2_ASAP7_75t_SL g412 ( .A(n_366), .Y(n_412) );
NAND4xp25_ASAP7_75t_SL g368 ( .A(n_369), .B(n_371), .C(n_372), .D(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI211xp5_ASAP7_75t_SL g375 ( .A1(n_374), .A2(n_376), .B(n_379), .C(n_385), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_377), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_377), .A2(n_418), .B1(n_420), .B2(n_422), .C(n_424), .Y(n_417) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI221xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_394), .B1(n_397), .B2(n_399), .C(n_401), .Y(n_392) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_400), .A2(n_423), .B1(n_425), .B2(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_413), .B2(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx4_ASAP7_75t_L g729 ( .A(n_438), .Y(n_729) );
XOR2xp5_ASAP7_75t_L g739 ( .A(n_438), .B(n_740), .Y(n_739) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR5x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_596), .C(n_674), .D(n_698), .E(n_715), .Y(n_439) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_473), .B(n_515), .C(n_573), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_452), .Y(n_441) );
AND2x2_ASAP7_75t_L g527 ( .A(n_442), .B(n_454), .Y(n_527) );
INVx5_ASAP7_75t_SL g555 ( .A(n_442), .Y(n_555) );
AND2x2_ASAP7_75t_L g591 ( .A(n_442), .B(n_576), .Y(n_591) );
OR2x2_ASAP7_75t_L g630 ( .A(n_442), .B(n_453), .Y(n_630) );
OR2x2_ASAP7_75t_L g661 ( .A(n_442), .B(n_552), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_442), .B(n_565), .Y(n_697) );
AND2x2_ASAP7_75t_L g709 ( .A(n_442), .B(n_552), .Y(n_709) );
OR2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_451), .Y(n_442) );
AND2x2_ASAP7_75t_L g708 ( .A(n_452), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g571 ( .A(n_453), .B(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_454), .B(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_454), .Y(n_564) );
INVx3_ASAP7_75t_L g579 ( .A(n_454), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_454), .B(n_463), .Y(n_603) );
OR2x2_ASAP7_75t_L g612 ( .A(n_454), .B(n_555), .Y(n_612) );
AND2x2_ASAP7_75t_L g616 ( .A(n_454), .B(n_576), .Y(n_616) );
AND2x2_ASAP7_75t_L g622 ( .A(n_454), .B(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_L g659 ( .A(n_454), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_454), .B(n_518), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_459), .A2(n_500), .B(n_501), .C(n_502), .Y(n_499) );
OR2x2_ASAP7_75t_L g565 ( .A(n_463), .B(n_518), .Y(n_565) );
AND2x2_ASAP7_75t_L g576 ( .A(n_463), .B(n_552), .Y(n_576) );
AND2x2_ASAP7_75t_L g588 ( .A(n_463), .B(n_579), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_463), .B(n_518), .Y(n_611) );
INVx1_ASAP7_75t_SL g623 ( .A(n_463), .Y(n_623) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g517 ( .A(n_464), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_464), .B(n_555), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B(n_472), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_472), .A2(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .Y(n_474) );
AND2x2_ASAP7_75t_L g536 ( .A(n_475), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_475), .B(n_495), .Y(n_540) );
AND2x2_ASAP7_75t_L g543 ( .A(n_475), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_475), .B(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g568 ( .A(n_475), .B(n_559), .Y(n_568) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_475), .Y(n_587) );
AND2x2_ASAP7_75t_L g608 ( .A(n_475), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g618 ( .A(n_475), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g664 ( .A(n_475), .B(n_547), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_475), .B(n_570), .Y(n_691) );
INVx5_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g561 ( .A(n_476), .Y(n_561) );
AND2x2_ASAP7_75t_L g627 ( .A(n_476), .B(n_559), .Y(n_627) );
AND2x2_ASAP7_75t_L g711 ( .A(n_476), .B(n_579), .Y(n_711) );
OR2x6_ASAP7_75t_L g476 ( .A(n_477), .B(n_483), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_485), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g700 ( .A(n_485), .Y(n_700) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
AND2x2_ASAP7_75t_L g530 ( .A(n_486), .B(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g539 ( .A(n_486), .B(n_537), .Y(n_539) );
INVx5_ASAP7_75t_L g547 ( .A(n_486), .Y(n_547) );
AND2x2_ASAP7_75t_L g570 ( .A(n_486), .B(n_506), .Y(n_570) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_486), .Y(n_607) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_L g648 ( .A(n_495), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_495), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g681 ( .A(n_495), .B(n_547), .Y(n_681) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_495), .A2(n_604), .B(n_711), .C(n_712), .Y(n_710) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
BUFx2_ASAP7_75t_L g531 ( .A(n_496), .Y(n_531) );
INVx2_ASAP7_75t_L g535 ( .A(n_496), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_503), .Y(n_497) );
INVx2_ASAP7_75t_L g537 ( .A(n_506), .Y(n_537) );
AND2x2_ASAP7_75t_L g544 ( .A(n_506), .B(n_535), .Y(n_544) );
AND2x2_ASAP7_75t_L g635 ( .A(n_506), .B(n_547), .Y(n_635) );
AOI211x1_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_528), .B(n_541), .C(n_566), .Y(n_515) );
INVx1_ASAP7_75t_L g632 ( .A(n_516), .Y(n_632) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
INVx5_ASAP7_75t_SL g552 ( .A(n_518), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_518), .B(n_622), .Y(n_621) );
AOI311xp33_ASAP7_75t_L g640 ( .A1(n_518), .A2(n_641), .A3(n_643), .B(n_644), .C(n_650), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g675 ( .A1(n_518), .A2(n_588), .B(n_676), .C(n_679), .Y(n_675) );
INVxp67_ASAP7_75t_L g595 ( .A(n_527), .Y(n_595) );
NAND4xp25_ASAP7_75t_SL g528 ( .A(n_529), .B(n_532), .C(n_538), .D(n_540), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_529), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g586 ( .A(n_530), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_533), .B(n_539), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_533), .B(n_546), .Y(n_666) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_534), .B(n_547), .Y(n_684) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g559 ( .A(n_535), .Y(n_559) );
INVxp67_ASAP7_75t_L g594 ( .A(n_536), .Y(n_594) );
AND2x4_ASAP7_75t_L g546 ( .A(n_537), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g620 ( .A(n_537), .B(n_559), .Y(n_620) );
INVx1_ASAP7_75t_L g647 ( .A(n_537), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_537), .B(n_634), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_538), .B(n_608), .Y(n_628) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_539), .B(n_561), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_539), .B(n_608), .Y(n_707) );
INVx1_ASAP7_75t_L g718 ( .A(n_540), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .B(n_548), .C(n_556), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g560 ( .A(n_544), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g598 ( .A(n_544), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g580 ( .A(n_545), .Y(n_580) );
AND2x2_ASAP7_75t_L g557 ( .A(n_546), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_546), .B(n_608), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_546), .B(n_627), .Y(n_651) );
OR2x2_ASAP7_75t_L g567 ( .A(n_547), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g599 ( .A(n_547), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_547), .B(n_559), .Y(n_614) );
AND2x2_ASAP7_75t_L g671 ( .A(n_547), .B(n_627), .Y(n_671) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_547), .Y(n_678) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_549), .A2(n_561), .B1(n_683), .B2(n_685), .C(n_688), .Y(n_682) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g572 ( .A(n_552), .B(n_555), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_552), .B(n_622), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_552), .B(n_579), .Y(n_687) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g672 ( .A(n_554), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g686 ( .A(n_554), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_555), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g583 ( .A(n_555), .B(n_576), .Y(n_583) );
AND2x2_ASAP7_75t_L g653 ( .A(n_555), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_555), .B(n_602), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_555), .B(n_703), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_560), .B(n_562), .Y(n_556) );
INVx2_ASAP7_75t_L g589 ( .A(n_557), .Y(n_589) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g609 ( .A(n_559), .Y(n_609) );
OR2x2_ASAP7_75t_L g613 ( .A(n_561), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g716 ( .A(n_561), .B(n_684), .Y(n_716) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AOI21xp33_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_569), .B(n_571), .Y(n_566) );
INVx1_ASAP7_75t_L g720 ( .A(n_567), .Y(n_720) );
INVx2_ASAP7_75t_SL g634 ( .A(n_568), .Y(n_634) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_571), .A2(n_652), .B(n_716), .C(n_717), .Y(n_715) );
OAI322xp33_ASAP7_75t_SL g584 ( .A1(n_572), .A2(n_585), .A3(n_588), .B1(n_589), .B2(n_590), .C1(n_592), .C2(n_595), .Y(n_584) );
INVx2_ASAP7_75t_L g604 ( .A(n_572), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_580), .B1(n_581), .B2(n_583), .C(n_584), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp33_ASAP7_75t_SL g650 ( .A1(n_575), .A2(n_651), .B1(n_652), .B2(n_655), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_576), .B(n_579), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_576), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g649 ( .A(n_578), .B(n_611), .Y(n_649) );
INVx1_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_583), .A2(n_693), .B(n_695), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g617 ( .A1(n_585), .A2(n_618), .B(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp67_ASAP7_75t_SL g646 ( .A(n_587), .B(n_647), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_587), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g703 ( .A(n_588), .Y(n_703) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_624), .C(n_640), .D(n_656), .Y(n_596) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_605), .C(n_617), .Y(n_597) );
INVx1_ASAP7_75t_L g689 ( .A(n_598), .Y(n_689) );
AND2x2_ASAP7_75t_L g637 ( .A(n_599), .B(n_620), .Y(n_637) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_604), .B(n_639), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_610), .B1(n_613), .B2(n_615), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_607), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g655 ( .A(n_608), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_608), .A2(n_647), .B(n_670), .C(n_672), .Y(n_669) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g654 ( .A(n_611), .Y(n_654) );
INVx1_ASAP7_75t_L g714 ( .A(n_612), .Y(n_714) );
NAND2xp33_ASAP7_75t_SL g704 ( .A(n_613), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g643 ( .A(n_622), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_628), .B(n_629), .C(n_631), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_636), .B2(n_638), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_634), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_639), .B(n_660), .Y(n_722) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI21xp33_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_648), .B(n_649), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_662), .B1(n_665), .B2(n_667), .C(n_669), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_672), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_688) );
NAND3xp33_ASAP7_75t_SL g674 ( .A(n_675), .B(n_682), .C(n_692), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_701), .C(n_710), .Y(n_698) );
INVx1_ASAP7_75t_L g719 ( .A(n_699), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_706), .B2(n_708), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
BUFx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g746 ( .A(n_736), .Y(n_746) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
BUFx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g750 ( .A(n_744), .Y(n_750) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
endmodule