module fake_jpeg_22977_n_240 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_240);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_17),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_33),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_40),
.B1(n_38),
.B2(n_34),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_65),
.B1(n_40),
.B2(n_36),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_38),
.B(n_36),
.C(n_18),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_60),
.A2(n_75),
.B(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_40),
.B1(n_21),
.B2(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_34),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_84),
.C(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_77),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_76),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_41),
.C(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_35),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_89),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_88),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_18),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_18),
.B(n_23),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_18),
.C(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_82),
.B1(n_92),
.B2(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_100),
.B1(n_111),
.B2(n_82),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_36),
.B1(n_23),
.B2(n_53),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_36),
.B1(n_51),
.B2(n_21),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_112),
.B1(n_115),
.B2(n_118),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_33),
.B(n_24),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_116),
.B(n_73),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_21),
.B1(n_33),
.B2(n_24),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_24),
.B1(n_26),
.B2(n_25),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_19),
.B(n_31),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_62),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_118)
);

OAI211xp5_ASAP7_75t_L g119 ( 
.A1(n_62),
.A2(n_32),
.B(n_29),
.C(n_22),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_63),
.B1(n_19),
.B2(n_20),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_62),
.A2(n_26),
.B1(n_29),
.B2(n_22),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_20),
.B1(n_89),
.B2(n_87),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_141),
.B1(n_146),
.B2(n_95),
.Y(n_166)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_124),
.Y(n_150)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_130),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_66),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_138),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_147),
.B1(n_111),
.B2(n_110),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_93),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_86),
.B1(n_85),
.B2(n_78),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_145),
.B(n_148),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_73),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_78),
.B1(n_77),
.B2(n_26),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_0),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_129),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_138),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_158),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_102),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_163),
.C(n_168),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_100),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_134),
.B(n_133),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_164),
.B(n_27),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_106),
.C(n_103),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_149),
.B(n_164),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_101),
.C(n_99),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_95),
.B(n_100),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_81),
.C(n_70),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_70),
.C(n_27),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_142),
.C(n_140),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_137),
.A3(n_147),
.B1(n_132),
.B2(n_128),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_180),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_168),
.C(n_157),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_139),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_123),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_188),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g197 ( 
.A(n_187),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_124),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_165),
.C(n_160),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_199),
.C(n_200),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_171),
.B1(n_167),
.B2(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_181),
.C(n_187),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_156),
.C(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_204),
.C(n_183),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_170),
.C(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_182),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_208),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_169),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_176),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_177),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_191),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_174),
.B1(n_178),
.B2(n_173),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_197),
.B1(n_201),
.B2(n_194),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_223),
.C(n_214),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_175),
.B(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_215),
.B(n_205),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_124),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_6),
.B(n_7),
.Y(n_227)
);

OAI322xp33_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_220),
.A2(n_4),
.B(n_5),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_227),
.B(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_226),
.B(n_228),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_10),
.C(n_12),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_221),
.B(n_216),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_231),
.A2(n_219),
.B(n_221),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_SL g235 ( 
.A1(n_233),
.A2(n_217),
.B(n_14),
.C(n_15),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_235),
.B(n_236),
.CI(n_16),
.CON(n_238),
.SN(n_238)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_16),
.B1(n_12),
.B2(n_14),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_230),
.C(n_238),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_16),
.Y(n_240)
);


endmodule