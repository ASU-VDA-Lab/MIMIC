module real_jpeg_31982_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_0),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_0),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g399 ( 
.A(n_0),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_1),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_1),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_1),
.B(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_1),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_1),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_1),
.B(n_260),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_1),
.B(n_481),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_3),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_4),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_4),
.B(n_121),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_4),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_4),
.B(n_142),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_4),
.B(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_4),
.B(n_260),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_49),
.Y(n_48)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_5),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_5),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_126),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_5),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_5),
.B(n_171),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_5),
.B(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_6),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_6),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_6),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_6),
.B(n_180),
.Y(n_179)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_6),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_6),
.B(n_474),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_7),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_9),
.Y(n_402)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_10),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_L g91 ( 
.A(n_11),
.B(n_92),
.Y(n_91)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_11),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_11),
.B(n_158),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_11),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_11),
.B(n_365),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_11),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_11),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_12),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_12),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_12),
.B(n_86),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_12),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_12),
.B(n_74),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_12),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_12),
.B(n_422),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_21),
.B(n_491),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_13),
.B(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_14),
.B(n_40),
.Y(n_100)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

NAND2x1_ASAP7_75t_SL g225 ( 
.A(n_14),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_14),
.B(n_478),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_40),
.Y(n_39)
);

NAND2x1_ASAP7_75t_L g170 ( 
.A(n_16),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_16),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_16),
.B(n_458),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_17),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_43),
.Y(n_42)
);

NAND2x1_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_18),
.B(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_18),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_18),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_18),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_18),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_18),
.B(n_397),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_35),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_19),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_19),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_19),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_19),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_19),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_446),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_284),
.B(n_443),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_235),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_25),
.A2(n_444),
.B(n_445),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_189),
.Y(n_25)
);

NOR2xp67_ASAP7_75t_L g445 ( 
.A(n_26),
.B(n_189),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_112),
.C(n_167),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_28),
.B(n_167),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_76),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_46),
.C(n_65),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_30),
.B(n_46),
.C(n_65),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_30),
.A2(n_31),
.B1(n_46),
.B2(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2x1_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_42),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_34),
.B(n_38),
.C(n_42),
.Y(n_176)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_37),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_38),
.A2(n_39),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_39),
.B(n_170),
.C(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_45),
.Y(n_482)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_57),
.B(n_63),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_50),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_53),
.B(n_64),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_56),
.Y(n_223)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_56),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_56),
.Y(n_465)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_57),
.Y(n_276)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_62),
.Y(n_458)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_65),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_73),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_70),
.C(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_72),
.Y(n_232)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_89),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_77),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_78),
.B(n_85),
.C(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_80),
.Y(n_205)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_85),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_85),
.B(n_200),
.C(n_202),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_86),
.Y(n_210)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_89),
.B(n_191),
.C(n_192),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_101),
.B(n_111),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_99),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_SL g164 ( 
.A(n_91),
.B(n_95),
.C(n_99),
.Y(n_164)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_98),
.Y(n_350)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_98),
.Y(n_378)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_107),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_107),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_107),
.Y(n_165)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_106),
.Y(n_274)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_106),
.Y(n_371)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_112),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_137),
.C(n_160),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_113),
.B(n_239),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_131),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_115),
.B(n_117),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_118),
.A2(n_119),
.B1(n_131),
.B2(n_132),
.Y(n_311)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_123),
.B(n_127),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_120),
.B(n_250),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_128),
.B(n_130),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_123),
.A2(n_124),
.B1(n_130),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_129),
.B(n_186),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_130),
.Y(n_251)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OA21x2_ASAP7_75t_SL g295 ( 
.A1(n_132),
.A2(n_133),
.B(n_136),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_138),
.A2(n_161),
.B1(n_162),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_138),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_151),
.C(n_156),
.Y(n_138)
);

XOR2x1_ASAP7_75t_L g280 ( 
.A(n_139),
.B(n_281),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.C(n_150),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_140),
.A2(n_141),
.B1(n_150),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_143),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_145),
.B(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g475 ( 
.A(n_159),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_176),
.C(n_177),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_172),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_172),
.B(n_209),
.C(n_212),
.Y(n_467)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_181),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_188),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_190),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_206),
.B2(n_234),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_R g487 ( 
.A(n_194),
.B(n_206),
.C(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_196),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_198),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_SL g449 ( 
.A(n_204),
.B(n_450),
.C(n_452),
.Y(n_449)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

XNOR2x2_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_208),
.B(n_218),
.C(n_219),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_212),
.A2(n_213),
.B1(n_457),
.B2(n_459),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_220),
.B(n_225),
.C(n_229),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_229),
.B1(n_230),
.B2(n_233),
.Y(n_224)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_282),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_236),
.B(n_282),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.C(n_246),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_238),
.B(n_242),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_246),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_275),
.C(n_278),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_247),
.A2(n_248),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_263),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_249),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_252),
.A2(n_263),
.B1(n_264),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_252),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_253),
.A2(n_254),
.B1(n_258),
.B2(n_259),
.Y(n_332)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_262),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_262),
.Y(n_424)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.C(n_271),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_265),
.A2(n_266),
.B1(n_271),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_270),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_279),
.B1(n_280),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_339),
.B(n_441),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_312),
.B(n_315),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_286),
.B(n_312),
.C(n_442),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_308),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_309),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.C(n_296),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_295),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_296),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.C(n_304),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_355),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_345)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_355)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_337),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_316),
.B(n_337),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.C(n_333),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_334),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.C(n_332),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_332),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.C(n_328),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_328),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_325),
.B(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_331),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_358),
.B(n_440),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_356),
.Y(n_340)
);

NAND2xp33_ASAP7_75t_SL g440 ( 
.A(n_341),
.B(n_356),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.C(n_354),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_342),
.B(n_438),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_344),
.B(n_354),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.C(n_347),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_346),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

AO22x1_ASAP7_75t_L g380 ( 
.A1(n_348),
.A2(n_349),
.B1(n_351),
.B2(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_435),
.B(n_439),
.Y(n_358)
);

OAI21x1_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_392),
.B(n_434),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_381),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_361),
.B(n_381),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_374),
.C(n_380),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_362),
.A2(n_363),
.B1(n_430),
.B2(n_432),
.Y(n_429)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_368),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_387),
.C(n_388),
.Y(n_386)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_372),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_374),
.A2(n_375),
.B1(n_380),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_379),
.Y(n_410)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_380),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_385),
.B2(n_391),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_386),
.C(n_389),
.Y(n_436)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_385),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_427),
.B(n_433),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_411),
.B(n_426),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_403),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_395),
.B(n_403),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_400),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_400),
.Y(n_419)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx8_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_400),
.B(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_410),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_407),
.B2(n_409),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_405),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_409),
.C(n_410),
.Y(n_428)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_420),
.B(n_425),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_419),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_419),
.Y(n_425)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_436),
.B(n_437),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_489),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_487),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_SL g490 ( 
.A(n_448),
.B(n_487),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_453),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_469),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_466),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_460),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_457),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_486),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_470)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_471),
.Y(n_485)
);

XNOR2x1_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_480),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_476),
.B1(n_477),
.B2(n_479),
.Y(n_472)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_473),
.Y(n_479)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);


endmodule