module fake_jpeg_8308_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_40),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_40),
.C(n_37),
.Y(n_68)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_53),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_32),
.B1(n_27),
.B2(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_32),
.B1(n_27),
.B2(n_40),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_35),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_37),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_76),
.B(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_62),
.B(n_72),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_69),
.B1(n_24),
.B2(n_34),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_40),
.B1(n_36),
.B2(n_32),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_67),
.A2(n_84),
.B1(n_47),
.B2(n_57),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_70),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_27),
.B1(n_32),
.B2(n_16),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_35),
.B(n_37),
.C(n_36),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_33),
.B(n_17),
.C(n_16),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_36),
.B1(n_17),
.B2(n_24),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_34),
.B1(n_47),
.B2(n_46),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_22),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_94),
.B1(n_107),
.B2(n_79),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_109),
.B1(n_80),
.B2(n_86),
.Y(n_118)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_90),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_30),
.B(n_22),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_93),
.B(n_97),
.Y(n_140)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_98),
.B(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_29),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_68),
.B(n_19),
.CI(n_39),
.CON(n_102),
.SN(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_31),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_70),
.B1(n_34),
.B2(n_65),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_152)
);

INVx6_ASAP7_75t_SL g116 ( 
.A(n_92),
.Y(n_116)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_117),
.B(n_125),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_28),
.B(n_26),
.Y(n_161)
);

AOI22x1_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_39),
.B1(n_85),
.B2(n_21),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_86),
.B1(n_65),
.B2(n_79),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_130),
.B1(n_133),
.B2(n_82),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_63),
.B1(n_22),
.B2(n_30),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_132),
.B1(n_126),
.B2(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_75),
.B1(n_63),
.B2(n_30),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_39),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_135),
.C(n_82),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_20),
.B1(n_25),
.B2(n_31),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_26),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_97),
.B1(n_109),
.B2(n_103),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_149),
.B1(n_154),
.B2(n_159),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_148),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_135),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_151),
.C(n_129),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_55),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_71),
.B1(n_25),
.B2(n_20),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_165),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_55),
.B(n_52),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_158),
.B(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_194)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_160),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_0),
.Y(n_158)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_39),
.B1(n_26),
.B2(n_23),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_52),
.B(n_23),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_43),
.B1(n_23),
.B2(n_21),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_9),
.Y(n_168)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_182),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_113),
.B1(n_128),
.B2(n_127),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_194),
.B1(n_162),
.B2(n_165),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_185),
.C(n_188),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_186),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_119),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_190),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_130),
.C(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_133),
.Y(n_187)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_81),
.C(n_23),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_193),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_21),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_152),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_198),
.C(n_201),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_192),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_158),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_193),
.B1(n_186),
.B2(n_191),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_202),
.A2(n_207),
.B1(n_210),
.B2(n_212),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_158),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_188),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_167),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_208),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_155),
.B1(n_150),
.B2(n_149),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_168),
.B(n_154),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_179),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_144),
.B1(n_166),
.B2(n_81),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_218),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_187),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_206),
.C(n_205),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_221),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_194),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_177),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_225),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_177),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_181),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_175),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_234),
.B(n_237),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_215),
.B1(n_214),
.B2(n_195),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_240),
.B1(n_243),
.B2(n_218),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_219),
.A2(n_204),
.B(n_209),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_183),
.B1(n_208),
.B2(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_7),
.B(n_3),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_211),
.B1(n_208),
.B2(n_3),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_221),
.B1(n_220),
.B2(n_217),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_8),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_250),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_239),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_255),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_238),
.C(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_254),
.C(n_12),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_11),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_12),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_11),
.C(n_4),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_11),
.B(n_4),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_244),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_258),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_233),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_253),
.B1(n_246),
.B2(n_13),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_248),
.B(n_12),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_0),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_265),
.C(n_15),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_260),
.B(n_263),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_13),
.B(n_14),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_257),
.B(n_15),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_271),
.Y(n_275)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_273),
.B(n_15),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_0),
.C(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_268),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_256),
.Y(n_279)
);


endmodule