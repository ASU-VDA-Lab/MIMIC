module fake_jpeg_2602_n_202 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_45),
.B(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_72),
.A2(n_65),
.B1(n_52),
.B2(n_57),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_87),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_54),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_60),
.B1(n_65),
.B2(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_52),
.B1(n_60),
.B2(n_63),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_55),
.B(n_54),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_101),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_67),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_62),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_64),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_59),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_47),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_6),
.C(n_7),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_78),
.B1(n_90),
.B2(n_49),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_129),
.B(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_83),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_66),
.B(n_53),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_150),
.B(n_9),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_93),
.B(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_122),
.B(n_117),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_96),
.B(n_101),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_146),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_103),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_134),
.C(n_135),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_99),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_50),
.B1(n_107),
.B2(n_90),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_139),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_50),
.C(n_39),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_151),
.C(n_117),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_20),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_156),
.B(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_158),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_22),
.B(n_37),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_7),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_17),
.C(n_36),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_149),
.B(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_166),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_140),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_11),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_133),
.A2(n_11),
.B(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_12),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_29),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_13),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_176),
.Y(n_186)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_147),
.B1(n_152),
.B2(n_16),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_162),
.B1(n_155),
.B2(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_178),
.B(n_159),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_171),
.C(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_187),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_162),
.B(n_167),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_182),
.B(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_181),
.C(n_180),
.Y(n_190)
);

OAI321xp33_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_160),
.A3(n_16),
.B1(n_15),
.B2(n_27),
.C(n_25),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_185),
.C(n_186),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_172),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_33),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_191),
.Y(n_199)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_197),
.B(n_198),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_34),
.Y(n_202)
);


endmodule