module fake_jpeg_14610_n_98 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_22),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_0),
.B1(n_3),
.B2(n_7),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_53),
.B(n_59),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_3),
.B1(n_11),
.B2(n_14),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_46),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_66),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_57),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_23),
.B1(n_29),
.B2(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_67),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_36),
.B(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_34),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_83),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_52),
.B1(n_49),
.B2(n_66),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_45),
.B1(n_28),
.B2(n_37),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_77),
.B1(n_63),
.B2(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_74),
.Y(n_88)
);

XNOR2x1_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_70),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_74),
.C(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_85),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_89),
.B(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_93),
.B(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.C(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_73),
.B1(n_43),
.B2(n_60),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_62),
.Y(n_98)
);


endmodule