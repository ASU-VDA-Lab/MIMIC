module fake_jpeg_9032_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_32),
.Y(n_58)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_29),
.B1(n_33),
.B2(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_38),
.B1(n_29),
.B2(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_46),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_53),
.B1(n_61),
.B2(n_16),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_16),
.B1(n_27),
.B2(n_18),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_63),
.A2(n_49),
.B1(n_34),
.B2(n_18),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_70),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_81),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_23),
.B1(n_30),
.B2(n_20),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_85),
.C(n_62),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_116),
.B(n_22),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_48),
.B1(n_56),
.B2(n_44),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_104),
.B1(n_105),
.B2(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_53),
.B1(n_48),
.B2(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_113),
.A2(n_69),
.B1(n_84),
.B2(n_81),
.Y(n_119)
);

MAJx3_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_34),
.C(n_42),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_24),
.B(n_31),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_25),
.B1(n_20),
.B2(n_26),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_55),
.C(n_24),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_122),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_24),
.B1(n_25),
.B2(n_76),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_82),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_136),
.B(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_123),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_125),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_115),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_87),
.B1(n_68),
.B2(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_137),
.B(n_138),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_142),
.B1(n_64),
.B2(n_25),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_26),
.B1(n_31),
.B2(n_18),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_97),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_26),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_86),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_93),
.B(n_114),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_154),
.B(n_160),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_114),
.B(n_116),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_98),
.B1(n_100),
.B2(n_94),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_159),
.B1(n_172),
.B2(n_142),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_144),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_100),
.B1(n_76),
.B2(n_92),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_164),
.B1(n_168),
.B2(n_125),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_100),
.B1(n_89),
.B2(n_112),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_106),
.B1(n_112),
.B2(n_102),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_102),
.B1(n_106),
.B2(n_90),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_24),
.CI(n_88),
.CON(n_165),
.SN(n_165)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_165),
.B(n_144),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_90),
.B1(n_97),
.B2(n_64),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_64),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_174),
.C(n_177),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_126),
.B(n_132),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_22),
.C(n_1),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_22),
.C(n_1),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_22),
.A3(n_8),
.B1(n_9),
.B2(n_15),
.Y(n_178)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_182),
.B(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_191),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_192),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_143),
.B(n_137),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_196),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_136),
.B1(n_131),
.B2(n_139),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_140),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_202),
.Y(n_214)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_199),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_122),
.B1(n_121),
.B2(n_141),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_198),
.B1(n_178),
.B2(n_151),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_148),
.A2(n_8),
.B(n_12),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_0),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_6),
.Y(n_202)
);

OR2x4_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_22),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_165),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_156),
.B(n_6),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_205),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_12),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_158),
.C(n_152),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_211),
.C(n_216),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_173),
.B1(n_169),
.B2(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_153),
.C(n_162),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_163),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_165),
.C(n_169),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_170),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_229),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_151),
.B1(n_168),
.B2(n_166),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_200),
.B1(n_190),
.B2(n_201),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_190),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_204),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_239),
.C(n_211),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_215),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_247),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_227),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_206),
.B1(n_201),
.B2(n_9),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_221),
.B1(n_220),
.B2(n_226),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_0),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_216),
.C(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_217),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_258),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_252),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_229),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_254),
.C(n_252),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_208),
.C(n_242),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_228),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_257),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_214),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_243),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_244),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_270),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_266),
.B1(n_262),
.B2(n_271),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_256),
.A2(n_245),
.B(n_233),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_241),
.C(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_269),
.C(n_9),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_232),
.B(n_243),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_246),
.C(n_231),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_235),
.B(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_234),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_263),
.B1(n_269),
.B2(n_248),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_278),
.B1(n_284),
.B2(n_3),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_226),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_281),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_214),
.B1(n_3),
.B2(n_4),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_10),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_10),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_284)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_12),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.C(n_284),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_282),
.A2(n_10),
.B(n_11),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_278),
.B(n_11),
.CI(n_3),
.CON(n_289),
.SN(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_283),
.C(n_280),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_286),
.B(n_290),
.C(n_279),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_297),
.A2(n_290),
.B(n_293),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_296),
.B(n_275),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_295),
.B(n_289),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_5),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_5),
.B(n_286),
.Y(n_302)
);


endmodule