module fake_ibex_1726_n_1612 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_9, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_211, n_218, n_314, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1612);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_9;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1612;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_1326;
wire n_971;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1558;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_422;
wire n_1609;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_1577;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1540;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_650;
wire n_409;
wire n_1575;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1460;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_1607;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_193),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_27),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_43),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_82),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_9),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_291),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_133),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_302),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_185),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_21),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_2),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_106),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_112),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_87),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_32),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_161),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_257),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_219),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_183),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_75),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_56),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_55),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_296),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_43),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_45),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_204),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_131),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_118),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_238),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_223),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_325),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_123),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_196),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_242),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_94),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_234),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_122),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_21),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_292),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_37),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_119),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_198),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_289),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_12),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_1),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_111),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_311),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_126),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_174),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_244),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_287),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_304),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_269),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_249),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_170),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_139),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_282),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_176),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_252),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_25),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_300),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_166),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_317),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_84),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_310),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_136),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_201),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_35),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_50),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_264),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_284),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_182),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_150),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_305),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_159),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_327),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_277),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_326),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_306),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_10),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_298),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_65),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_149),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_35),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_77),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_259),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_73),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_299),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_281),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_260),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_7),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_106),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_162),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_107),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_233),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_266),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_216),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_301),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_308),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_128),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_76),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_123),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_297),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_239),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_218),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_138),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_221),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_276),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_2),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_68),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_28),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_267),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_19),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_271),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_199),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_61),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_120),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_274),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_17),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_137),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_255),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_235),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_253),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_1),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_226),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_144),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_236),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_273),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_208),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_39),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_246),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_141),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_225),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_323),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_275),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_184),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_82),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_261),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_270),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_142),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_102),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_157),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_124),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_206),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_102),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_130),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_247),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_313),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_316),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_288),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_293),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_171),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_286),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_77),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_280),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_272),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_319),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_85),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_214),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_19),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_27),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_94),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_228),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_107),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_40),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_314),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_303),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_44),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_30),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_11),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_165),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_232),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_135),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_104),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_5),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_265),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_8),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_168),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_122),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_140),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_52),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_179),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_258),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_207),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_187),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_322),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_262),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_101),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_101),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_241),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_307),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_70),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_98),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_321),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_42),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_86),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_209),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_210),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_256),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_312),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_57),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_117),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_294),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_156),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_15),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_279),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_126),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_268),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_158),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_290),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_181),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_120),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_240),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_180),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_33),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_263),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_63),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_190),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_315),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_213),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_251),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_295),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_3),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_145),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_254),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_188),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_100),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_117),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_11),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_116),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_0),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_99),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_248),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_250),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_278),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_32),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_5),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_186),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_97),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_55),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_91),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_84),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_283),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_81),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_59),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_227),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_344),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_384),
.B(n_0),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_339),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_371),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_339),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_553),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_349),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_344),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_540),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_381),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_569),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_569),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_333),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_386),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_333),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_355),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_404),
.B(n_3),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_422),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_425),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_442),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_439),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_442),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_355),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_407),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_509),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_493),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_555),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_573),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_573),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_475),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_345),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_529),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_532),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_366),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_414),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_434),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_398),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_330),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_340),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_409),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_342),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_343),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_350),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_493),
.Y(n_624)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_523),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_358),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_567),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_351),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_500),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_500),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_369),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_450),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_380),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_502),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_329),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_450),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_401),
.Y(n_637)
);

INVxp33_ASAP7_75t_SL g638 ( 
.A(n_352),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_502),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_416),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_424),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_426),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_452),
.B(n_4),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_433),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_480),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_480),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_524),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_537),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_504),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_407),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_559),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_561),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_568),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_572),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_504),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_390),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_390),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_574),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_520),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_520),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_535),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_582),
.Y(n_663)
);

CKINVDCx16_ASAP7_75t_R g664 ( 
.A(n_625),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_585),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_662),
.B(n_510),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_584),
.B(n_512),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_587),
.B(n_412),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_611),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_588),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_614),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_628),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_592),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_596),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_610),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_615),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_635),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_581),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_651),
.B(n_349),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_583),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_597),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_638),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_585),
.Y(n_683)
);

BUFx8_ASAP7_75t_L g684 ( 
.A(n_616),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_599),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_590),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_591),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_589),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_612),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_657),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_619),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_621),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_613),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_593),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_606),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_598),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_R g698 ( 
.A(n_638),
.B(n_354),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_623),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_618),
.B(n_412),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_600),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_632),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_636),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_658),
.B(n_362),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_645),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_647),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_626),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_631),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_601),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_633),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_617),
.B(n_329),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_604),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_579),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_637),
.B(n_370),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_640),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_605),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_650),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_642),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_607),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_606),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_656),
.Y(n_721)
);

OA21x2_ASAP7_75t_L g722 ( 
.A1(n_641),
.A2(n_464),
.B(n_405),
.Y(n_722)
);

CKINVDCx6p67_ASAP7_75t_R g723 ( 
.A(n_579),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_620),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_624),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_608),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_627),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_624),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_609),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_644),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_646),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_648),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_629),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_629),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_649),
.B(n_652),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_654),
.B(n_329),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_653),
.B(n_412),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_655),
.B(n_405),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_659),
.B(n_372),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_630),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_580),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_595),
.B(n_331),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_643),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_586),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_586),
.B(n_535),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_630),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_594),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_602),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_602),
.B(n_376),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_634),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_634),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_661),
.B(n_378),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_639),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_639),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_660),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_660),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_661),
.B(n_464),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_638),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_657),
.B(n_328),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_611),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_585),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_611),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_628),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_638),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_606),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_585),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_582),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_611),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_635),
.B(n_535),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_662),
.B(n_467),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_611),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_606),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_611),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_SL g776 ( 
.A(n_635),
.B(n_554),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_R g778 ( 
.A(n_638),
.B(n_392),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_611),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_606),
.Y(n_780)
);

OA21x2_ASAP7_75t_L g781 ( 
.A1(n_585),
.A2(n_538),
.B(n_467),
.Y(n_781)
);

AND2x6_ASAP7_75t_L g782 ( 
.A(n_662),
.B(n_479),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_603),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_662),
.B(n_396),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_628),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_635),
.B(n_554),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_662),
.B(n_400),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_582),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_SL g789 ( 
.A1(n_606),
.A2(n_534),
.B1(n_377),
.B2(n_448),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_SL g790 ( 
.A1(n_606),
.A2(n_534),
.B1(n_445),
.B2(n_417),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_603),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_611),
.Y(n_792)
);

OA21x2_ASAP7_75t_L g793 ( 
.A1(n_585),
.A2(n_551),
.B(n_538),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_603),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_603),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_582),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_611),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_582),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_603),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_611),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_611),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_675),
.B(n_554),
.Y(n_802)
);

BUFx4f_ASAP7_75t_L g803 ( 
.A(n_770),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_722),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_682),
.Y(n_805)
);

INVx5_ASAP7_75t_L g806 ( 
.A(n_762),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_722),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_722),
.Y(n_808)
);

AND2x6_ASAP7_75t_L g809 ( 
.A(n_786),
.B(n_479),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_799),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_737),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_668),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_715),
.B(n_335),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_759),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_682),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_737),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_675),
.B(n_741),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_715),
.B(n_336),
.Y(n_818)
);

BUFx10_ASAP7_75t_L g819 ( 
.A(n_677),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_718),
.B(n_337),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_718),
.B(n_558),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_736),
.A2(n_419),
.B1(n_441),
.B2(n_423),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_743),
.B(n_341),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_668),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_688),
.B(n_797),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_765),
.B(n_443),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_700),
.A2(n_412),
.B1(n_334),
.B2(n_338),
.Y(n_827)
);

AND2x6_ASAP7_75t_L g828 ( 
.A(n_711),
.B(n_700),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_672),
.B(n_449),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_801),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_764),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_785),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_687),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_669),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_799),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_691),
.B(n_347),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_800),
.Y(n_837)
);

AND2x6_ASAP7_75t_L g838 ( 
.A(n_745),
.B(n_332),
.Y(n_838)
);

INVx8_ASAP7_75t_L g839 ( 
.A(n_782),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_692),
.B(n_348),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_671),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_677),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_776),
.B(n_451),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_753),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_690),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_694),
.B(n_353),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_704),
.B(n_558),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_676),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_687),
.Y(n_849)
);

NAND2x1p5_ASAP7_75t_L g850 ( 
.A(n_713),
.B(n_373),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_690),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_687),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_687),
.Y(n_853)
);

AND2x6_ASAP7_75t_L g854 ( 
.A(n_772),
.B(n_356),
.Y(n_854)
);

AND2x6_ASAP7_75t_L g855 ( 
.A(n_772),
.B(n_359),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_784),
.B(n_357),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_695),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_761),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_724),
.B(n_456),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_742),
.A2(n_469),
.B1(n_473),
.B2(n_462),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_763),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_753),
.Y(n_862)
);

AND2x6_ASAP7_75t_L g863 ( 
.A(n_699),
.B(n_363),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_787),
.B(n_361),
.Y(n_864)
);

AND3x2_ASAP7_75t_L g865 ( 
.A(n_724),
.B(n_368),
.C(n_364),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_663),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_695),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_769),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_735),
.B(n_477),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_707),
.B(n_365),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_783),
.Y(n_871)
);

NOR2x1p5_ASAP7_75t_L g872 ( 
.A(n_723),
.B(n_486),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_730),
.B(n_708),
.Y(n_873)
);

AND2x2_ASAP7_75t_SL g874 ( 
.A(n_664),
.B(n_382),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_710),
.B(n_367),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_771),
.B(n_492),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_727),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_714),
.B(n_374),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_773),
.B(n_775),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_791),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_794),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_731),
.B(n_494),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_795),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_744),
.B(n_383),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_746),
.B(n_385),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_732),
.B(n_739),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_781),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_667),
.B(n_375),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_666),
.B(n_379),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_709),
.B(n_387),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_684),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_777),
.B(n_388),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_695),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_695),
.Y(n_894)
);

BUFx10_ASAP7_75t_L g895 ( 
.A(n_758),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_709),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_L g897 ( 
.A1(n_779),
.A2(n_497),
.B(n_496),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_SL g898 ( 
.A1(n_696),
.A2(n_506),
.B1(n_507),
.B2(n_501),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_665),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_665),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_792),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_686),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_684),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_782),
.B(n_394),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_697),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_696),
.Y(n_906)
);

AND2x6_ASAP7_75t_L g907 ( 
.A(n_678),
.B(n_389),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_680),
.B(n_395),
.Y(n_908)
);

NOR2x1p5_ASAP7_75t_L g909 ( 
.A(n_670),
.B(n_511),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_701),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_782),
.B(n_712),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_758),
.B(n_513),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_738),
.B(n_528),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_767),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_701),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_782),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_750),
.B(n_360),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_698),
.B(n_525),
.C(n_521),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_701),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_716),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_748),
.B(n_539),
.Y(n_921)
);

CKINVDCx16_ASAP7_75t_R g922 ( 
.A(n_698),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_673),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_719),
.B(n_527),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_781),
.Y(n_925)
);

AND2x6_ASAP7_75t_L g926 ( 
.A(n_683),
.B(n_397),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_738),
.B(n_533),
.Y(n_927)
);

XOR2xp5_ASAP7_75t_L g928 ( 
.A(n_720),
.B(n_544),
.Y(n_928)
);

AND3x4_ASAP7_75t_L g929 ( 
.A(n_789),
.B(n_551),
.C(n_549),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_702),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_726),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_729),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_679),
.B(n_547),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_679),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_703),
.B(n_399),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_705),
.B(n_560),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_778),
.A2(n_563),
.B1(n_564),
.B2(n_562),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_749),
.A2(n_576),
.B1(n_577),
.B2(n_571),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_781),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_760),
.B(n_391),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_793),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_793),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_793),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_706),
.B(n_406),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_778),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_717),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_721),
.B(n_393),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_674),
.B(n_457),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_681),
.B(n_685),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_689),
.B(n_402),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_752),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_693),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_754),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_768),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_788),
.B(n_796),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_798),
.B(n_415),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_728),
.B(n_418),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_733),
.B(n_403),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_734),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_790),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_740),
.B(n_550),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_751),
.Y(n_962)
);

INVxp33_ASAP7_75t_L g963 ( 
.A(n_755),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_756),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_757),
.Y(n_965)
);

INVxp67_ASAP7_75t_SL g966 ( 
.A(n_780),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_720),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_725),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_725),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_747),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_747),
.B(n_408),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_766),
.B(n_410),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_766),
.B(n_420),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_774),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_774),
.A2(n_431),
.B1(n_440),
.B2(n_427),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_682),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_677),
.B(n_4),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_668),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_715),
.B(n_411),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_799),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_718),
.B(n_413),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_677),
.B(n_6),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_668),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_668),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_675),
.B(n_454),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_799),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_718),
.B(n_421),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_799),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_715),
.B(n_428),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_675),
.B(n_429),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_668),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_668),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_799),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_715),
.B(n_430),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_668),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_668),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_715),
.B(n_432),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_682),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_668),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_770),
.B(n_461),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_759),
.B(n_578),
.Y(n_1001)
);

BUFx4f_ASAP7_75t_L g1002 ( 
.A(n_770),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_759),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_799),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_668),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_668),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_675),
.B(n_487),
.C(n_478),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_759),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_675),
.B(n_435),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_675),
.B(n_437),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_759),
.B(n_488),
.Y(n_1011)
);

AND2x6_ASAP7_75t_L g1012 ( 
.A(n_770),
.B(n_499),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_815),
.B(n_438),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_814),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_832),
.B(n_6),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_998),
.A2(n_976),
.B1(n_1008),
.B2(n_1003),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_985),
.B(n_444),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_830),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_805),
.B(n_447),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_834),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_851),
.B(n_7),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_876),
.A2(n_515),
.B1(n_516),
.B2(n_508),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_SL g1023 ( 
.A(n_916),
.B(n_453),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_985),
.B(n_455),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_825),
.B(n_458),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_819),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_825),
.A2(n_556),
.B1(n_557),
.B2(n_542),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_831),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_916),
.B(n_459),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_869),
.B(n_460),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_886),
.A2(n_570),
.B1(n_465),
.B2(n_468),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_837),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_879),
.B(n_463),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_819),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_841),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_879),
.B(n_471),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_842),
.B(n_472),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_845),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_803),
.B(n_474),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_829),
.B(n_8),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_873),
.B(n_924),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_803),
.B(n_476),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_876),
.A2(n_482),
.B1(n_483),
.B2(n_481),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_927),
.B(n_484),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1011),
.B(n_575),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_839),
.B(n_485),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_927),
.B(n_489),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_874),
.A2(n_495),
.B1(n_498),
.B2(n_491),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_1002),
.B(n_503),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_859),
.B(n_9),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1002),
.B(n_505),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_848),
.B(n_514),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_850),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_858),
.B(n_517),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_861),
.B(n_518),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_813),
.B(n_522),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_826),
.B(n_526),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_868),
.A2(n_436),
.B(n_446),
.C(n_346),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_804),
.A2(n_531),
.B(n_530),
.Y(n_1059)
);

CKINVDCx11_ASAP7_75t_R g1060 ( 
.A(n_891),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_968),
.B(n_10),
.Y(n_1061)
);

NOR2x2_ASAP7_75t_L g1062 ( 
.A(n_960),
.B(n_13),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_818),
.B(n_566),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_979),
.B(n_989),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_901),
.B(n_536),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_994),
.B(n_997),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_921),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_933),
.B(n_541),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_839),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_804),
.A2(n_545),
.B(n_543),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_933),
.B(n_546),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_932),
.B(n_548),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_817),
.B(n_13),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_827),
.B(n_436),
.C(n_346),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_953),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_810),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_945),
.B(n_552),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_871),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_882),
.B(n_565),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1001),
.B(n_346),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_896),
.B(n_14),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_854),
.B(n_16),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_854),
.B(n_17),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_807),
.A2(n_446),
.B(n_436),
.Y(n_1084)
);

AND2x6_ASAP7_75t_SL g1085 ( 
.A(n_949),
.B(n_18),
.Y(n_1085)
);

NAND3xp33_ASAP7_75t_L g1086 ( 
.A(n_1007),
.B(n_466),
.C(n_446),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_854),
.A2(n_470),
.B1(n_519),
.B2(n_466),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_930),
.B(n_18),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_855),
.B(n_20),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_912),
.A2(n_470),
.B1(n_466),
.B2(n_519),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_L g1091 ( 
.A(n_863),
.B(n_466),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_880),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_855),
.B(n_20),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_855),
.B(n_22),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_903),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_810),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_812),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_967),
.B(n_23),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_977),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_824),
.Y(n_1100)
);

NOR2x2_ASAP7_75t_L g1101 ( 
.A(n_884),
.B(n_885),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_881),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_902),
.A2(n_519),
.B(n_470),
.C(n_25),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_810),
.B(n_470),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_835),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_981),
.B(n_23),
.Y(n_1106)
);

NAND2x1_ASAP7_75t_L g1107 ( 
.A(n_833),
.B(n_519),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_895),
.B(n_24),
.Y(n_1108)
);

BUFx5_ASAP7_75t_L g1109 ( 
.A(n_887),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1000),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_835),
.B(n_26),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_953),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_835),
.B(n_29),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_988),
.B(n_31),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_895),
.B(n_33),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_956),
.B(n_34),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_987),
.B(n_34),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_955),
.B(n_36),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_883),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_899),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_913),
.B(n_36),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_936),
.B(n_877),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_978),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_947),
.B(n_37),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_913),
.B(n_38),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_821),
.B(n_38),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_988),
.B(n_39),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_956),
.B(n_40),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_822),
.B(n_41),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_928),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_988),
.B(n_41),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1000),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_944),
.B(n_46),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_843),
.B(n_46),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_966),
.B(n_47),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_838),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_983),
.Y(n_1137)
);

AO22x1_ASAP7_75t_L g1138 ( 
.A1(n_929),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_809),
.B(n_51),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_925),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_809),
.B(n_51),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_838),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_948),
.B(n_53),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_809),
.B(n_54),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_900),
.B(n_56),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_944),
.B(n_57),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_809),
.B(n_58),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_820),
.B(n_58),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_905),
.B(n_59),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_951),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_984),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_860),
.B(n_60),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_991),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_884),
.B(n_63),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_807),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_920),
.B(n_64),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1000),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_838),
.A2(n_70),
.B1(n_67),
.B2(n_69),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_823),
.B(n_69),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_808),
.A2(n_132),
.B(n_129),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_931),
.B(n_71),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_802),
.B(n_72),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_849),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_828),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_969),
.B(n_74),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_925),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_992),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_890),
.B(n_78),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_863),
.B(n_78),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_995),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_925),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_917),
.B(n_79),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_836),
.B(n_79),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_840),
.B(n_846),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_863),
.B(n_80),
.Y(n_1175)
);

AO22x1_ASAP7_75t_L g1176 ( 
.A1(n_866),
.A2(n_83),
.B1(n_80),
.B2(n_81),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_863),
.B(n_907),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_857),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_914),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_808),
.B(n_134),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1000),
.A2(n_86),
.B1(n_83),
.B2(n_85),
.Y(n_1181)
);

NOR2xp67_ASAP7_75t_L g1182 ( 
.A(n_962),
.B(n_87),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_973),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_969),
.B(n_88),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_870),
.B(n_88),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_923),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1012),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_907),
.B(n_89),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_887),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_907),
.B(n_92),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_907),
.B(n_93),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1069),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1041),
.B(n_1012),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1014),
.B(n_922),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1014),
.B(n_1012),
.Y(n_1195)
);

INVx8_ASAP7_75t_L g1196 ( 
.A(n_1073),
.Y(n_1196)
);

BUFx8_ASAP7_75t_SL g1197 ( 
.A(n_1186),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1018),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1060),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1020),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1095),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1032),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1028),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1067),
.B(n_963),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1069),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1026),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1067),
.A2(n_973),
.B1(n_1012),
.B2(n_957),
.Y(n_1207)
);

NOR3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1129),
.B(n_954),
.C(n_862),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1034),
.Y(n_1209)
);

NOR3xp33_ASAP7_75t_L g1210 ( 
.A(n_1138),
.B(n_964),
.C(n_959),
.Y(n_1210)
);

NOR3xp33_ASAP7_75t_SL g1211 ( 
.A(n_1154),
.B(n_844),
.C(n_898),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1099),
.B(n_970),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1038),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1122),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1073),
.A2(n_973),
.B1(n_957),
.B2(n_828),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1145),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1035),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1016),
.B(n_828),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1050),
.B(n_828),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1118),
.B(n_909),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1140),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_R g1222 ( 
.A(n_1046),
.B(n_906),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1084),
.A2(n_942),
.B(n_941),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1023),
.B(n_946),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1097),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1100),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1099),
.B(n_982),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_SL g1228 ( 
.A(n_1053),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1123),
.Y(n_1229)
);

XNOR2xp5_ASAP7_75t_L g1230 ( 
.A(n_1130),
.B(n_872),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1140),
.Y(n_1231)
);

INVx6_ASAP7_75t_L g1232 ( 
.A(n_1085),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1152),
.B(n_970),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1137),
.Y(n_1234)
);

INVx4_ASAP7_75t_L g1235 ( 
.A(n_1145),
.Y(n_1235)
);

INVx5_ASAP7_75t_L g1236 ( 
.A(n_1076),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1015),
.B(n_937),
.Y(n_1237)
);

OR2x4_ASAP7_75t_L g1238 ( 
.A(n_1101),
.B(n_974),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1183),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1151),
.Y(n_1240)
);

NOR3xp33_ASAP7_75t_L g1241 ( 
.A(n_1108),
.B(n_959),
.C(n_952),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1037),
.A2(n_973),
.B1(n_972),
.B2(n_965),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1062),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1140),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1023),
.B(n_918),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1153),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1167),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1076),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_R g1249 ( 
.A(n_1046),
.B(n_865),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1166),
.Y(n_1250)
);

BUFx4f_ASAP7_75t_L g1251 ( 
.A(n_1162),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1166),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1096),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1040),
.B(n_847),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1043),
.B(n_904),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1162),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1109),
.B(n_938),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1120),
.B(n_885),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_1088),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1166),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1170),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1048),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1165),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1146),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1184),
.Y(n_1265)
);

OR2x6_ASAP7_75t_SL g1266 ( 
.A(n_1098),
.B(n_875),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1022),
.B(n_975),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_R g1268 ( 
.A(n_1091),
.B(n_961),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1171),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1013),
.B(n_911),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1116),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1149),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1124),
.B(n_996),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_1171),
.B(n_943),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1156),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_L g1276 ( 
.A(n_1172),
.B(n_940),
.C(n_971),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1161),
.Y(n_1277)
);

CKINVDCx6p67_ASAP7_75t_R g1278 ( 
.A(n_1135),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_SL g1279 ( 
.A(n_1177),
.B(n_990),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1078),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1121),
.Y(n_1281)
);

OR2x6_ASAP7_75t_L g1282 ( 
.A(n_1176),
.B(n_1182),
.Y(n_1282)
);

NOR3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1128),
.B(n_958),
.C(n_935),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1179),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1096),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1105),
.Y(n_1286)
);

NAND2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1045),
.B(n_1105),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1171),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1092),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1143),
.B(n_878),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1102),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1061),
.Y(n_1292)
);

BUFx4f_ASAP7_75t_L g1293 ( 
.A(n_1119),
.Y(n_1293)
);

NOR3xp33_ASAP7_75t_SL g1294 ( 
.A(n_1133),
.B(n_950),
.C(n_897),
.Y(n_1294)
);

BUFx10_ASAP7_75t_L g1295 ( 
.A(n_1115),
.Y(n_1295)
);

CKINVDCx16_ASAP7_75t_R g1296 ( 
.A(n_1110),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1125),
.B(n_999),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1134),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1021),
.B(n_1009),
.Y(n_1299)
);

NAND2xp33_ASAP7_75t_SL g1300 ( 
.A(n_1082),
.B(n_1010),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_R g1301 ( 
.A(n_1139),
.B(n_939),
.Y(n_1301)
);

AND3x2_ASAP7_75t_SL g1302 ( 
.A(n_1112),
.B(n_1157),
.C(n_1132),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1081),
.Y(n_1303)
);

NAND2x1_ASAP7_75t_L g1304 ( 
.A(n_1163),
.B(n_852),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1178),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1141),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1075),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1019),
.B(n_888),
.Y(n_1308)
);

AOI211xp5_ASAP7_75t_L g1309 ( 
.A1(n_1057),
.A2(n_889),
.B(n_856),
.C(n_864),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1064),
.A2(n_1066),
.B1(n_1148),
.B2(n_811),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1030),
.B(n_1005),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1103),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1033),
.B(n_806),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1027),
.B(n_1044),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1174),
.B(n_892),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1155),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1223),
.A2(n_1084),
.B(n_939),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1199),
.B(n_1189),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1267),
.B(n_1047),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1251),
.B(n_1180),
.Y(n_1320)
);

O2A1O1Ixp5_ASAP7_75t_L g1321 ( 
.A1(n_1245),
.A2(n_1159),
.B(n_1168),
.C(n_1113),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1198),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1312),
.A2(n_1058),
.A3(n_1089),
.B(n_1083),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_SL g1324 ( 
.A1(n_1282),
.A2(n_1160),
.B(n_1180),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1257),
.A2(n_1117),
.B(n_1106),
.Y(n_1325)
);

AOI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1316),
.A2(n_1094),
.B(n_1093),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1314),
.A2(n_1070),
.B(n_1059),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_1251),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1196),
.B(n_1150),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1304),
.A2(n_1104),
.B(n_1107),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1282),
.A2(n_1175),
.B(n_1169),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1270),
.A2(n_1126),
.B(n_1080),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1286),
.A2(n_1114),
.B(n_1111),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1307),
.A2(n_1187),
.B(n_1181),
.C(n_1090),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1201),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1227),
.B(n_1068),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1255),
.A2(n_1185),
.B(n_1173),
.Y(n_1337)
);

NAND2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1293),
.B(n_811),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1216),
.B(n_1144),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1286),
.A2(n_1131),
.B(n_1127),
.Y(n_1340)
);

AOI221x1_ASAP7_75t_L g1341 ( 
.A1(n_1316),
.A2(n_1191),
.B1(n_1190),
.B2(n_1188),
.C(n_1147),
.Y(n_1341)
);

NAND2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1293),
.B(n_816),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1228),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1198),
.Y(n_1344)
);

OAI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1243),
.A2(n_1042),
.B1(n_1049),
.B2(n_1039),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1272),
.A2(n_1277),
.B(n_1275),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1300),
.A2(n_1054),
.B(n_1052),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1305),
.A2(n_1087),
.B(n_910),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1214),
.B(n_1071),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1221),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1217),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1217),
.A2(n_893),
.A3(n_934),
.B(n_980),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1313),
.A2(n_894),
.B(n_853),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1253),
.A2(n_894),
.B(n_853),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1203),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1256),
.A2(n_1196),
.B1(n_1296),
.B2(n_1210),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_L g1357 ( 
.A1(n_1224),
.A2(n_1029),
.B(n_1063),
.C(n_1056),
.Y(n_1357)
);

AOI211x1_ASAP7_75t_L g1358 ( 
.A1(n_1193),
.A2(n_1074),
.B(n_1086),
.C(n_1065),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1253),
.A2(n_993),
.B(n_986),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1197),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1289),
.A2(n_1004),
.B(n_1086),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1254),
.A2(n_1055),
.B(n_1074),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1200),
.B(n_1079),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1281),
.A2(n_1031),
.A3(n_1006),
.B(n_1077),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1202),
.B(n_1025),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1291),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1213),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1291),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1276),
.A2(n_1311),
.B(n_1273),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1279),
.A2(n_1024),
.B(n_1017),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1287),
.A2(n_1164),
.B(n_1142),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1247),
.Y(n_1372)
);

AO21x1_ASAP7_75t_L g1373 ( 
.A1(n_1216),
.A2(n_1036),
.B(n_816),
.Y(n_1373)
);

AO21x1_ASAP7_75t_L g1374 ( 
.A1(n_1235),
.A2(n_1072),
.B(n_908),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1204),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1297),
.A2(n_1158),
.B(n_1136),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1219),
.A2(n_915),
.B(n_867),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1284),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1247),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1225),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1280),
.A2(n_919),
.B(n_806),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1221),
.A2(n_1051),
.B(n_926),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1205),
.A2(n_926),
.B(n_146),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1294),
.A2(n_926),
.B(n_97),
.C(n_95),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1231),
.A2(n_1250),
.B(n_1244),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1266),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1263),
.A2(n_95),
.B(n_96),
.Y(n_1387)
);

CKINVDCx14_ASAP7_75t_R g1388 ( 
.A(n_1360),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1320),
.B(n_1235),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1386),
.B(n_1262),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1326),
.A2(n_1301),
.B(n_1218),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1375),
.B(n_1238),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1380),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1341),
.A2(n_1229),
.A3(n_1234),
.B(n_1226),
.Y(n_1394)
);

OR2x6_ASAP7_75t_L g1395 ( 
.A(n_1324),
.B(n_1318),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1380),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1336),
.B(n_1233),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1318),
.A2(n_1241),
.B1(n_1215),
.B2(n_1222),
.Y(n_1398)
);

OA21x2_ASAP7_75t_L g1399 ( 
.A1(n_1317),
.A2(n_1310),
.B(n_1195),
.Y(n_1399)
);

NAND2x1p5_ASAP7_75t_L g1400 ( 
.A(n_1343),
.B(n_1192),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1339),
.B(n_1236),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1319),
.B(n_1346),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1355),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1325),
.A2(n_1244),
.B(n_1231),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1384),
.A2(n_1207),
.B(n_1242),
.C(n_1290),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1348),
.A2(n_1274),
.B(n_1246),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1334),
.A2(n_1261),
.A3(n_1240),
.B(n_1265),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1385),
.A2(n_1239),
.B(n_1285),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1339),
.B(n_1236),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1362),
.A2(n_1347),
.B(n_1337),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1322),
.B(n_1237),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1378),
.B(n_1278),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1377),
.A2(n_1244),
.B(n_1231),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1376),
.A2(n_1290),
.B(n_1212),
.Y(n_1414)
);

OAI222xp33_ASAP7_75t_L g1415 ( 
.A1(n_1329),
.A2(n_1259),
.B1(n_1302),
.B2(n_1299),
.C1(n_1298),
.C2(n_1264),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1329),
.B(n_1248),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1369),
.A2(n_1232),
.B1(n_1220),
.B2(n_1271),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1361),
.A2(n_1315),
.B(n_1283),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1322),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1331),
.B(n_1248),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1370),
.A2(n_1308),
.B(n_1309),
.Y(n_1421)
);

AOI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_1363),
.A2(n_1220),
.B1(n_1315),
.B2(n_1258),
.C(n_1208),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1344),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1349),
.B(n_1194),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1367),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1350),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1419),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1393),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1395),
.B(n_1344),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1396),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1395),
.A2(n_1249),
.B1(n_1232),
.B2(n_1328),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1420),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1395),
.B(n_1351),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1423),
.B(n_1351),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1403),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1414),
.A2(n_1374),
.B1(n_1373),
.B2(n_1345),
.Y(n_1436)
);

AO31x2_ASAP7_75t_L g1437 ( 
.A1(n_1410),
.A2(n_1372),
.A3(n_1379),
.B(n_1368),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1394),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1414),
.A2(n_1421),
.B1(n_1398),
.B2(n_1422),
.Y(n_1439)
);

CKINVDCx9p33_ASAP7_75t_R g1440 ( 
.A(n_1390),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1420),
.B(n_1382),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1401),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1415),
.B(n_1230),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1388),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1405),
.A2(n_1321),
.B(n_1387),
.Y(n_1445)
);

INVx5_ASAP7_75t_L g1446 ( 
.A(n_1420),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_SL g1447 ( 
.A(n_1417),
.B(n_1356),
.C(n_1268),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_SL g1448 ( 
.A(n_1417),
.B(n_1211),
.C(n_1209),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1407),
.B(n_1372),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1407),
.B(n_1379),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1416),
.A2(n_1292),
.B1(n_1295),
.B2(n_1303),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1416),
.A2(n_1292),
.B1(n_1258),
.B2(n_1368),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1427),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1445),
.A2(n_1404),
.B(n_1413),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1439),
.A2(n_1416),
.B1(n_1424),
.B2(n_1402),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1452),
.A2(n_1392),
.B(n_1397),
.C(n_1411),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1450),
.B(n_1394),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1446),
.A2(n_1391),
.B(n_1426),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1427),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1447),
.A2(n_1418),
.B1(n_1327),
.B2(n_1306),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1438),
.A2(n_1406),
.B(n_1408),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1450),
.B(n_1394),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1432),
.A2(n_1401),
.B1(n_1409),
.B2(n_1418),
.Y(n_1463)
);

INVx5_ASAP7_75t_L g1464 ( 
.A(n_1446),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1429),
.A2(n_1389),
.B1(n_1409),
.B2(n_1295),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1434),
.B(n_1366),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1448),
.A2(n_1365),
.B1(n_1206),
.B2(n_1425),
.C(n_1357),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1435),
.B(n_1428),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1431),
.A2(n_1389),
.B1(n_1412),
.B2(n_1400),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1437),
.B(n_1399),
.Y(n_1470)
);

BUFx4f_ASAP7_75t_SL g1471 ( 
.A(n_1444),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1429),
.A2(n_1399),
.B1(n_1391),
.B2(n_1371),
.Y(n_1472)
);

OAI322xp33_ASAP7_75t_L g1473 ( 
.A1(n_1443),
.A2(n_1332),
.A3(n_98),
.B1(n_99),
.B2(n_100),
.C1(n_103),
.C2(n_104),
.Y(n_1473)
);

AOI33xp33_ASAP7_75t_L g1474 ( 
.A1(n_1451),
.A2(n_96),
.A3(n_103),
.B1(n_105),
.B2(n_108),
.B3(n_109),
.Y(n_1474)
);

INVx5_ASAP7_75t_SL g1475 ( 
.A(n_1440),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1446),
.A2(n_1299),
.B1(n_1426),
.B2(n_1236),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1446),
.A2(n_1338),
.B1(n_1342),
.B2(n_1358),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1468),
.B(n_1430),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_L g1479 ( 
.A(n_1469),
.B(n_1432),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1457),
.B(n_1446),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1457),
.B(n_1437),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1453),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1453),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1462),
.B(n_1459),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1462),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1429),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1466),
.B(n_1437),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1461),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1470),
.B(n_1437),
.Y(n_1489)
);

AO21x1_ASAP7_75t_SL g1490 ( 
.A1(n_1465),
.A2(n_1442),
.B(n_1449),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1464),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1464),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1464),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1464),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_R g1495 ( 
.A(n_1492),
.B(n_1444),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1485),
.B(n_1470),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1492),
.A2(n_1475),
.B1(n_1456),
.B2(n_1433),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1478),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1485),
.B(n_1475),
.Y(n_1499)
);

NAND3xp33_ASAP7_75t_L g1500 ( 
.A(n_1479),
.B(n_1467),
.C(n_1436),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1493),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1493),
.A2(n_1475),
.B1(n_1455),
.B2(n_1463),
.Y(n_1502)
);

AOI33xp33_ASAP7_75t_L g1503 ( 
.A1(n_1481),
.A2(n_1460),
.A3(n_1433),
.B1(n_1434),
.B2(n_1476),
.B3(n_1472),
.Y(n_1503)
);

AOI211xp5_ASAP7_75t_L g1504 ( 
.A1(n_1491),
.A2(n_1473),
.B(n_1477),
.C(n_1433),
.Y(n_1504)
);

CKINVDCx10_ASAP7_75t_R g1505 ( 
.A(n_1494),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1488),
.A2(n_1454),
.B(n_1458),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1480),
.A2(n_1475),
.B1(n_1441),
.B2(n_1471),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1484),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1484),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1503),
.A2(n_1494),
.B(n_1474),
.C(n_1486),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1509),
.B(n_1481),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1495),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1501),
.B(n_1486),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1502),
.B(n_1486),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1496),
.B(n_1489),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1508),
.B(n_1489),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1498),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1501),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1480),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1500),
.B(n_1480),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1501),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1495),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1506),
.B(n_1487),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1506),
.B(n_1482),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1506),
.B(n_1490),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1517),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_R g1527 ( 
.A(n_1522),
.B(n_1505),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1512),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1516),
.B(n_1483),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1511),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1524),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1511),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1515),
.Y(n_1533)
);

OAI21xp33_ASAP7_75t_L g1534 ( 
.A1(n_1528),
.A2(n_1514),
.B(n_1520),
.Y(n_1534)
);

OR3x1_ASAP7_75t_L g1535 ( 
.A(n_1527),
.B(n_1520),
.C(n_1510),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1528),
.B(n_1520),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1526),
.Y(n_1537)
);

AOI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1535),
.A2(n_1523),
.B1(n_1510),
.B2(n_1531),
.C(n_1525),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1536),
.B(n_1523),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1537),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1538),
.B(n_1534),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1539),
.A2(n_1535),
.B1(n_1520),
.B2(n_1525),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1540),
.B(n_1531),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1540),
.B(n_1530),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1543),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1544),
.Y(n_1546)
);

XNOR2xp5_ASAP7_75t_L g1547 ( 
.A(n_1541),
.B(n_1497),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1542),
.B(n_1532),
.Y(n_1548)
);

XNOR2xp5_ASAP7_75t_L g1549 ( 
.A(n_1541),
.B(n_1507),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1541),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1543),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1545),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1550),
.B(n_1533),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1546),
.B(n_1503),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1551),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1547),
.B(n_1335),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1545),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_SL g1560 ( 
.A(n_1546),
.B(n_1504),
.C(n_1518),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1560),
.A2(n_1557),
.B1(n_1554),
.B2(n_1553),
.Y(n_1561)
);

O2A1O1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1552),
.A2(n_1559),
.B(n_1555),
.C(n_1560),
.Y(n_1562)
);

OAI31xp33_ASAP7_75t_L g1563 ( 
.A1(n_1558),
.A2(n_1513),
.A3(n_1519),
.B(n_1529),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1556),
.B(n_1513),
.Y(n_1564)
);

AOI211x1_ASAP7_75t_SL g1565 ( 
.A1(n_1553),
.A2(n_112),
.B(n_108),
.C(n_110),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_R g1566 ( 
.A(n_1552),
.B(n_110),
.Y(n_1566)
);

AOI221x1_ASAP7_75t_L g1567 ( 
.A1(n_1552),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.C(n_116),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1556),
.B(n_114),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1568),
.B(n_115),
.Y(n_1569)
);

OAI21xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1561),
.A2(n_1441),
.B(n_1490),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1565),
.B(n_119),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1562),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1567),
.Y(n_1573)
);

OAI211xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1563),
.A2(n_127),
.B(n_121),
.C(n_125),
.Y(n_1574)
);

OAI322xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1564),
.A2(n_127),
.A3(n_1441),
.B1(n_1437),
.B2(n_1364),
.C1(n_1383),
.C2(n_1323),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1566),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1568),
.Y(n_1577)
);

AOI211xp5_ASAP7_75t_L g1578 ( 
.A1(n_1572),
.A2(n_1340),
.B(n_1333),
.C(n_1353),
.Y(n_1578)
);

AO22x1_ASAP7_75t_L g1579 ( 
.A1(n_1573),
.A2(n_1269),
.B1(n_1252),
.B2(n_1260),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_SL g1580 ( 
.A(n_1571),
.B(n_143),
.C(n_147),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1569),
.A2(n_1260),
.B1(n_1269),
.B2(n_1288),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1576),
.B(n_148),
.Y(n_1582)
);

AO22x2_ASAP7_75t_L g1583 ( 
.A1(n_1577),
.A2(n_1364),
.B1(n_1323),
.B2(n_1352),
.Y(n_1583)
);

NOR3xp33_ASAP7_75t_L g1584 ( 
.A(n_1574),
.B(n_1330),
.C(n_1354),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1575),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1570),
.B(n_151),
.Y(n_1586)
);

NAND4xp25_ASAP7_75t_L g1587 ( 
.A(n_1586),
.B(n_152),
.C(n_153),
.D(n_154),
.Y(n_1587)
);

AOI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1580),
.A2(n_155),
.B1(n_160),
.B2(n_163),
.C(n_164),
.Y(n_1588)
);

XNOR2xp5_ASAP7_75t_L g1589 ( 
.A(n_1585),
.B(n_167),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1582),
.B(n_1381),
.C(n_1359),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1579),
.B(n_169),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1584),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.C(n_177),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1589),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1587),
.A2(n_1578),
.B(n_1581),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1591),
.B(n_1583),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1588),
.B(n_1583),
.C(n_178),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1590),
.B(n_189),
.Y(n_1597)
);

CKINVDCx16_ASAP7_75t_R g1598 ( 
.A(n_1592),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_L g1599 ( 
.A(n_1596),
.B(n_1593),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1598),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1597),
.Y(n_1601)
);

NOR2xp67_ASAP7_75t_L g1602 ( 
.A(n_1595),
.B(n_191),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1602),
.A2(n_1594),
.B(n_192),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1600),
.A2(n_1352),
.B1(n_194),
.B2(n_195),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1603),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_SL g1606 ( 
.A(n_1604),
.B(n_1601),
.C(n_1599),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1605),
.Y(n_1607)
);

AOI222xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1607),
.A2(n_1606),
.B1(n_197),
.B2(n_200),
.C1(n_202),
.C2(n_203),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1608),
.B(n_205),
.C(n_211),
.Y(n_1609)
);

AOI322xp5_ASAP7_75t_L g1610 ( 
.A1(n_1608),
.A2(n_212),
.A3(n_215),
.B1(n_217),
.B2(n_220),
.C1(n_222),
.C2(n_224),
.Y(n_1610)
);

AOI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1609),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.C(n_237),
.Y(n_1611)
);

AOI211xp5_ASAP7_75t_L g1612 ( 
.A1(n_1611),
.A2(n_1610),
.B(n_243),
.C(n_245),
.Y(n_1612)
);


endmodule