module real_aes_10079_n_15 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_15);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_15;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_55;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_33;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_54;
wire n_51;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_50;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_53;
wire n_36;
NOR2xp33_ASAP7_75t_R g22 ( .A(n_0), .B(n_5), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_1), .B(n_7), .C(n_21), .Y(n_20) );
NOR3xp33_ASAP7_75t_SL g51 ( .A(n_1), .B(n_10), .C(n_52), .Y(n_51) );
NAND2xp33_ASAP7_75t_R g21 ( .A(n_2), .B(n_22), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g54 ( .A(n_2), .Y(n_54) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_3), .Y(n_23) );
NOR4xp25_ASAP7_75t_SL g49 ( .A(n_3), .B(n_50), .C(n_53), .D(n_54), .Y(n_49) );
NOR4xp25_ASAP7_75t_SL g18 ( .A(n_4), .B(n_19), .C(n_23), .D(n_24), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g53 ( .A(n_4), .Y(n_53) );
NOR2xp33_ASAP7_75t_R g17 ( .A(n_6), .B(n_11), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g28 ( .A(n_6), .B(n_11), .Y(n_28) );
NAND2xp33_ASAP7_75t_SL g33 ( .A(n_6), .B(n_34), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g38 ( .A(n_6), .B(n_34), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g55 ( .A(n_7), .Y(n_55) );
AOI322xp5_ASAP7_75t_SL g31 ( .A1(n_8), .A2(n_13), .A3(n_18), .B1(n_32), .B2(n_35), .C1(n_39), .C2(n_46), .Y(n_31) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_9), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_10), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_11), .Y(n_34) );
BUFx2_ASAP7_75t_L g45 ( .A(n_12), .Y(n_45) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_14), .Y(n_30) );
OAI221xp5_ASAP7_75t_L g15 ( .A1(n_16), .A2(n_25), .B1(n_26), .B2(n_30), .C(n_31), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_17), .B(n_18), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g47 ( .A(n_17), .Y(n_47) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_18), .Y(n_29) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_18), .B(n_38), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g52 ( .A(n_22), .Y(n_52) );
INVxp33_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
NOR2xp33_ASAP7_75t_R g27 ( .A(n_28), .B(n_29), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
INVx1_ASAP7_75t_SL g39 ( .A(n_40), .Y(n_39) );
INVx1_ASAP7_75t_SL g40 ( .A(n_41), .Y(n_40) );
INVx5_ASAP7_75t_L g41 ( .A(n_42), .Y(n_41) );
BUFx8_ASAP7_75t_SL g42 ( .A(n_43), .Y(n_42) );
INVx2_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
BUFx2_ASAP7_75t_L g44 ( .A(n_45), .Y(n_44) );
NOR2xp33_ASAP7_75t_R g46 ( .A(n_47), .B(n_48), .Y(n_46) );
NAND2xp33_ASAP7_75t_R g48 ( .A(n_49), .B(n_55), .Y(n_48) );
CKINVDCx5p33_ASAP7_75t_R g50 ( .A(n_51), .Y(n_50) );
endmodule