module fake_jpeg_12055_n_479 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_479);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_479;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_50),
.Y(n_152)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_56),
.Y(n_104)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_74),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_23),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_62),
.B(n_69),
.Y(n_135)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_91),
.Y(n_101)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_81),
.Y(n_141)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_84),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_0),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_20),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_89),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NAND2x1_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_93),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_20),
.A2(n_14),
.B(n_3),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_30),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_2),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_19),
.B1(n_41),
.B2(n_30),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_98),
.A2(n_108),
.B1(n_118),
.B2(n_124),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_45),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_100),
.B(n_105),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_19),
.B1(n_41),
.B2(n_48),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_35),
.B1(n_41),
.B2(n_38),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_110),
.A2(n_126),
.B1(n_139),
.B2(n_150),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_35),
.B1(n_41),
.B2(n_38),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_132),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_17),
.B1(n_46),
.B2(n_31),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_115),
.A2(n_116),
.B1(n_140),
.B2(n_85),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_51),
.B1(n_81),
.B2(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_131),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_76),
.A2(n_48),
.B1(n_25),
.B2(n_43),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_46),
.B1(n_27),
.B2(n_31),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_82),
.A2(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_58),
.A2(n_42),
.B(n_40),
.C(n_39),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_130),
.B(n_144),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_39),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_34),
.B1(n_28),
.B2(n_25),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_84),
.A2(n_34),
.B1(n_28),
.B2(n_5),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_95),
.B1(n_97),
.B2(n_79),
.Y(n_160)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_59),
.B(n_2),
.CON(n_144),
.SN(n_144)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_65),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_64),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_61),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_154),
.B(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_5),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_175),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_71),
.B1(n_68),
.B2(n_57),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_158),
.A2(n_140),
.B1(n_114),
.B2(n_134),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_159),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_186),
.B1(n_188),
.B2(n_100),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_190),
.Y(n_236)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_169),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_122),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_170),
.B(n_184),
.Y(n_244)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_171),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_6),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_6),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_203),
.Y(n_207)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_104),
.B(n_92),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_137),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_101),
.A2(n_92),
.B1(n_85),
.B2(n_73),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_121),
.B(n_73),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_189),
.B(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

BUFx16f_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_115),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_123),
.B(n_138),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_105),
.B(n_65),
.C(n_61),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_202),
.C(n_144),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_137),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_197),
.B(n_200),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_116),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_199),
.B1(n_127),
.B2(n_134),
.Y(n_209)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_135),
.B(n_7),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_201),
.B(n_125),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_100),
.B(n_9),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_135),
.B(n_10),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_204),
.A2(n_243),
.B1(n_246),
.B2(n_202),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_146),
.B1(n_116),
.B2(n_127),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_205),
.A2(n_210),
.B1(n_226),
.B2(n_201),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_135),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_215),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_102),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_102),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_235),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_202),
.C(n_182),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_107),
.B1(n_142),
.B2(n_133),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_141),
.B(n_113),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_231),
.A2(n_237),
.B(n_194),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_190),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_234),
.B(n_245),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_157),
.B(n_107),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_194),
.A2(n_113),
.B1(n_136),
.B2(n_138),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_162),
.A2(n_174),
.B1(n_168),
.B2(n_175),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_162),
.A2(n_142),
.B1(n_133),
.B2(n_129),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_263),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_257),
.C(n_285),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_166),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_251),
.Y(n_303)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_182),
.C(n_196),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_264),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_259),
.A2(n_276),
.B1(n_283),
.B2(n_223),
.Y(n_299)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_180),
.B(n_182),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_261),
.A2(n_250),
.B(n_256),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_262),
.A2(n_270),
.B1(n_268),
.B2(n_282),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_191),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_211),
.A2(n_161),
.B(n_195),
.C(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_195),
.B1(n_178),
.B2(n_179),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_277),
.B1(n_278),
.B2(n_226),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_217),
.B1(n_232),
.B2(n_204),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_274),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_216),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_273),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_216),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_164),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_210),
.A2(n_185),
.B1(n_155),
.B2(n_173),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_215),
.A2(n_193),
.B1(n_199),
.B2(n_167),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_233),
.A2(n_171),
.B1(n_125),
.B2(n_136),
.Y(n_278)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_214),
.B(n_181),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_282),
.Y(n_308)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_236),
.A2(n_123),
.B1(n_176),
.B2(n_172),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_222),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_206),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_159),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_206),
.B(n_163),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_207),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_291),
.B(n_265),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_231),
.B(n_237),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_295),
.A2(n_298),
.B(n_300),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_271),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_302),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_241),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_299),
.A2(n_277),
.B1(n_253),
.B2(n_278),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_274),
.A2(n_225),
.B(n_222),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_306),
.A2(n_309),
.B(n_319),
.Y(n_342)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_269),
.A2(n_241),
.B(n_225),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_320),
.B1(n_283),
.B2(n_276),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_321),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_259),
.A2(n_207),
.B1(n_219),
.B2(n_230),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_315),
.A2(n_299),
.B1(n_321),
.B2(n_308),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_257),
.B(n_208),
.C(n_219),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_323),
.C(n_293),
.Y(n_339)
);

AO22x1_ASAP7_75t_L g319 ( 
.A1(n_264),
.A2(n_242),
.B1(n_224),
.B2(n_223),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_262),
.A2(n_218),
.B1(n_224),
.B2(n_227),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_287),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_261),
.B(n_242),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_324),
.A2(n_325),
.B1(n_333),
.B2(n_337),
.Y(n_363)
);

OAI221xp5_ASAP7_75t_L g325 ( 
.A1(n_306),
.A2(n_280),
.B1(n_256),
.B2(n_267),
.C(n_260),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_290),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_326),
.B(n_327),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_288),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_329),
.B(n_331),
.Y(n_381)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_255),
.B1(n_267),
.B2(n_266),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_275),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_339),
.C(n_345),
.Y(n_373)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_336),
.B(n_340),
.Y(n_372)
);

AOI22x1_ASAP7_75t_L g337 ( 
.A1(n_316),
.A2(n_255),
.B1(n_252),
.B2(n_254),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_343),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_291),
.B(n_249),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_305),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_273),
.C(n_272),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_281),
.Y(n_346)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_347),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g348 ( 
.A1(n_316),
.A2(n_238),
.B(n_213),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_348),
.A2(n_319),
.B(n_312),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_308),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_349),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_279),
.Y(n_350)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_315),
.A2(n_279),
.B1(n_218),
.B2(n_227),
.Y(n_351)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_323),
.B(n_227),
.Y(n_352)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_314),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_248),
.Y(n_354)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_353),
.B(n_303),
.C(n_300),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_355),
.B(n_359),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_327),
.B(n_326),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_338),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_344),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_328),
.A2(n_298),
.B1(n_295),
.B2(n_309),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_360),
.A2(n_369),
.B1(n_376),
.B2(n_332),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_362),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_298),
.B1(n_301),
.B2(n_318),
.Y(n_364)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_316),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_366),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_331),
.A2(n_301),
.B1(n_322),
.B2(n_318),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_319),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_382),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_324),
.A2(n_344),
.B1(n_349),
.B2(n_333),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_377),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_322),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_383),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_357),
.A2(n_329),
.B1(n_346),
.B2(n_350),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_384),
.A2(n_390),
.B1(n_392),
.B2(n_400),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_361),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_387),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_341),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_389),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_345),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_341),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_357),
.A2(n_354),
.B1(n_342),
.B2(n_337),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_381),
.A2(n_342),
.B1(n_337),
.B2(n_352),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_381),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g406 ( 
.A(n_394),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_336),
.C(n_348),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_397),
.C(n_398),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_366),
.C(n_382),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_347),
.C(n_335),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_351),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_405),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_362),
.A2(n_313),
.B1(n_307),
.B2(n_312),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_402),
.A2(n_370),
.B1(n_368),
.B2(n_367),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_358),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_404),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_379),
.Y(n_405)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_391),
.B(n_372),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_410),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_363),
.Y(n_410)
);

AO21x1_ASAP7_75t_L g411 ( 
.A1(n_395),
.A2(n_368),
.B(n_367),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_411),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_399),
.A2(n_370),
.B1(n_376),
.B2(n_377),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_401),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_380),
.C(n_374),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_420),
.C(n_398),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_395),
.A2(n_371),
.B(n_289),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_419),
.A2(n_390),
.B(n_402),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_289),
.C(n_292),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_296),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_405),
.Y(n_432)
);

AO221x1_ASAP7_75t_L g423 ( 
.A1(n_388),
.A2(n_296),
.B1(n_292),
.B2(n_228),
.C(n_238),
.Y(n_423)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_435),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_418),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_430),
.Y(n_442)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_429),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_421),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_412),
.A2(n_393),
.B1(n_396),
.B2(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_431),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_410),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_433),
.A2(n_416),
.B(n_407),
.Y(n_450)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_437),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_413),
.A2(n_392),
.B1(n_403),
.B2(n_247),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_403),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_228),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_438),
.A2(n_419),
.B(n_427),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_414),
.C(n_420),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_447),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_417),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_441),
.A2(n_446),
.B(n_449),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_228),
.Y(n_460)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_415),
.C(n_409),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_448),
.B(n_425),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_436),
.A2(n_415),
.B(n_409),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_450),
.A2(n_422),
.B(n_432),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_428),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_453),
.B(n_458),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_443),
.A2(n_433),
.B1(n_436),
.B2(n_428),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_454),
.A2(n_455),
.B1(n_441),
.B2(n_451),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_450),
.A2(n_413),
.B1(n_429),
.B2(n_438),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_460),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_442),
.B(n_408),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_440),
.A2(n_216),
.B(n_191),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_445),
.C(n_448),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_447),
.Y(n_463)
);

OAI221xp5_ASAP7_75t_L g470 ( 
.A1(n_463),
.A2(n_464),
.B1(n_467),
.B2(n_459),
.C(n_462),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_451),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_466),
.C(n_444),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g469 ( 
.A1(n_468),
.A2(n_467),
.B(n_457),
.Y(n_469)
);

A2O1A1O1Ixp25_ASAP7_75t_L g473 ( 
.A1(n_469),
.A2(n_471),
.B(n_472),
.C(n_452),
.D(n_460),
.Y(n_473)
);

OAI311xp33_ASAP7_75t_L g474 ( 
.A1(n_470),
.A2(n_213),
.A3(n_12),
.B1(n_13),
.C1(n_14),
.Y(n_474)
);

NOR2x1_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_455),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_473),
.B(n_474),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

AOI221xp5_ASAP7_75t_L g477 ( 
.A1(n_475),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_476),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_11),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_11),
.Y(n_479)
);


endmodule