module fake_jpeg_12818_n_393 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_393);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_393;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_46),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_29),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g107 ( 
.A(n_50),
.Y(n_107)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_10),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_59),
.B(n_64),
.Y(n_112)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_30),
.B(n_7),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_68),
.B(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2x1_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_7),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_75),
.Y(n_91)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_38),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_0),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_41),
.B1(n_37),
.B2(n_33),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_90),
.B1(n_106),
.B2(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_44),
.A2(n_38),
.B1(n_41),
.B2(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_18),
.B1(n_19),
.B2(n_38),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_95),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_42),
.B1(n_40),
.B2(n_34),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_41),
.B1(n_33),
.B2(n_37),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_96),
.A2(n_99),
.B1(n_101),
.B2(n_17),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_37),
.B1(n_33),
.B2(n_40),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_73),
.A2(n_27),
.B1(n_39),
.B2(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_109),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_45),
.A2(n_32),
.B1(n_17),
.B2(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_36),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_47),
.A2(n_17),
.B1(n_32),
.B2(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_0),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_32),
.B1(n_17),
.B2(n_11),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_121),
.A2(n_62),
.B1(n_46),
.B2(n_66),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_50),
.B(n_11),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_50),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_0),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_79),
.B1(n_77),
.B2(n_76),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_128),
.A2(n_150),
.B1(n_86),
.B2(n_126),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_136),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_1),
.B(n_2),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_154),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_133),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_135),
.A2(n_98),
.B1(n_115),
.B2(n_82),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_91),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_145),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_147),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_92),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_1),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_153),
.Y(n_183)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_17),
.B1(n_32),
.B2(n_1),
.Y(n_150)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_3),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_119),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_157),
.Y(n_184)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_15),
.Y(n_205)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_87),
.B(n_89),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_4),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_163),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_92),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_4),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_4),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_126),
.B1(n_105),
.B2(n_108),
.Y(n_171)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_83),
.B(n_5),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_7),
.Y(n_188)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_16),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_93),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_175),
.C(n_209),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_83),
.C(n_95),
.Y(n_175)
);

AND2x4_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_108),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_192),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_127),
.A2(n_104),
.B1(n_82),
.B2(n_118),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_138),
.B1(n_169),
.B2(n_152),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_86),
.B(n_98),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_127),
.B(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_188),
.B(n_207),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_206),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_197),
.A2(n_198),
.B1(n_189),
.B2(n_192),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_134),
.A2(n_120),
.B1(n_118),
.B2(n_85),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_200),
.B1(n_151),
.B2(n_149),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_130),
.A2(n_120),
.B1(n_13),
.B2(n_14),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_143),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_137),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_139),
.B(n_16),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_212),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_182),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_233),
.B(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_231),
.B1(n_238),
.B2(n_206),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_132),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_219),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_141),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_139),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_223),
.B(n_227),
.Y(n_267)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_173),
.B(n_148),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_183),
.B(n_153),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_228),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_173),
.B(n_154),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_189),
.B1(n_199),
.B2(n_205),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_175),
.A2(n_142),
.B1(n_158),
.B2(n_157),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_180),
.A2(n_179),
.B(n_195),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_167),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_209),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_237),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_177),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_179),
.A2(n_156),
.B1(n_159),
.B2(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_194),
.B(n_187),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_197),
.B1(n_199),
.B2(n_202),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_176),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_184),
.Y(n_261)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_244),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_190),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_252),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_172),
.C(n_195),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_266),
.C(n_239),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_234),
.B1(n_214),
.B2(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_258),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_210),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_220),
.Y(n_252)
);

BUFx8_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_254),
.A2(n_257),
.B1(n_268),
.B2(n_272),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_210),
.A2(n_230),
.B1(n_243),
.B2(n_232),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_220),
.Y(n_258)
);

BUFx12_ASAP7_75t_L g259 ( 
.A(n_211),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_219),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_201),
.C(n_184),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_242),
.A2(n_196),
.B1(n_201),
.B2(n_202),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_274),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_196),
.B1(n_191),
.B2(n_181),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_191),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_203),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_275),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_273),
.A2(n_264),
.B(n_257),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_274),
.Y(n_320)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_260),
.B1(n_252),
.B2(n_268),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_269),
.A2(n_232),
.B1(n_236),
.B2(n_210),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_296),
.B(n_260),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_288),
.C(n_290),
.Y(n_306)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_294),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_235),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_219),
.B(n_236),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_271),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_250),
.A2(n_213),
.B(n_216),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_228),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_231),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_225),
.C(n_254),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_265),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_258),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_307),
.A2(n_303),
.B1(n_291),
.B2(n_302),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_262),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_310),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_270),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_317),
.C(n_290),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_282),
.B(n_262),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_312),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_278),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_246),
.Y(n_314)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_296),
.Y(n_315)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_217),
.Y(n_316)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_225),
.C(n_212),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_248),
.Y(n_318)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_319),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_320),
.B(n_287),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_221),
.Y(n_322)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_326),
.C(n_329),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_299),
.C(n_292),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_292),
.C(n_281),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_309),
.C(n_313),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_331),
.B(n_338),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_314),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_304),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_336),
.A2(n_307),
.B(n_303),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_311),
.A2(n_295),
.B1(n_280),
.B2(n_293),
.Y(n_337)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_302),
.A2(n_293),
.B1(n_287),
.B2(n_284),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_328),
.B(n_305),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_341),
.B(n_351),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_320),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_344),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_304),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_348),
.C(n_335),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_346),
.B(n_350),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_310),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_314),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_330),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_352),
.B(n_353),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_301),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_334),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_340),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_347),
.A2(n_340),
.B1(n_324),
.B2(n_325),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_361),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_349),
.C(n_350),
.Y(n_367)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_363),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_349),
.B(n_332),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_339),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_364),
.B(n_316),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_338),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_370),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_368),
.B(n_369),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_365),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_342),
.C(n_343),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_360),
.A2(n_329),
.B(n_279),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_371),
.A2(n_372),
.B(n_373),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_364),
.A2(n_279),
.B(n_259),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_355),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_359),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_375),
.A2(n_357),
.B(n_359),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_377),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_321),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_382),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_316),
.B1(n_300),
.B2(n_289),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_381),
.A2(n_368),
.B1(n_286),
.B2(n_265),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_383),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_386),
.B(n_382),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_379),
.B(n_256),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_389),
.C(n_253),
.Y(n_390)
);

OAI311xp33_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_380),
.A3(n_259),
.B1(n_253),
.C1(n_256),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_390),
.A2(n_387),
.B(n_222),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_203),
.B(n_208),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_208),
.Y(n_393)
);


endmodule