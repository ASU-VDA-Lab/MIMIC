module fake_jpeg_27637_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_9),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_16),
.CON(n_57),
.SN(n_57)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_24),
.C(n_27),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_41),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_61),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_31),
.B1(n_23),
.B2(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_61)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_39),
.C(n_35),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_65),
.B(n_75),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_46),
.B1(n_50),
.B2(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_80),
.B1(n_37),
.B2(n_38),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_84),
.B(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_76),
.B(n_85),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_34),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_37),
.B1(n_38),
.B2(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_45),
.Y(n_94)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_88),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_39),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_85),
.B(n_60),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_44),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_37),
.B1(n_38),
.B2(n_36),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_110),
.B1(n_117),
.B2(n_49),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_100),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_26),
.B(n_17),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_97),
.A2(n_107),
.B(n_116),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_37),
.B1(n_38),
.B2(n_62),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_104),
.B1(n_106),
.B2(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_82),
.B1(n_70),
.B2(n_56),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_27),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_32),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_41),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_66),
.B1(n_79),
.B2(n_76),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_37),
.B1(n_39),
.B2(n_59),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_39),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_87),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_37),
.B1(n_39),
.B2(n_51),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_90),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_69),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_39),
.B1(n_58),
.B2(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_118),
.B(n_69),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_125),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_99),
.B1(n_112),
.B2(n_67),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_130),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_104),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_127),
.B1(n_146),
.B2(n_101),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_64),
.B1(n_84),
.B2(n_73),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_65),
.B(n_70),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_141),
.B(n_16),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_41),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_19),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_41),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_140),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_58),
.B1(n_90),
.B2(n_19),
.Y(n_178)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_143),
.B(n_63),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_0),
.B(n_1),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_32),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_9),
.C(n_15),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_19),
.B(n_25),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_51),
.B1(n_78),
.B2(n_67),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_32),
.C(n_24),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_98),
.C(n_107),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_151),
.B1(n_170),
.B2(n_134),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_40),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_158),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_91),
.C(n_107),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_168),
.C(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_122),
.B1(n_138),
.B2(n_136),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_178),
.B1(n_90),
.B2(n_25),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_166),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_25),
.B(n_33),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_171),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_91),
.C(n_95),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_95),
.C(n_35),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_92),
.B1(n_112),
.B2(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_93),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_179),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_112),
.B1(n_78),
.B2(n_89),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_175),
.A2(n_123),
.B1(n_147),
.B2(n_139),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_18),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_32),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_183),
.B(n_185),
.Y(n_208)
);

AO32x1_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_134),
.A3(n_139),
.B1(n_141),
.B2(n_135),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_188),
.B1(n_192),
.B2(n_200),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_123),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_194),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_195),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_165),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_18),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_206),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_28),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_160),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_16),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_17),
.B1(n_33),
.B2(n_29),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_207),
.A2(n_160),
.B1(n_17),
.B2(n_33),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_168),
.C(n_149),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_215),
.C(n_219),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_213),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_163),
.B(n_153),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_221),
.B1(n_207),
.B2(n_204),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_154),
.C(n_179),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_198),
.B(n_180),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_167),
.C(n_40),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_152),
.B1(n_29),
.B2(n_18),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_40),
.C(n_35),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_226),
.C(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_40),
.C(n_35),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_40),
.C(n_152),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_40),
.C(n_24),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_231),
.C(n_205),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_28),
.C(n_29),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_196),
.Y(n_246)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_234),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_188),
.B1(n_206),
.B2(n_183),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_184),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_242),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_185),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_251),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_181),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_250),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_248),
.A2(n_208),
.B1(n_231),
.B2(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_252),
.C(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_193),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_187),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_12),
.B1(n_10),
.B2(n_8),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_14),
.C(n_13),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_209),
.C(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_265),
.C(n_241),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_215),
.C(n_219),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_223),
.C(n_229),
.Y(n_258)
);

OAI22x1_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_28),
.B1(n_10),
.B2(n_8),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_225),
.B(n_2),
.C(n_3),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_239),
.B(n_244),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_20),
.C(n_26),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_20),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_251),
.C(n_233),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_276),
.C(n_261),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_278),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_280),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_236),
.B1(n_245),
.B2(n_248),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_246),
.C(n_26),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_13),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_12),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_261),
.B1(n_10),
.B2(n_8),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_2),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_273),
.A2(n_267),
.B1(n_268),
.B2(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_282),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_289),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_264),
.C(n_2),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_291),
.Y(n_301)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_264),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_7),
.C(n_2),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_1),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_5),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_269),
.B1(n_3),
.B2(n_4),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_299),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_3),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_300),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_4),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_289),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.Y(n_304)
);

OAI21x1_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_283),
.B(n_285),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_305),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_301),
.C(n_287),
.Y(n_311)
);

AOI31xp33_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.A3(n_309),
.B(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_290),
.C(n_293),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_310),
.B(n_304),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_6),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_7),
.Y(n_317)
);


endmodule