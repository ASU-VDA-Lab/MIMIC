module fake_jpeg_23530_n_114 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx5_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_19),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_24),
.C(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_19),
.B1(n_13),
.B2(n_21),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_17),
.B1(n_13),
.B2(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_44),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_20),
.B1(n_26),
.B2(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_34),
.B1(n_33),
.B2(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_35),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_47),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_43),
.B1(n_46),
.B2(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_58),
.B(n_48),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_14),
.B(n_12),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_23),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_29),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_15),
.C(n_11),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_56),
.A3(n_23),
.B1(n_29),
.B2(n_14),
.C1(n_12),
.C2(n_11),
.Y(n_77)
);

OA21x2_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_65),
.B(n_66),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_80),
.B(n_0),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_87),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_62),
.B1(n_63),
.B2(n_29),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_74),
.B1(n_70),
.B2(n_71),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_61),
.C(n_29),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_83),
.C(n_88),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

OAI322xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_78),
.A3(n_85),
.B1(n_88),
.B2(n_82),
.C1(n_86),
.C2(n_89),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_9),
.B(n_8),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_96),
.C(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_9),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_39),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_91),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_106),
.C(n_4),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

OAI31xp33_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_4),
.C(n_5),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_105),
.B(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_107),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_111),
.C(n_104),
.Y(n_114)
);


endmodule