module real_jpeg_25059_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_34),
.B1(n_39),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_34),
.B1(n_73),
.B2(n_75),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_34),
.B1(n_54),
.B2(n_57),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_46),
.B1(n_54),
.B2(n_57),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_46),
.B1(n_68),
.B2(n_73),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_2),
.A2(n_65),
.B(n_129),
.C(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_2),
.B(n_63),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_2),
.A2(n_52),
.B(n_54),
.C(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_2),
.B(n_23),
.C(n_42),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_2),
.B(n_152),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_82),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_2),
.B(n_44),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_25),
.B1(n_39),
.B2(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_54),
.B1(n_57),
.B2(n_69),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_39),
.B1(n_43),
.B2(n_69),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_69),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_135),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_134),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_111),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_16),
.B(n_111),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_77),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_49),
.C(n_61),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_18),
.A2(n_19),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_35),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_28),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_21),
.A2(n_86),
.B(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_22),
.A2(n_23),
.B1(n_41),
.B2(n_42),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_23),
.B(n_221),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_33),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_26),
.A2(n_85),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_26),
.B(n_85),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_26),
.B(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_27),
.Y(n_132)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_27),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_29),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_29),
.B(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_47),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_36),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_45),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_37),
.B(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_37),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_43),
.B1(n_52),
.B2(n_56),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_39),
.B(n_197),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_43),
.A2(n_46),
.B(n_56),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_44),
.B(n_184),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_45),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_46),
.A2(n_54),
.B(n_64),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_47),
.A2(n_89),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_47),
.B(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_49),
.A2(n_61),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_49),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_58),
.B(n_59),
.Y(n_49)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_50),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_50),
.B(n_100),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_54),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_59),
.Y(n_126)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_63),
.B(n_74),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_65),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_71),
.Y(n_96)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_95),
.Y(n_144)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_104),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_87),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_87),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_81),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_86),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_109),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_88),
.B(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_90),
.B(n_194),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_99),
.B(n_123),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_102),
.B(n_151),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_105),
.A2(n_110),
.B1(n_178),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.C(n_133),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_112),
.A2(n_113),
.B1(n_133),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_118),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_131),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_133),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_171),
.B(n_246),
.C(n_251),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_159),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_137),
.B(n_159),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_155),
.B2(n_158),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_153),
.B2(n_154),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_140),
.B(n_154),
.C(n_158),
.Y(n_247)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_148),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_143),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.C(n_166),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_161),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_166),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.C(n_169),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_245),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_188),
.B(n_244),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_185),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_174),
.B(n_185),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_180),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_180),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_178),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_239),
.B(n_243),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_230),
.B(n_238),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_211),
.B(n_229),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_192),
.B(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_193),
.A2(n_195),
.B1(n_196),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_205),
.B2(n_210),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_201),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_204),
.C(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_218),
.B(n_228),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_224),
.B(n_227),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_232),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_240),
.B(n_241),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);


endmodule