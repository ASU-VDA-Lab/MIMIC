module real_aes_16222_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_858, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_858;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_0), .Y(n_569) );
AND2x4_ASAP7_75t_L g854 ( .A(n_1), .B(n_855), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g113 ( .A1(n_2), .A2(n_114), .B1(n_115), .B2(n_474), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_2), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_3), .A2(n_4), .B1(n_230), .B2(n_231), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_5), .A2(n_22), .B1(n_131), .B2(n_143), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_6), .A2(n_52), .B1(n_163), .B2(n_164), .Y(n_162) );
BUFx3_ASAP7_75t_L g526 ( .A(n_7), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_8), .A2(n_14), .B1(n_140), .B2(n_180), .Y(n_195) );
INVx1_ASAP7_75t_L g855 ( .A(n_9), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_10), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_11), .B(n_187), .Y(n_511) );
OR2x2_ASAP7_75t_L g108 ( .A(n_12), .B(n_31), .Y(n_108) );
BUFx2_ASAP7_75t_L g851 ( .A(n_12), .Y(n_851) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_13), .Y(n_132) );
OAI22xp33_ASAP7_75t_SL g479 ( .A1(n_15), .A2(n_480), .B1(n_481), .B2(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_15), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_15), .A2(n_480), .B1(n_494), .B2(n_831), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_16), .B(n_170), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_17), .B(n_208), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_18), .A2(n_84), .B1(n_143), .B2(n_170), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_19), .Y(n_109) );
OAI21x1_ASAP7_75t_L g125 ( .A1(n_20), .A2(n_48), .B(n_126), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_21), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_23), .B(n_131), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_24), .B(n_138), .Y(n_254) );
INVx4_ASAP7_75t_R g216 ( .A(n_25), .Y(n_216) );
AO32x2_ASAP7_75t_L g572 ( .A1(n_26), .A2(n_149), .A3(n_150), .B1(n_573), .B2(n_576), .Y(n_572) );
AO32x1_ASAP7_75t_L g609 ( .A1(n_26), .A2(n_149), .A3(n_150), .B1(n_573), .B2(n_576), .Y(n_609) );
INVx1_ASAP7_75t_L g235 ( .A(n_27), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_28), .B(n_131), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_SL g139 ( .A1(n_29), .A2(n_140), .B(n_141), .C(n_144), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_30), .A2(n_45), .B1(n_140), .B2(n_198), .Y(n_303) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_31), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_32), .Y(n_135) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_33), .A2(n_51), .B1(n_131), .B2(n_217), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_34), .A2(n_89), .B1(n_143), .B2(n_198), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_35), .B(n_513), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_36), .B(n_548), .Y(n_598) );
INVx1_ASAP7_75t_L g257 ( .A(n_37), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_38), .B(n_140), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_39), .A2(n_66), .B1(n_198), .B2(n_581), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_40), .Y(n_181) );
INVx2_ASAP7_75t_L g477 ( .A(n_41), .Y(n_477) );
INVx1_ASAP7_75t_L g106 ( .A(n_42), .Y(n_106) );
BUFx3_ASAP7_75t_L g492 ( .A(n_42), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_43), .A2(n_100), .B1(n_844), .B2(n_856), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_44), .B(n_600), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_46), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_47), .A2(n_83), .B1(n_140), .B2(n_198), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_49), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_50), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_53), .A2(n_77), .B1(n_172), .B2(n_548), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_54), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_55), .A2(n_81), .B1(n_143), .B2(n_170), .Y(n_522) );
INVx1_ASAP7_75t_L g126 ( .A(n_56), .Y(n_126) );
AND2x4_ASAP7_75t_L g146 ( .A(n_57), .B(n_147), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_58), .A2(n_88), .B1(n_198), .B2(n_228), .Y(n_227) );
AO22x1_ASAP7_75t_L g168 ( .A1(n_59), .A2(n_71), .B1(n_169), .B2(n_171), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_60), .B(n_143), .Y(n_510) );
INVx1_ASAP7_75t_L g147 ( .A(n_61), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_62), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_63), .B(n_149), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_64), .A2(n_160), .B(n_163), .C(n_568), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_65), .B(n_143), .C(n_515), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_67), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_68), .B(n_163), .Y(n_188) );
AND2x2_ASAP7_75t_L g570 ( .A(n_69), .B(n_221), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_70), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_72), .B(n_131), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_73), .A2(n_94), .B1(n_170), .B2(n_172), .Y(n_550) );
INVx2_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_75), .B(n_183), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_76), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_78), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_79), .B(n_149), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_80), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_82), .B(n_124), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_85), .B(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_86), .A2(n_98), .B1(n_198), .B2(n_217), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_87), .B(n_548), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_90), .B(n_149), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_91), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g487 ( .A(n_91), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_92), .B(n_208), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_93), .A2(n_163), .B(n_200), .C(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g220 ( .A(n_95), .B(n_221), .Y(n_220) );
NAND2xp33_ASAP7_75t_L g186 ( .A(n_96), .B(n_187), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_97), .Y(n_531) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_110), .Y(n_100) );
AOI21x1_ASAP7_75t_L g111 ( .A1(n_101), .A2(n_112), .B(n_113), .Y(n_111) );
NOR2xp33_ASAP7_75t_SL g101 ( .A(n_102), .B(n_109), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_103), .Y(n_112) );
AND2x6_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_107), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_108), .B(n_492), .Y(n_843) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_475), .B(n_478), .Y(n_110) );
INVx1_ASAP7_75t_L g474 ( .A(n_115), .Y(n_474) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g482 ( .A(n_116), .Y(n_482) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_374), .Y(n_116) );
NAND3xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_276), .C(n_336), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_151), .B1(n_263), .B2(n_269), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g333 ( .A(n_120), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_120), .B(n_250), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_120), .B(n_296), .Y(n_444) );
AND2x2_ASAP7_75t_L g450 ( .A(n_120), .B(n_275), .Y(n_450) );
INVxp67_ASAP7_75t_L g455 ( .A(n_120), .Y(n_455) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g267 ( .A(n_121), .Y(n_267) );
AOI21x1_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .B(n_148), .Y(n_121) );
AO31x2_ASAP7_75t_L g225 ( .A1(n_122), .A2(n_226), .A3(n_232), .B(n_234), .Y(n_225) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_123), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g221 ( .A(n_123), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_123), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_123), .B(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_123), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g174 ( .A1(n_124), .A2(n_145), .B(n_166), .Y(n_174) );
INVx2_ASAP7_75t_L g201 ( .A(n_124), .Y(n_201) );
INVx2_ASAP7_75t_L g209 ( .A(n_124), .Y(n_209) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_125), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_139), .B(n_145), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B(n_136), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_131), .A2(n_217), .B1(n_564), .B2(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g581 ( .A(n_131), .Y(n_581) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g134 ( .A(n_132), .Y(n_134) );
INVx3_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
INVx2_ASAP7_75t_L g143 ( .A(n_132), .Y(n_143) );
INVx1_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
INVx1_ASAP7_75t_L g217 ( .A(n_132), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
INVx2_ASAP7_75t_L g231 ( .A(n_134), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g530 ( .A1(n_136), .A2(n_231), .B(n_531), .C(n_532), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_136), .A2(n_144), .B1(n_574), .B2(n_575), .Y(n_573) );
BUFx4f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_137), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g515 ( .A(n_137), .Y(n_515) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx8_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx2_ASAP7_75t_L g161 ( .A(n_138), .Y(n_161) );
INVx1_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
INVx4_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
INVx2_ASAP7_75t_SL g548 ( .A(n_143), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_144), .B(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_144), .A2(n_186), .B(n_188), .Y(n_185) );
INVx6_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_144), .A2(n_158), .B(n_168), .C(n_174), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_144), .A2(n_510), .B(n_511), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_144), .A2(n_196), .B1(n_522), .B2(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_145), .A2(n_562), .B(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx10_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
BUFx10_ASAP7_75t_L g202 ( .A(n_146), .Y(n_202) );
INVx1_ASAP7_75t_L g233 ( .A(n_146), .Y(n_233) );
AO31x2_ASAP7_75t_L g578 ( .A1(n_146), .A2(n_545), .A3(n_579), .B(n_583), .Y(n_578) );
NOR2x1_ASAP7_75t_L g189 ( .A(n_149), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g304 ( .A(n_149), .Y(n_304) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g261 ( .A(n_150), .B(n_191), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_150), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g528 ( .A(n_150), .Y(n_528) );
BUFx3_ASAP7_75t_L g545 ( .A(n_150), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_150), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_SL g592 ( .A(n_150), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_222), .B(n_236), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_192), .Y(n_153) );
INVx1_ASAP7_75t_L g371 ( .A(n_154), .Y(n_371) );
AND2x2_ASAP7_75t_L g400 ( .A(n_154), .B(n_362), .Y(n_400) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_175), .Y(n_154) );
AND2x2_ASAP7_75t_L g293 ( .A(n_155), .B(n_206), .Y(n_293) );
INVx1_ASAP7_75t_L g349 ( .A(n_155), .Y(n_349) );
AND2x2_ASAP7_75t_L g399 ( .A(n_155), .B(n_205), .Y(n_399) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g273 ( .A(n_156), .B(n_205), .Y(n_273) );
AND2x4_ASAP7_75t_L g418 ( .A(n_156), .B(n_206), .Y(n_418) );
AOI21x1_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_167), .B(n_173), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_166), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_159), .A2(n_259), .B(n_260), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_159), .A2(n_196), .B1(n_302), .B2(n_303), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_159), .A2(n_196), .B1(n_580), .B2(n_582), .Y(n_579) );
AOI21x1_ASAP7_75t_L g594 ( .A1(n_159), .A2(n_595), .B(n_596), .Y(n_594) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g184 ( .A(n_161), .Y(n_184) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_165), .B(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g600 ( .A(n_170), .Y(n_600) );
OAI21xp33_ASAP7_75t_SL g253 ( .A1(n_171), .A2(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_172), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx2_ASAP7_75t_L g343 ( .A(n_175), .Y(n_343) );
AND2x2_ASAP7_75t_L g412 ( .A(n_175), .B(n_206), .Y(n_412) );
AND2x2_ASAP7_75t_L g419 ( .A(n_175), .B(n_244), .Y(n_419) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
BUFx3_ASAP7_75t_L g275 ( .A(n_176), .Y(n_275) );
AND2x2_ASAP7_75t_L g286 ( .A(n_176), .B(n_272), .Y(n_286) );
AND2x2_ASAP7_75t_L g350 ( .A(n_176), .B(n_193), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_176), .B(n_206), .Y(n_355) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
OAI21x1_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_185), .B(n_189), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_183), .Y(n_179) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_184), .A2(n_534), .B1(n_535), .B2(n_536), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g215 ( .A1(n_187), .A2(n_216), .B1(n_217), .B2(n_218), .Y(n_215) );
INVx2_ASAP7_75t_L g228 ( .A(n_187), .Y(n_228) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AO31x2_ASAP7_75t_L g300 ( .A1(n_191), .A2(n_301), .A3(n_304), .B(n_305), .Y(n_300) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_191), .A2(n_509), .B(n_512), .Y(n_508) );
AOI31xp67_ASAP7_75t_L g520 ( .A1(n_191), .A2(n_304), .A3(n_521), .B(n_524), .Y(n_520) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_191), .A2(n_530), .B(n_533), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_192), .B(n_361), .Y(n_463) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_205), .Y(n_192) );
INVx2_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
OR2x2_ASAP7_75t_L g247 ( .A(n_193), .B(n_206), .Y(n_247) );
INVx2_ASAP7_75t_L g272 ( .A(n_193), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_193), .B(n_242), .Y(n_288) );
AND2x2_ASAP7_75t_L g362 ( .A(n_193), .B(n_206), .Y(n_362) );
AO31x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_201), .A3(n_202), .B(n_203), .Y(n_193) );
OAI22x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_199), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_196), .A2(n_199), .B1(n_227), .B2(n_229), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_196), .A2(n_547), .B1(n_549), .B2(n_550), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_196), .A2(n_598), .B(n_599), .Y(n_597) );
INVx2_ASAP7_75t_L g230 ( .A(n_198), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_198), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g513 ( .A(n_198), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_199), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_SL g549 ( .A(n_200), .Y(n_549) );
INVx1_ASAP7_75t_L g566 ( .A(n_200), .Y(n_566) );
INVx2_ASAP7_75t_L g507 ( .A(n_201), .Y(n_507) );
INVx2_ASAP7_75t_L g219 ( .A(n_202), .Y(n_219) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g289 ( .A(n_206), .Y(n_289) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_210), .B(n_220), .Y(n_206) );
AOI21x1_ASAP7_75t_L g560 ( .A1(n_207), .A2(n_561), .B(n_570), .Y(n_560) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_219), .Y(n_210) );
INVx1_ASAP7_75t_L g535 ( .A(n_217), .Y(n_535) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_223), .B(n_325), .Y(n_471) );
BUFx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g262 ( .A(n_225), .Y(n_262) );
AND2x2_ASAP7_75t_L g268 ( .A(n_225), .B(n_250), .Y(n_268) );
INVx1_ASAP7_75t_L g317 ( .A(n_225), .Y(n_317) );
OR2x2_ASAP7_75t_L g322 ( .A(n_225), .B(n_300), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_225), .B(n_300), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_225), .B(n_299), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_225), .B(n_267), .Y(n_407) );
AO31x2_ASAP7_75t_L g544 ( .A1(n_232), .A2(n_545), .A3(n_546), .B(n_551), .Y(n_544) );
INVx2_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_SL g576 ( .A(n_233), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_245), .B(n_248), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
OR2x2_ASAP7_75t_L g246 ( .A(n_239), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g398 ( .A(n_239), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g428 ( .A(n_239), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_240), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g396 ( .A(n_240), .Y(n_396) );
OR2x2_ASAP7_75t_L g309 ( .A(n_241), .B(n_310), .Y(n_309) );
INVxp33_ASAP7_75t_L g427 ( .A(n_241), .Y(n_427) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
INVx2_ASAP7_75t_L g331 ( .A(n_242), .Y(n_331) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g284 ( .A(n_244), .Y(n_284) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_246), .A2(n_318), .B1(n_323), .B2(n_394), .C(n_397), .Y(n_393) );
OR2x2_ASAP7_75t_L g380 ( .A(n_247), .B(n_331), .Y(n_380) );
INVx2_ASAP7_75t_L g429 ( .A(n_247), .Y(n_429) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g329 ( .A(n_249), .Y(n_329) );
OR2x2_ASAP7_75t_L g332 ( .A(n_249), .B(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_249), .Y(n_373) );
OR2x2_ASAP7_75t_L g386 ( .A(n_249), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_262), .Y(n_249) );
NAND2x1p5_ASAP7_75t_SL g281 ( .A(n_250), .B(n_266), .Y(n_281) );
INVx3_ASAP7_75t_L g296 ( .A(n_250), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_250), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
AND2x2_ASAP7_75t_L g401 ( .A(n_250), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g408 ( .A(n_250), .B(n_315), .Y(n_408) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_258), .B(n_261), .Y(n_252) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
AND2x2_ASAP7_75t_L g460 ( .A(n_264), .B(n_319), .Y(n_460) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g364 ( .A(n_266), .B(n_334), .Y(n_364) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g298 ( .A(n_267), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g325 ( .A(n_267), .B(n_300), .Y(n_325) );
AND2x4_ASAP7_75t_L g422 ( .A(n_268), .B(n_392), .Y(n_422) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g341 ( .A(n_273), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_274), .B(n_362), .Y(n_446) );
AND2x2_ASAP7_75t_L g453 ( .A(n_274), .B(n_413), .Y(n_453) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g378 ( .A(n_275), .Y(n_378) );
AOI321xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_290), .A3(n_307), .B1(n_308), .B2(n_311), .C(n_326), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_278), .B(n_287), .Y(n_277) );
AOI21xp33_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_283), .B(n_285), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI21xp33_ASAP7_75t_L g290 ( .A1(n_280), .A2(n_291), .B(n_294), .Y(n_290) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
OR2x2_ASAP7_75t_L g390 ( .A(n_281), .B(n_322), .Y(n_390) );
INVx1_ASAP7_75t_L g382 ( .A(n_282), .Y(n_382) );
INVx2_ASAP7_75t_L g367 ( .A(n_283), .Y(n_367) );
OAI32xp33_ASAP7_75t_L g470 ( .A1(n_283), .A2(n_432), .A3(n_443), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g385 ( .A(n_284), .Y(n_385) );
INVx1_ASAP7_75t_L g335 ( .A(n_285), .Y(n_335) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_SL g423 ( .A(n_286), .B(n_330), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_287), .B(n_291), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_287), .A2(n_364), .B1(n_425), .B2(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g413 ( .A(n_288), .Y(n_413) );
INVx1_ASAP7_75t_L g310 ( .A(n_289), .Y(n_310) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g395 ( .A(n_293), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g311 ( .A(n_294), .B(n_312), .C(n_318), .D(n_323), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVxp67_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
AND2x2_ASAP7_75t_L g416 ( .A(n_295), .B(n_325), .Y(n_416) );
OR2x2_ASAP7_75t_L g425 ( .A(n_295), .B(n_298), .Y(n_425) );
AND2x2_ASAP7_75t_L g449 ( .A(n_295), .B(n_321), .Y(n_449) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g363 ( .A(n_296), .B(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g370 ( .A(n_296), .B(n_317), .Y(n_370) );
INVx1_ASAP7_75t_L g434 ( .A(n_297), .Y(n_434) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g342 ( .A(n_298), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g392 ( .A(n_298), .Y(n_392) );
INVx1_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g315 ( .A(n_300), .Y(n_315) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AND2x4_ASAP7_75t_L g328 ( .A(n_314), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_316), .Y(n_433) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g324 ( .A(n_320), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g410 ( .A(n_322), .Y(n_410) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g387 ( .A(n_325), .Y(n_387) );
AND2x2_ASAP7_75t_L g430 ( .A(n_325), .B(n_370), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_330), .B(n_332), .C(n_335), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g441 ( .A(n_330), .B(n_419), .Y(n_441) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g345 ( .A(n_333), .Y(n_345) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_351), .C(n_365), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_340), .A2(n_448), .B(n_451), .Y(n_447) );
INVx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g361 ( .A(n_343), .Y(n_361) );
AND2x2_ASAP7_75t_L g421 ( .A(n_343), .B(n_418), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g440 ( .A(n_348), .Y(n_440) );
AND2x2_ASAP7_75t_L g466 ( .A(n_348), .B(n_429), .Y(n_466) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g354 ( .A(n_349), .Y(n_354) );
INVx2_ASAP7_75t_L g405 ( .A(n_350), .Y(n_405) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_350), .B(n_440), .Y(n_439) );
AOI33xp33_ASAP7_75t_L g457 ( .A1(n_350), .A2(n_370), .A3(n_408), .B1(n_418), .B2(n_450), .B3(n_858), .Y(n_457) );
OAI22xp33_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_356), .B1(n_359), .B2(n_363), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
AND2x2_ASAP7_75t_L g384 ( .A(n_355), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_356), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g469 ( .A(n_358), .B(n_403), .Y(n_469) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
OAI22xp33_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_368), .B1(n_371), .B2(n_372), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_369), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_369), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g391 ( .A(n_370), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g456 ( .A(n_370), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_435), .Y(n_374) );
NOR4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_393), .C(n_414), .D(n_431), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_383), .B2(n_386), .C(n_388), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_SL g431 ( .A1(n_377), .A2(n_432), .B(n_433), .C(n_434), .Y(n_431) );
NAND2x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g464 ( .A(n_380), .Y(n_464) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_384), .A2(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x6_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
O2A1O1Ixp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_401), .C(n_404), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g443 ( .A(n_403), .B(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_403), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_409), .B2(n_411), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
OAI211xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B(n_420), .C(n_426), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_418), .A2(n_466), .B1(n_467), .B2(n_468), .C(n_470), .Y(n_465) );
INVx3_ASAP7_75t_L g473 ( .A(n_418), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_420) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g432 ( .A(n_429), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_458), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_447), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B(n_442), .C(n_445), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_441), .B(n_462), .C(n_464), .Y(n_461) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B(n_457), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_461), .B(n_465), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_SL g489 ( .A(n_476), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_477), .B(n_841), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_483), .B1(n_493), .B2(n_833), .C(n_836), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NOR2xp67_ASAP7_75t_SL g483 ( .A(n_484), .B(n_488), .Y(n_483) );
INVx4_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g842 ( .A(n_486), .B(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g835 ( .A(n_487), .Y(n_835) );
NOR2x1_ASAP7_75t_R g833 ( .A(n_488), .B(n_834), .Y(n_833) );
INVx5_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NOR3x1_ASAP7_75t_L g852 ( .A(n_492), .B(n_835), .C(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_496), .Y(n_832) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_741), .Y(n_496) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_498), .B(n_646), .C(n_673), .D(n_709), .Y(n_497) );
AOI221x1_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_557), .B1(n_585), .B2(n_621), .C(n_625), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_538), .C(n_555), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_518), .Y(n_502) );
INVx2_ASAP7_75t_L g586 ( .A(n_503), .Y(n_586) );
AND2x2_ASAP7_75t_L g759 ( .A(n_503), .B(n_703), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_503), .B(n_556), .Y(n_768) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g774 ( .A(n_504), .Y(n_774) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g619 ( .A(n_505), .Y(n_619) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g702 ( .A(n_506), .B(n_554), .Y(n_702) );
OAI21x1_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_517), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g631 ( .A1(n_507), .A2(n_508), .B(n_517), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_516), .Y(n_512) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_518), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_518), .B(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g772 ( .A(n_518), .Y(n_772) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
AND2x2_ASAP7_75t_L g556 ( .A(n_519), .B(n_544), .Y(n_556) );
INVx2_ASAP7_75t_L g628 ( .A(n_519), .Y(n_628) );
AND2x2_ASAP7_75t_L g693 ( .A(n_519), .B(n_631), .Y(n_693) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g620 ( .A(n_527), .Y(n_620) );
AND2x2_ASAP7_75t_L g630 ( .A(n_527), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g692 ( .A(n_527), .B(n_544), .Y(n_692) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .B(n_537), .Y(n_527) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_528), .A2(n_529), .B(n_537), .Y(n_541) );
INVx1_ASAP7_75t_L g657 ( .A(n_538), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_540), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_540), .B(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_540), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_540), .B(n_727), .Y(n_734) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g703 ( .A(n_541), .B(n_678), .Y(n_703) );
OR2x2_ASAP7_75t_L g705 ( .A(n_541), .B(n_631), .Y(n_705) );
INVx1_ASAP7_75t_L g764 ( .A(n_541), .Y(n_764) );
BUFx2_ASAP7_75t_L g778 ( .A(n_541), .Y(n_778) );
OR2x2_ASAP7_75t_L g806 ( .A(n_541), .B(n_544), .Y(n_806) );
INVx1_ASAP7_75t_L g825 ( .A(n_542), .Y(n_825) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g672 ( .A(n_543), .Y(n_672) );
OR2x2_ASAP7_75t_L g685 ( .A(n_543), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g704 ( .A(n_543), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_553), .Y(n_543) );
INVx2_ASAP7_75t_L g624 ( .A(n_544), .Y(n_624) );
AND2x2_ASAP7_75t_L g640 ( .A(n_544), .B(n_553), .Y(n_640) );
INVx1_ASAP7_75t_L g678 ( .A(n_544), .Y(n_678) );
INVx1_ASAP7_75t_L g721 ( .A(n_544), .Y(n_721) );
AND2x2_ASAP7_75t_L g763 ( .A(n_544), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g819 ( .A(n_555), .Y(n_819) );
AND2x4_ASAP7_75t_L g757 ( .A(n_556), .B(n_617), .Y(n_757) );
INVx2_ASAP7_75t_L g786 ( .A(n_556), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_556), .B(n_778), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_557), .B(n_776), .Y(n_775) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_571), .Y(n_557) );
AND2x2_ASAP7_75t_L g697 ( .A(n_558), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g718 ( .A(n_558), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g589 ( .A(n_559), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g613 ( .A(n_559), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g644 ( .A(n_559), .Y(n_644) );
AND2x2_ASAP7_75t_L g684 ( .A(n_559), .B(n_577), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_559), .B(n_668), .Y(n_725) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g637 ( .A(n_560), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_563), .B(n_566), .Y(n_562) );
INVx3_ASAP7_75t_L g603 ( .A(n_571), .Y(n_603) );
AND2x2_ASAP7_75t_L g648 ( .A(n_571), .B(n_643), .Y(n_648) );
AND2x2_ASAP7_75t_L g803 ( .A(n_571), .B(n_607), .Y(n_803) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g654 ( .A(n_572), .Y(n_654) );
AND2x2_ASAP7_75t_L g682 ( .A(n_572), .B(n_590), .Y(n_682) );
OAI21x1_ASAP7_75t_L g593 ( .A1(n_576), .A2(n_594), .B(n_597), .Y(n_593) );
AND2x4_ASAP7_75t_L g635 ( .A(n_577), .B(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g608 ( .A(n_578), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g645 ( .A(n_578), .B(n_609), .Y(n_645) );
AND2x2_ASAP7_75t_L g655 ( .A(n_578), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_578), .B(n_590), .Y(n_707) );
AND2x2_ASAP7_75t_L g713 ( .A(n_578), .B(n_637), .Y(n_713) );
OAI21xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_604), .Y(n_585) );
OAI21xp33_ASAP7_75t_L g746 ( .A1(n_586), .A2(n_747), .B(n_751), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_586), .B(n_777), .Y(n_824) );
NAND2x1_ASAP7_75t_SL g587 ( .A(n_588), .B(n_602), .Y(n_587) );
INVx1_ASAP7_75t_L g830 ( .A(n_588), .Y(n_830) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g607 ( .A(n_590), .Y(n_607) );
INVx2_ASAP7_75t_L g612 ( .A(n_590), .Y(n_612) );
INVxp67_ASAP7_75t_L g633 ( .A(n_590), .Y(n_633) );
AND2x2_ASAP7_75t_L g653 ( .A(n_590), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g664 ( .A(n_590), .B(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g668 ( .A(n_590), .Y(n_668) );
INVx1_ASAP7_75t_L g686 ( .A(n_590), .Y(n_686) );
OR2x2_ASAP7_75t_L g719 ( .A(n_590), .B(n_654), .Y(n_719) );
INVx1_ASAP7_75t_L g790 ( .A(n_590), .Y(n_790) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_601), .Y(n_591) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_610), .B(n_615), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_606), .A2(n_729), .B1(n_731), .B2(n_734), .Y(n_728) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_607), .B(n_655), .Y(n_689) );
BUFx2_ASAP7_75t_L g748 ( .A(n_607), .Y(n_748) );
INVx2_ASAP7_75t_L g698 ( .A(n_608), .Y(n_698) );
OR2x2_ASAP7_75t_L g782 ( .A(n_608), .B(n_612), .Y(n_782) );
INVx1_ASAP7_75t_L g614 ( .A(n_609), .Y(n_614) );
INVx1_ASAP7_75t_L g663 ( .A(n_609), .Y(n_663) );
NOR2x1p5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_612), .Y(n_733) );
OR2x2_ASAP7_75t_L g817 ( .A(n_612), .B(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g820 ( .A(n_612), .B(n_655), .Y(n_820) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_613), .Y(n_783) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_617), .B(n_677), .Y(n_739) );
AND2x2_ASAP7_75t_L g829 ( .A(n_617), .B(n_627), .Y(n_829) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g738 ( .A(n_618), .B(n_627), .Y(n_738) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AND2x2_ASAP7_75t_L g695 ( .A(n_619), .B(n_628), .Y(n_695) );
AND2x2_ASAP7_75t_L g730 ( .A(n_619), .B(n_624), .Y(n_730) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g649 ( .A(n_622), .B(n_630), .Y(n_649) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g789 ( .A(n_624), .B(n_790), .Y(n_789) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_632), .B1(n_638), .B2(n_641), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g826 ( .A1(n_626), .A2(n_827), .B(n_828), .C(n_830), .Y(n_826) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g677 ( .A(n_628), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g745 ( .A(n_628), .Y(n_745) );
OR2x2_ASAP7_75t_L g792 ( .A(n_629), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
AND2x2_ASAP7_75t_L g647 ( .A(n_633), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g750 ( .A(n_636), .Y(n_750) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g656 ( .A(n_637), .Y(n_656) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_637), .Y(n_665) );
INVx1_ASAP7_75t_L g737 ( .A(n_637), .Y(n_737) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g793 ( .A(n_640), .Y(n_793) );
AND2x2_ASAP7_75t_L g815 ( .A(n_640), .B(n_778), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_641), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g667 ( .A(n_645), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g723 ( .A(n_645), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g818 ( .A(n_645), .Y(n_818) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_650), .B2(n_657), .C(n_658), .Y(n_646) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx2_ASAP7_75t_L g740 ( .A(n_653), .Y(n_740) );
BUFx2_ASAP7_75t_L g760 ( .A(n_655), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_666), .B(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .Y(n_660) );
AND2x2_ASAP7_75t_L g802 ( .A(n_661), .B(n_724), .Y(n_802) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g708 ( .A(n_663), .Y(n_708) );
AND2x2_ASAP7_75t_L g798 ( .A(n_663), .B(n_668), .Y(n_798) );
INVx1_ASAP7_75t_L g681 ( .A(n_665), .Y(n_681) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_687), .C(n_699), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B1(n_683), .B2(n_685), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
BUFx2_ASAP7_75t_L g715 ( .A(n_682), .Y(n_715) );
AND2x2_ASAP7_75t_L g808 ( .A(n_682), .B(n_750), .Y(n_808) );
OAI21xp33_ASAP7_75t_L g811 ( .A1(n_683), .A2(n_812), .B(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B1(n_694), .B2(n_696), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_690), .B(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g762 ( .A(n_695), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g749 ( .A(n_698), .B(n_750), .Y(n_749) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_698), .Y(n_765) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B(n_706), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
AND2x2_ASAP7_75t_L g776 ( .A(n_701), .B(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g813 ( .A(n_701), .B(n_778), .Y(n_813) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g727 ( .A(n_702), .Y(n_727) );
OR2x2_ASAP7_75t_L g805 ( .A(n_702), .B(n_806), .Y(n_805) );
OR2x2_ASAP7_75t_L g720 ( .A(n_705), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g752 ( .A(n_705), .Y(n_752) );
OR2x2_ASAP7_75t_L g785 ( .A(n_705), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g756 ( .A(n_706), .Y(n_756) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_728), .C(n_735), .Y(n_709) );
OAI322xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_714), .A3(n_716), .B1(n_718), .B2(n_720), .C1(n_722), .C2(n_726), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g787 ( .A1(n_712), .A2(n_752), .B(n_788), .C(n_791), .Y(n_787) );
BUFx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g732 ( .A(n_713), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g769 ( .A(n_713), .Y(n_769) );
AND2x4_ASAP7_75t_L g797 ( .A(n_713), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI32xp33_ASAP7_75t_L g766 ( .A1(n_715), .A2(n_753), .A3(n_767), .B1(n_769), .B2(n_770), .Y(n_766) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g753 ( .A(n_719), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_721), .B(n_774), .Y(n_773) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
O2A1O1Ixp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B(n_739), .C(n_740), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_742), .B(n_799), .Y(n_741) );
AOI211xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B(n_754), .C(n_779), .Y(n_742) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_SL g821 ( .A1(n_747), .A2(n_822), .B(n_823), .C(n_825), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
OAI31xp33_ASAP7_75t_L g801 ( .A1(n_749), .A2(n_802), .A3(n_803), .B(n_804), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g761 ( .A(n_753), .Y(n_761) );
NAND4xp25_ASAP7_75t_SL g754 ( .A(n_755), .B(n_758), .C(n_766), .D(n_775), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
AOI32xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .A3(n_761), .B1(n_762), .B2(n_765), .Y(n_758) );
INVx1_ASAP7_75t_L g810 ( .A(n_762), .Y(n_810) );
INVx1_ASAP7_75t_L g822 ( .A(n_765), .Y(n_822) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OR2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_787), .C(n_794), .Y(n_779) );
OAI21xp5_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_783), .B(n_784), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx3_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_SL g812 ( .A(n_788), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NOR4xp25_ASAP7_75t_L g799 ( .A(n_800), .B(n_811), .C(n_821), .D(n_826), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_807), .Y(n_800) );
OAI21xp33_ASAP7_75t_L g807 ( .A1(n_802), .A2(n_808), .B(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_819), .B2(n_820), .Y(n_814) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_818), .Y(n_827) );
INVxp67_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx6f_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx6_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
BUFx10_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx4f_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx8_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx8_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_847), .Y(n_856) );
AND2x6_ASAP7_75t_L g847 ( .A(n_848), .B(n_852), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
INVx2_ASAP7_75t_SL g853 ( .A(n_854), .Y(n_853) );
endmodule