module fake_ariane_3069_n_1354 (n_295, n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_289, n_288, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_294, n_47, n_110, n_304, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_299, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_281, n_209, n_49, n_262, n_291, n_20, n_292, n_174, n_275, n_100, n_305, n_17, n_283, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_297, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_290, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_286, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_287, n_302, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_284, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_282, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_301, n_184, n_177, n_135, n_258, n_73, n_77, n_293, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_303, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_279, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_280, n_215, n_252, n_142, n_251, n_161, n_285, n_300, n_14, n_163, n_88, n_186, n_141, n_296, n_298, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1354);

input n_295;
input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_289;
input n_288;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_294;
input n_47;
input n_110;
input n_304;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_299;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_281;
input n_209;
input n_49;
input n_262;
input n_291;
input n_20;
input n_292;
input n_174;
input n_275;
input n_100;
input n_305;
input n_17;
input n_283;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_297;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_290;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_286;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_287;
input n_302;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_284;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_282;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_301;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_293;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_303;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_279;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_280;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_285;
input n_300;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_296;
input n_298;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1354;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1341;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_222),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_180),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_170),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_46),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_300),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_101),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_286),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_103),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_132),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_236),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_261),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_247),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_107),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_40),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_111),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_279),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_17),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_302),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_93),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_189),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_96),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_79),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_223),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_242),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_268),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_46),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_262),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_144),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_159),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_243),
.Y(n_337)
);

BUFx2_ASAP7_75t_R g338 ( 
.A(n_177),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_39),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_229),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_40),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_259),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_190),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_125),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_15),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_16),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_166),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_109),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_130),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_272),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_42),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_246),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_209),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_44),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_257),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_34),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_27),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_292),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_290),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_171),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_120),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_24),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_75),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_219),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_182),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_287),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_32),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_283),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_207),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_136),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_117),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_49),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_258),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_25),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_16),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_4),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_291),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_56),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_151),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_285),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_17),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_244),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_217),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_12),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_212),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_34),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_206),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_43),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_13),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_274),
.Y(n_390)
);

INVx4_ASAP7_75t_R g391 ( 
.A(n_23),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_239),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_80),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_226),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_30),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_255),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_167),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_240),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_77),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_245),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_24),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_188),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_138),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_79),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_227),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_104),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_158),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_264),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_41),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_225),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_234),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_168),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_208),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_121),
.Y(n_414)
);

BUFx10_ASAP7_75t_L g415 ( 
.A(n_6),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_175),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_216),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_275),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_76),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_124),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_237),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_69),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_127),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_105),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_67),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_87),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_253),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_71),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_281),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_25),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_9),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_66),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_81),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_60),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_29),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_211),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_295),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_22),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_174),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_298),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_85),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_94),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_238),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_39),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_80),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_230),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_224),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_202),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_181),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_143),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_92),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_256),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_232),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_164),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_187),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_270),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_172),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_102),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_59),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_195),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_65),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_169),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_278),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_135),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_152),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_178),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_186),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_131),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_173),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_288),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_6),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_299),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_241),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_148),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_64),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_63),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_210),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_215),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_150),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_97),
.Y(n_480)
);

BUFx5_ASAP7_75t_L g481 ( 
.A(n_45),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_54),
.Y(n_482)
);

BUFx5_ASAP7_75t_L g483 ( 
.A(n_20),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_199),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_89),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_139),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_198),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_303),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_7),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_265),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_147),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_7),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_157),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_31),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_140),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_137),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_191),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_304),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_2),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_75),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_266),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_231),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_33),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_115),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_213),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_45),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_254),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_252),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_194),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g510 ( 
.A(n_145),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_42),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_192),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_28),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_337),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_0),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_0),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_337),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_337),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_315),
.B(n_1),
.Y(n_521)
);

CKINVDCx6p67_ASAP7_75t_R g522 ( 
.A(n_309),
.Y(n_522)
);

INVx6_ASAP7_75t_L g523 ( 
.A(n_417),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_337),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_481),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_481),
.B(n_1),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_321),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_374),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_374),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_345),
.B(n_2),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_496),
.B(n_3),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_336),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_437),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_327),
.B(n_3),
.Y(n_534)
);

BUFx8_ASAP7_75t_SL g535 ( 
.A(n_432),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_329),
.B(n_4),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_437),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_336),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_481),
.B(n_5),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_481),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_372),
.B(n_5),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_333),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_339),
.Y(n_544)
);

BUFx12f_ASAP7_75t_L g545 ( 
.A(n_372),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_348),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_360),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_372),
.B(n_415),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_360),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_450),
.Y(n_550)
);

BUFx12f_ASAP7_75t_L g551 ( 
.A(n_415),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_450),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_328),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_481),
.B(n_8),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_483),
.B(n_8),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_483),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_354),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_330),
.B(n_9),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_415),
.B(n_10),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_483),
.B(n_10),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_335),
.B(n_11),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_343),
.B(n_347),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_345),
.B(n_11),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_398),
.Y(n_564)
);

BUFx8_ASAP7_75t_L g565 ( 
.A(n_436),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_362),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_483),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_354),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_369),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_362),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_483),
.B(n_13),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_354),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_354),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_483),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_388),
.B(n_14),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_388),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_324),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_422),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_356),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_311),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_379),
.B(n_14),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_422),
.B(n_15),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_341),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_489),
.B(n_18),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_392),
.B(n_18),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_489),
.B(n_19),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_357),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_311),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_403),
.B(n_19),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_319),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_410),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_319),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_320),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_376),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_412),
.B(n_20),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_378),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_381),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_320),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_351),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_426),
.B(n_433),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_340),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_340),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_384),
.B(n_21),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_463),
.B(n_21),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_361),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_439),
.B(n_22),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_389),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_399),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_441),
.B(n_23),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_463),
.B(n_26),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_443),
.B(n_27),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_314),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_508),
.B(n_29),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_404),
.B(n_30),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_449),
.B(n_31),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_332),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_361),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_430),
.B(n_32),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_364),
.Y(n_620)
);

BUFx12f_ASAP7_75t_L g621 ( 
.A(n_363),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_364),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_476),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_451),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_508),
.B(n_510),
.Y(n_625)
);

BUFx8_ASAP7_75t_SL g626 ( 
.A(n_432),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_455),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_396),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_396),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_418),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_482),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_500),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_418),
.B(n_446),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_511),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_367),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_375),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_513),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_510),
.B(n_33),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_458),
.B(n_462),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_446),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_467),
.B(n_35),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_467),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_464),
.B(n_35),
.Y(n_643)
);

BUFx12f_ASAP7_75t_L g644 ( 
.A(n_386),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_306),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_491),
.B(n_36),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_493),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_307),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_308),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_495),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_498),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_504),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_505),
.B(n_36),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_393),
.B(n_37),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_401),
.B(n_37),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_310),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_444),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_507),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_509),
.B(n_38),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_411),
.B(n_38),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_395),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_409),
.B(n_41),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_313),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_424),
.B(n_43),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_316),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_469),
.B(n_44),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_338),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_605),
.A2(n_331),
.B1(n_484),
.B2(n_465),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_523),
.B(n_548),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_545),
.B(n_346),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_593),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_611),
.A2(n_331),
.B1(n_484),
.B2(n_465),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_531),
.A2(n_428),
.B1(n_431),
.B2(n_425),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_L g675 ( 
.A1(n_522),
.A2(n_419),
.B1(n_368),
.B2(n_390),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_557),
.Y(n_676)
);

NAND3x1_ASAP7_75t_L g677 ( 
.A(n_536),
.B(n_391),
.C(n_387),
.Y(n_677)
);

NAND3x1_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_427),
.C(n_408),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_593),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_568),
.Y(n_680)
);

AO22x2_ASAP7_75t_L g681 ( 
.A1(n_531),
.A2(n_473),
.B1(n_312),
.B2(n_421),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_568),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_568),
.Y(n_683)
);

OA22x2_ASAP7_75t_L g684 ( 
.A1(n_658),
.A2(n_435),
.B1(n_438),
.B2(n_434),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_613),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_614),
.A2(n_486),
.B1(n_459),
.B2(n_461),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_SL g687 ( 
.A1(n_617),
.A2(n_471),
.B1(n_475),
.B2(n_445),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_542),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_523),
.B(n_518),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_572),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_572),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_572),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_638),
.A2(n_494),
.B1(n_499),
.B2(n_492),
.Y(n_693)
);

AO22x1_ASAP7_75t_L g694 ( 
.A1(n_641),
.A2(n_506),
.B1(n_503),
.B2(n_318),
.Y(n_694)
);

AOI22x1_ASAP7_75t_L g695 ( 
.A1(n_641),
.A2(n_322),
.B1(n_323),
.B2(n_317),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_SL g696 ( 
.A1(n_655),
.A2(n_663),
.B1(n_523),
.B2(n_515),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_573),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_SL g698 ( 
.A1(n_655),
.A2(n_326),
.B1(n_334),
.B2(n_325),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_593),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_573),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_535),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_515),
.A2(n_344),
.B1(n_349),
.B2(n_342),
.Y(n_702)
);

OAI22xp33_ASAP7_75t_L g703 ( 
.A1(n_662),
.A2(n_352),
.B1(n_353),
.B2(n_350),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_532),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_662),
.A2(n_358),
.B1(n_359),
.B2(n_355),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_551),
.B(n_519),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_533),
.B(n_537),
.Y(n_707)
);

AO22x2_ASAP7_75t_L g708 ( 
.A1(n_559),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_708)
);

AO22x2_ASAP7_75t_L g709 ( 
.A1(n_530),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_656),
.A2(n_544),
.B1(n_600),
.B2(n_584),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_594),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_665),
.A2(n_366),
.B1(n_370),
.B2(n_365),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_532),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_635),
.A2(n_636),
.B1(n_654),
.B2(n_562),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_654),
.A2(n_562),
.B1(n_661),
.B2(n_563),
.Y(n_715)
);

AO22x2_ASAP7_75t_L g716 ( 
.A1(n_530),
.A2(n_563),
.B1(n_585),
.B2(n_575),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_665),
.A2(n_373),
.B1(n_377),
.B2(n_371),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_667),
.A2(n_382),
.B1(n_383),
.B2(n_380),
.Y(n_718)
);

AO22x2_ASAP7_75t_L g719 ( 
.A1(n_575),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_719)
);

OAI22x1_ASAP7_75t_L g720 ( 
.A1(n_626),
.A2(n_587),
.B1(n_585),
.B2(n_604),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_533),
.B(n_385),
.Y(n_721)
);

AO22x2_ASAP7_75t_L g722 ( 
.A1(n_587),
.A2(n_604),
.B1(n_619),
.B2(n_615),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_573),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_525),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_517),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_537),
.B(n_394),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_661),
.A2(n_400),
.B1(n_402),
.B2(n_397),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_667),
.A2(n_406),
.B1(n_407),
.B2(n_405),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_SL g729 ( 
.A1(n_608),
.A2(n_414),
.B1(n_416),
.B2(n_413),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_540),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_537),
.A2(n_512),
.B1(n_502),
.B2(n_501),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_532),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_615),
.A2(n_466),
.B1(n_490),
.B2(n_488),
.Y(n_733)
);

AND2x2_ASAP7_75t_SL g734 ( 
.A(n_583),
.B(n_619),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_R g735 ( 
.A1(n_521),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_735)
);

AO22x2_ASAP7_75t_L g736 ( 
.A1(n_601),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_621),
.A2(n_497),
.B1(n_487),
.B2(n_485),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_594),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_537),
.B(n_420),
.Y(n_739)
);

NAND3x1_ASAP7_75t_L g740 ( 
.A(n_582),
.B(n_55),
.C(n_57),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_543),
.B(n_423),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_601),
.A2(n_480),
.B1(n_479),
.B2(n_477),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_543),
.A2(n_474),
.B1(n_472),
.B2(n_468),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_528),
.B(n_429),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_528),
.B(n_440),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_582),
.B(n_442),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_556),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_594),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_529),
.B(n_447),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_538),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_599),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_664),
.B(n_448),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_552),
.B(n_452),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_599),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_666),
.B(n_453),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_590),
.A2(n_460),
.B1(n_457),
.B2(n_456),
.Y(n_756)
);

BUFx6f_ASAP7_75t_SL g757 ( 
.A(n_706),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_724),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_R g759 ( 
.A(n_668),
.B(n_595),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_730),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_755),
.B(n_546),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_747),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_676),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_670),
.B(n_546),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_685),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_672),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_746),
.B(n_734),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_689),
.Y(n_768)
);

XNOR2xp5_ASAP7_75t_L g769 ( 
.A(n_669),
.B(n_588),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_672),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_679),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_679),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_716),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_673),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_699),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_711),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_753),
.B(n_553),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_707),
.B(n_565),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_738),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_688),
.B(n_569),
.Y(n_780)
);

XNOR2x2_ASAP7_75t_L g781 ( 
.A(n_681),
.B(n_521),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_696),
.B(n_516),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_752),
.B(n_546),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_744),
.B(n_564),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_738),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_748),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_745),
.B(n_592),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_716),
.B(n_624),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_748),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_735),
.B(n_644),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_751),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_751),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_754),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_754),
.Y(n_794)
);

HAxp5_ASAP7_75t_SL g795 ( 
.A(n_735),
.B(n_578),
.CON(n_795),
.SN(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_704),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_713),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_732),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_722),
.B(n_627),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_750),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_750),
.Y(n_801)
);

XOR2xp5_ASAP7_75t_L g802 ( 
.A(n_687),
.B(n_527),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_710),
.B(n_527),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_722),
.B(n_714),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_680),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_682),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_686),
.B(n_659),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_749),
.A2(n_526),
.B(n_516),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_683),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_706),
.Y(n_810)
);

XOR2x2_ASAP7_75t_L g811 ( 
.A(n_678),
.B(n_639),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_715),
.B(n_566),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_693),
.B(n_566),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_701),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_690),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_691),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_692),
.Y(n_817)
);

AND2x6_ASAP7_75t_L g818 ( 
.A(n_721),
.B(n_526),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_697),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_700),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_723),
.Y(n_821)
);

XOR2x2_ASAP7_75t_L g822 ( 
.A(n_677),
.B(n_577),
.Y(n_822)
);

XNOR2xp5_ASAP7_75t_L g823 ( 
.A(n_675),
.B(n_577),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_725),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_725),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_684),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_733),
.B(n_564),
.Y(n_828)
);

NOR2x1p5_ASAP7_75t_L g829 ( 
.A(n_709),
.B(n_595),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_726),
.A2(n_567),
.B(n_574),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_698),
.B(n_539),
.Y(n_831)
);

BUFx6f_ASAP7_75t_SL g832 ( 
.A(n_671),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_739),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_727),
.B(n_538),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_741),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_721),
.Y(n_836)
);

AND2x2_ASAP7_75t_SL g837 ( 
.A(n_709),
.B(n_590),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_808),
.A2(n_702),
.B(n_695),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_767),
.A2(n_681),
.B1(n_719),
.B2(n_694),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_833),
.B(n_712),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_787),
.B(n_717),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_773),
.B(n_719),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_835),
.B(n_718),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_766),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_765),
.B(n_703),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_780),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_766),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_773),
.B(n_708),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_767),
.A2(n_708),
.B1(n_728),
.B2(n_756),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_799),
.Y(n_850)
);

AND2x2_ASAP7_75t_SL g851 ( 
.A(n_837),
.B(n_596),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_770),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_834),
.B(n_695),
.Y(n_853)
);

BUFx12f_ASAP7_75t_L g854 ( 
.A(n_814),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_830),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_760),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_812),
.B(n_608),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_760),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_768),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_770),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_788),
.B(n_646),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_834),
.B(n_705),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_772),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_772),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_764),
.B(n_731),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_837),
.B(n_596),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_789),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_789),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_777),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_758),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_807),
.B(n_648),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_813),
.B(n_652),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_762),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_777),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_771),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_829),
.B(n_653),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_782),
.A2(n_729),
.B1(n_674),
.B2(n_720),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_818),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_836),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_804),
.B(n_637),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_827),
.B(n_623),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_782),
.B(n_637),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_803),
.B(n_769),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_831),
.B(n_828),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_775),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_763),
.B(n_580),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_811),
.B(n_597),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_818),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_764),
.B(n_598),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_828),
.B(n_742),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_818),
.B(n_784),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_831),
.B(n_609),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_802),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_823),
.B(n_634),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_776),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_778),
.B(n_737),
.Y(n_896)
);

AND2x2_ASAP7_75t_SL g897 ( 
.A(n_781),
.B(n_610),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_779),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_784),
.B(n_743),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_759),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_816),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_785),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_816),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_759),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_R g905 ( 
.A(n_796),
.B(n_631),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_786),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_824),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_783),
.B(n_610),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_757),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_791),
.Y(n_910)
);

AND2x2_ASAP7_75t_SL g911 ( 
.A(n_795),
.B(n_616),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_792),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_795),
.B(n_616),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_793),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_783),
.B(n_660),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_794),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_822),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_797),
.B(n_632),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_822),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_810),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_817),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_817),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_876),
.B(n_798),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_847),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_854),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_876),
.B(n_800),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_856),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_869),
.B(n_874),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_869),
.B(n_801),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_844),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_847),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_858),
.B(n_790),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_857),
.B(n_774),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_884),
.B(n_761),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_854),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_844),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_888),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_888),
.Y(n_938)
);

AND2x6_ASAP7_75t_L g939 ( 
.A(n_878),
.B(n_819),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_860),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_857),
.B(n_774),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_883),
.B(n_671),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_860),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_920),
.B(n_757),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_859),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_871),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_852),
.Y(n_947)
);

BUFx12f_ASAP7_75t_L g948 ( 
.A(n_874),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_863),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_863),
.Y(n_950)
);

BUFx12f_ASAP7_75t_L g951 ( 
.A(n_881),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_880),
.B(n_805),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_856),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_871),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_880),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_862),
.B(n_761),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_894),
.B(n_570),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_864),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_894),
.B(n_579),
.Y(n_959)
);

INVx6_ASAP7_75t_L g960 ( 
.A(n_881),
.Y(n_960)
);

AND2x6_ASAP7_75t_L g961 ( 
.A(n_878),
.B(n_806),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_872),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_842),
.B(n_861),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_856),
.Y(n_964)
);

INVx4_ASAP7_75t_SL g965 ( 
.A(n_842),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_864),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_861),
.B(n_809),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_887),
.B(n_736),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_867),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_848),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_882),
.B(n_815),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_856),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_856),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_846),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_848),
.B(n_820),
.Y(n_975)
);

BUFx12f_ASAP7_75t_L g976 ( 
.A(n_881),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_858),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_879),
.B(n_821),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_868),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_900),
.B(n_660),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_904),
.B(n_534),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_867),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_886),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_891),
.B(n_825),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_882),
.B(n_576),
.Y(n_985)
);

NAND2x1_ASAP7_75t_SL g986 ( 
.A(n_845),
.B(n_839),
.Y(n_986)
);

INVx6_ASAP7_75t_L g987 ( 
.A(n_918),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_868),
.Y(n_988)
);

AND2x2_ASAP7_75t_SL g989 ( 
.A(n_911),
.B(n_832),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_879),
.B(n_826),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_921),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_908),
.B(n_633),
.Y(n_992)
);

BUFx8_ASAP7_75t_L g993 ( 
.A(n_887),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_889),
.B(n_534),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_988),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_945),
.Y(n_996)
);

BUFx12f_ASAP7_75t_L g997 ( 
.A(n_935),
.Y(n_997)
);

BUFx4_ASAP7_75t_SL g998 ( 
.A(n_925),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_961),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_944),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_963),
.Y(n_1001)
);

INVx6_ASAP7_75t_L g1002 ( 
.A(n_951),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_991),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_956),
.B(n_851),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_976),
.Y(n_1005)
);

INVx6_ASAP7_75t_L g1006 ( 
.A(n_948),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_944),
.Y(n_1007)
);

INVx5_ASAP7_75t_L g1008 ( 
.A(n_961),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_987),
.A2(n_911),
.B1(n_913),
.B2(n_897),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_988),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_968),
.A2(n_913),
.B1(n_897),
.B2(n_866),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_973),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_974),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_973),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_993),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_993),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_932),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_988),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_991),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_977),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_924),
.Y(n_1021)
);

CKINVDCx11_ASAP7_75t_R g1022 ( 
.A(n_977),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_989),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_927),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_934),
.B(n_851),
.Y(n_1025)
);

INVx6_ASAP7_75t_SL g1026 ( 
.A(n_975),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_937),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_950),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_987),
.A2(n_866),
.B1(n_849),
.B2(n_890),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_927),
.Y(n_1030)
);

BUFx24_ASAP7_75t_L g1031 ( 
.A(n_963),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_937),
.Y(n_1032)
);

CKINVDCx16_ASAP7_75t_R g1033 ( 
.A(n_933),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_924),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_983),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_960),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_960),
.Y(n_1037)
);

BUFx2_ASAP7_75t_SL g1038 ( 
.A(n_928),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_931),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_938),
.B(n_907),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_SL g1041 ( 
.A(n_955),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_962),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_942),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_927),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_941),
.B(n_850),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_934),
.A2(n_838),
.B1(n_915),
.B2(n_853),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_950),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_940),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_940),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_938),
.B(n_907),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_975),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_953),
.Y(n_1052)
);

OAI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1009),
.A2(n_877),
.B1(n_899),
.B2(n_917),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1011),
.A2(n_917),
.B1(n_919),
.B2(n_957),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_996),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1003),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_1045),
.B(n_970),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1019),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_1021),
.Y(n_1059)
);

OAI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1029),
.A2(n_994),
.B1(n_841),
.B2(n_865),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_1002),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1025),
.A2(n_898),
.B1(n_906),
.B2(n_875),
.Y(n_1062)
);

INVx6_ASAP7_75t_L g1063 ( 
.A(n_1002),
.Y(n_1063)
);

INVx6_ASAP7_75t_L g1064 ( 
.A(n_1017),
.Y(n_1064)
);

BUFx8_ASAP7_75t_L g1065 ( 
.A(n_1005),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_SL g1066 ( 
.A1(n_1033),
.A2(n_832),
.B1(n_893),
.B2(n_986),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_1022),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_1026),
.Y(n_1068)
);

INVx6_ASAP7_75t_L g1069 ( 
.A(n_1006),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_1038),
.Y(n_1070)
);

OAI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1025),
.A2(n_843),
.B1(n_840),
.B2(n_954),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_998),
.Y(n_1072)
);

BUFx12f_ASAP7_75t_L g1073 ( 
.A(n_997),
.Y(n_1073)
);

BUFx12f_ASAP7_75t_L g1074 ( 
.A(n_1006),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_998),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_1014),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1034),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_999),
.B(n_1008),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1011),
.A2(n_959),
.B1(n_946),
.B2(n_967),
.Y(n_1079)
);

INVx6_ASAP7_75t_L g1080 ( 
.A(n_1043),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_1014),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1004),
.B(n_943),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1039),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_1035),
.Y(n_1084)
);

INVx8_ASAP7_75t_L g1085 ( 
.A(n_1014),
.Y(n_1085)
);

BUFx8_ASAP7_75t_L g1086 ( 
.A(n_1015),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1028),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1048),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_1016),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1047),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1049),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1001),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1046),
.A2(n_992),
.B(n_985),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_1037),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1051),
.Y(n_1095)
);

OAI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1013),
.A2(n_980),
.B1(n_896),
.B2(n_981),
.Y(n_1096)
);

BUFx12f_ASAP7_75t_L g1097 ( 
.A(n_1000),
.Y(n_1097)
);

INVx8_ASAP7_75t_L g1098 ( 
.A(n_999),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1026),
.A2(n_952),
.B1(n_870),
.B2(n_1042),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1046),
.B(n_943),
.Y(n_1100)
);

BUFx8_ASAP7_75t_L g1101 ( 
.A(n_1007),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_1023),
.Y(n_1102)
);

INVx3_ASAP7_75t_SL g1103 ( 
.A(n_1020),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1013),
.A2(n_978),
.B1(n_990),
.B2(n_926),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1036),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1031),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_1072),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1053),
.A2(n_892),
.B1(n_870),
.B2(n_873),
.Y(n_1108)
);

OAI222xp33_ASAP7_75t_L g1109 ( 
.A1(n_1053),
.A2(n_1054),
.B1(n_1079),
.B2(n_1066),
.C1(n_1106),
.C2(n_1060),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1060),
.A2(n_892),
.B1(n_873),
.B2(n_885),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1059),
.A2(n_875),
.B1(n_906),
.B2(n_898),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1106),
.A2(n_1031),
.B1(n_1008),
.B2(n_999),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1056),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1059),
.A2(n_1041),
.B1(n_910),
.B2(n_916),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1094),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_1064),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1057),
.B(n_965),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1058),
.Y(n_1118)
);

OAI21xp33_ASAP7_75t_L g1119 ( 
.A1(n_1100),
.A2(n_561),
.B(n_558),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1077),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1104),
.A2(n_910),
.B1(n_916),
.B2(n_1008),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1100),
.A2(n_1008),
.B1(n_740),
.B2(n_971),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1071),
.B(n_889),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1096),
.A2(n_1012),
.B1(n_1032),
.B2(n_1027),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1070),
.A2(n_586),
.B1(n_607),
.B2(n_558),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1083),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_1062),
.A2(n_643),
.B(n_612),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1092),
.B(n_966),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1075),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1101),
.Y(n_1130)
);

BUFx4f_ASAP7_75t_L g1131 ( 
.A(n_1094),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1082),
.A2(n_647),
.B1(n_555),
.B2(n_560),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1087),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1093),
.A2(n_1010),
.B(n_995),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_SL g1135 ( 
.A1(n_1099),
.A2(n_571),
.B(n_554),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1082),
.A2(n_1091),
.B1(n_1088),
.B2(n_1093),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1090),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_SL g1138 ( 
.A1(n_1070),
.A2(n_984),
.B1(n_961),
.B2(n_939),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1055),
.B(n_923),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1089),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_1098),
.A2(n_984),
.B1(n_961),
.B2(n_939),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1055),
.B(n_926),
.Y(n_1142)
);

OAI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1067),
.A2(n_1012),
.B1(n_1050),
.B2(n_1040),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1094),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1095),
.Y(n_1145)
);

OAI222xp33_ASAP7_75t_L g1146 ( 
.A1(n_1105),
.A2(n_982),
.B1(n_969),
.B2(n_912),
.C1(n_914),
.C2(n_902),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1080),
.A2(n_895),
.B1(n_912),
.B2(n_902),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1102),
.A2(n_936),
.B1(n_947),
.B2(n_930),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1076),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1097),
.A2(n_958),
.B1(n_949),
.B2(n_985),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1084),
.B(n_909),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1103),
.B(n_918),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1068),
.A2(n_1050),
.B(n_1040),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1078),
.A2(n_1032),
.B(n_1027),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1076),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1069),
.A2(n_992),
.B1(n_979),
.B2(n_995),
.Y(n_1156)
);

BUFx8_ASAP7_75t_L g1157 ( 
.A(n_1073),
.Y(n_1157)
);

OAI211xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1119),
.A2(n_1081),
.B(n_905),
.C(n_1086),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1125),
.A2(n_1061),
.B1(n_1063),
.B2(n_1074),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1113),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1123),
.A2(n_549),
.B1(n_550),
.B2(n_547),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1118),
.B(n_1101),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1120),
.B(n_1126),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1137),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1127),
.B(n_651),
.C(n_1065),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1145),
.B(n_1065),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1150),
.A2(n_547),
.B1(n_868),
.B2(n_651),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1108),
.A2(n_868),
.B1(n_903),
.B2(n_901),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1121),
.A2(n_922),
.B1(n_903),
.B2(n_929),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1136),
.B(n_57),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1111),
.A2(n_1018),
.B(n_1024),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1136),
.B(n_1018),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_SL g1173 ( 
.A1(n_1122),
.A2(n_1085),
.B1(n_630),
.B2(n_602),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1122),
.A2(n_1148),
.B1(n_1133),
.B2(n_1142),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1114),
.A2(n_979),
.B1(n_964),
.B2(n_972),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1139),
.A2(n_922),
.B1(n_629),
.B2(n_620),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1115),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1110),
.A2(n_629),
.B1(n_630),
.B2(n_628),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1132),
.A2(n_630),
.B1(n_628),
.B2(n_642),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1128),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1149),
.B(n_1024),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1152),
.A2(n_939),
.B1(n_1085),
.B2(n_964),
.Y(n_1182)
);

OAI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_1135),
.A2(n_972),
.B1(n_454),
.B2(n_953),
.C(n_642),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1109),
.A2(n_642),
.B1(n_602),
.B2(n_606),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1155),
.B(n_1024),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1147),
.A2(n_622),
.B1(n_620),
.B2(n_618),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1124),
.A2(n_606),
.B1(n_618),
.B2(n_622),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1134),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1117),
.B(n_1030),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1115),
.B(n_1030),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1156),
.A2(n_633),
.B1(n_1018),
.B2(n_1030),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1156),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1112),
.A2(n_633),
.B1(n_855),
.B2(n_589),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1115),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1130),
.B(n_58),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1153),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1144),
.A2(n_1052),
.B1(n_1044),
.B2(n_603),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1143),
.B(n_1044),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1144),
.A2(n_1052),
.B1(n_603),
.B2(n_591),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1116),
.A2(n_1052),
.B1(n_855),
.B2(n_657),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1138),
.A2(n_591),
.B1(n_581),
.B2(n_640),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1141),
.A2(n_591),
.B1(n_581),
.B2(n_640),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1154),
.B(n_60),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1131),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1151),
.B(n_61),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1170),
.B(n_1140),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1163),
.Y(n_1207)
);

OAI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1170),
.A2(n_1129),
.B(n_1107),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1160),
.B(n_62),
.Y(n_1209)
);

AOI221xp5_ASAP7_75t_L g1210 ( 
.A1(n_1165),
.A2(n_1205),
.B1(n_1196),
.B2(n_1180),
.C(n_1172),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1188),
.B(n_62),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1188),
.B(n_63),
.Y(n_1212)
);

AND2x2_ASAP7_75t_SL g1213 ( 
.A(n_1192),
.B(n_1131),
.Y(n_1213)
);

OAI221xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1183),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.C(n_69),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1203),
.B(n_70),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1159),
.A2(n_1157),
.B(n_1146),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1166),
.B(n_1195),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1164),
.B(n_72),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1194),
.B(n_73),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1194),
.B(n_74),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1189),
.B(n_77),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1162),
.B(n_78),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1171),
.B(n_78),
.Y(n_1223)
);

OAI221xp5_ASAP7_75t_SL g1224 ( 
.A1(n_1171),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.C(n_86),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1177),
.B(n_517),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1181),
.B(n_524),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1184),
.A2(n_657),
.B1(n_650),
.B2(n_649),
.Y(n_1227)
);

OA211x2_ASAP7_75t_L g1228 ( 
.A1(n_1198),
.A2(n_88),
.B(n_90),
.C(n_91),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1185),
.B(n_95),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1173),
.A2(n_657),
.B1(n_650),
.B2(n_649),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1158),
.A2(n_98),
.B(n_99),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1177),
.B(n_100),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1174),
.B(n_1198),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1161),
.B(n_640),
.C(n_589),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1190),
.B(n_106),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1169),
.A2(n_650),
.B1(n_649),
.B2(n_645),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1191),
.B(n_108),
.Y(n_1237)
);

OAI221xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1179),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.C(n_114),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1182),
.B(n_589),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1204),
.B(n_640),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1178),
.A2(n_645),
.B1(n_520),
.B2(n_514),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1175),
.A2(n_645),
.B1(n_520),
.B2(n_514),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1207),
.B(n_1200),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1233),
.A2(n_1167),
.B1(n_1176),
.B2(n_1168),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1210),
.A2(n_1187),
.B(n_1197),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1211),
.B(n_1199),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1212),
.B(n_1201),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1212),
.B(n_1193),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1217),
.B(n_1202),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1206),
.B(n_1186),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_L g1251 ( 
.A(n_1214),
.B(n_116),
.C(n_118),
.Y(n_1251)
);

NAND4xp75_ASAP7_75t_L g1252 ( 
.A(n_1213),
.B(n_119),
.C(n_122),
.D(n_123),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1213),
.B(n_1208),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1223),
.B(n_126),
.Y(n_1254)
);

NAND2xp33_ASAP7_75t_R g1255 ( 
.A(n_1223),
.B(n_1233),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1209),
.B(n_128),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1209),
.B(n_129),
.Y(n_1257)
);

XNOR2xp5_ASAP7_75t_L g1258 ( 
.A(n_1215),
.B(n_1222),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1226),
.B(n_133),
.Y(n_1259)
);

AO21x2_ASAP7_75t_L g1260 ( 
.A1(n_1240),
.A2(n_134),
.B(n_141),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1221),
.B(n_142),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1218),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1219),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1220),
.B(n_146),
.Y(n_1264)
);

NAND4xp25_ASAP7_75t_L g1265 ( 
.A(n_1231),
.B(n_149),
.C(n_153),
.D(n_154),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1216),
.A2(n_155),
.B1(n_156),
.B2(n_160),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_L g1267 ( 
.A(n_1224),
.B(n_161),
.C(n_162),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1225),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1229),
.B(n_163),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1263),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1263),
.B(n_1229),
.Y(n_1271)
);

AND2x4_ASAP7_75t_SL g1272 ( 
.A(n_1253),
.B(n_1232),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1262),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1268),
.B(n_1246),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1243),
.Y(n_1275)
);

XNOR2xp5_ASAP7_75t_L g1276 ( 
.A(n_1258),
.B(n_1228),
.Y(n_1276)
);

XOR2x2_ASAP7_75t_L g1277 ( 
.A(n_1251),
.B(n_1238),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1246),
.B(n_1235),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1250),
.B(n_1239),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1248),
.Y(n_1280)
);

NAND4xp75_ASAP7_75t_SL g1281 ( 
.A(n_1254),
.B(n_1237),
.C(n_1242),
.D(n_1230),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1249),
.B(n_1254),
.Y(n_1282)
);

XNOR2xp5_ASAP7_75t_L g1283 ( 
.A(n_1266),
.B(n_1236),
.Y(n_1283)
);

XNOR2xp5_ASAP7_75t_L g1284 ( 
.A(n_1269),
.B(n_1227),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1247),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1255),
.B(n_1234),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1256),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1276),
.B(n_1261),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1280),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1275),
.B(n_1257),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1273),
.Y(n_1291)
);

XOR2x2_ASAP7_75t_L g1292 ( 
.A(n_1277),
.B(n_1251),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1270),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1282),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1272),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1271),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1272),
.B(n_1259),
.Y(n_1297)
);

XOR2x2_ASAP7_75t_L g1298 ( 
.A(n_1283),
.B(n_1267),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1297),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1289),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1294),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1295),
.A2(n_1282),
.B1(n_1278),
.B2(n_1286),
.Y(n_1302)
);

INVx6_ASAP7_75t_L g1303 ( 
.A(n_1297),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1288),
.A2(n_1286),
.B1(n_1279),
.B2(n_1284),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1296),
.Y(n_1305)
);

XOR2x2_ASAP7_75t_L g1306 ( 
.A(n_1292),
.B(n_1284),
.Y(n_1306)
);

AOI22x1_ASAP7_75t_L g1307 ( 
.A1(n_1298),
.A2(n_1245),
.B1(n_1281),
.B2(n_1279),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1288),
.A2(n_1287),
.B1(n_1271),
.B2(n_1285),
.Y(n_1308)
);

AOI22x1_ASAP7_75t_L g1309 ( 
.A1(n_1291),
.A2(n_1265),
.B1(n_1264),
.B2(n_1274),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1290),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1306),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1300),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1301),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1307),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1299),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1305),
.Y(n_1316)
);

OA22x2_ASAP7_75t_L g1317 ( 
.A1(n_1314),
.A2(n_1304),
.B1(n_1310),
.B2(n_1302),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1312),
.Y(n_1318)
);

OAI322xp33_ASAP7_75t_L g1319 ( 
.A1(n_1313),
.A2(n_1309),
.A3(n_1308),
.B1(n_1293),
.B2(n_1303),
.C1(n_1252),
.C2(n_1244),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1315),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1316),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1311),
.A2(n_1260),
.B1(n_1241),
.B2(n_179),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1318),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1317),
.A2(n_1241),
.B1(n_176),
.B2(n_183),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1322),
.A2(n_165),
.B1(n_184),
.B2(n_185),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1321),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1320),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1319),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_1328)
);

NOR4xp25_ASAP7_75t_L g1329 ( 
.A(n_1327),
.B(n_1319),
.C(n_201),
.D(n_203),
.Y(n_1329)
);

AO22x2_ASAP7_75t_L g1330 ( 
.A1(n_1328),
.A2(n_200),
.B1(n_204),
.B2(n_205),
.Y(n_1330)
);

AOI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1324),
.A2(n_214),
.B1(n_218),
.B2(n_221),
.C(n_228),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1323),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1329),
.A2(n_1325),
.B1(n_1326),
.B2(n_233),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1332),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1333),
.A2(n_1330),
.B1(n_1331),
.B2(n_235),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1334),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1336),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1335),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1337),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1338),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1338),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1340),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1341),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1339),
.Y(n_1344)
);

AOI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1342),
.A2(n_260),
.B1(n_263),
.B2(n_267),
.C(n_269),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1343),
.A2(n_271),
.B1(n_273),
.B2(n_276),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1346),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1345),
.Y(n_1348)
);

AO22x1_ASAP7_75t_L g1349 ( 
.A1(n_1348),
.A2(n_1344),
.B1(n_280),
.B2(n_282),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1347),
.A2(n_277),
.B1(n_284),
.B2(n_289),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1349),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1350),
.Y(n_1352)
);

AOI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1351),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.C(n_297),
.Y(n_1353)
);

AOI211xp5_ASAP7_75t_L g1354 ( 
.A1(n_1353),
.A2(n_1352),
.B(n_301),
.C(n_305),
.Y(n_1354)
);


endmodule