module fake_jpeg_30925_n_422 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_422);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_422;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_5),
.B(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_46),
.Y(n_95)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_62),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_51),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_12),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_65),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_24),
.B1(n_42),
.B2(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx12f_ASAP7_75t_SL g59 ( 
.A(n_32),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_67),
.Y(n_119)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_11),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_11),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_88),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_24),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_89),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_0),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_97),
.B1(n_56),
.B2(n_80),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_24),
.B1(n_84),
.B2(n_71),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_100),
.A2(n_109),
.B(n_115),
.C(n_133),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_40),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_70),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_129),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_46),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_23),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_23),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_51),
.B(n_42),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_30),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_54),
.A2(n_40),
.B1(n_20),
.B2(n_43),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_16),
.C(n_17),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_28),
.C(n_17),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_26),
.B1(n_39),
.B2(n_30),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_36),
.B1(n_21),
.B2(n_43),
.Y(n_184)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_40),
.B1(n_20),
.B2(n_16),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_184),
.B1(n_21),
.B2(n_68),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_147),
.B(n_149),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_47),
.B1(n_77),
.B2(n_64),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_151),
.Y(n_186)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_31),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_159),
.Y(n_220)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_111),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_110),
.Y(n_164)
);

OR2x2_ASAP7_75t_SL g165 ( 
.A(n_119),
.B(n_46),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_38),
.C(n_113),
.Y(n_205)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_93),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_170),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_31),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_173),
.Y(n_195)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_26),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_119),
.B(n_28),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_175),
.Y(n_217)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_53),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_178),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_95),
.B(n_53),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_98),
.B(n_38),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_180),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_36),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_112),
.B(n_38),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_94),
.Y(n_218)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_100),
.A2(n_36),
.B1(n_43),
.B2(n_31),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_191),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_133),
.B(n_96),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_188),
.A2(n_159),
.B(n_164),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_21),
.B(n_102),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_205),
.B(n_159),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_109),
.B(n_115),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_113),
.B(n_82),
.C(n_37),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_192),
.A2(n_120),
.B1(n_170),
.B2(n_166),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_134),
.B1(n_105),
.B2(n_74),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_117),
.C(n_137),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_162),
.A2(n_131),
.B1(n_121),
.B2(n_103),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_117),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_105),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_145),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_180),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_227),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_153),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_222),
.C(n_209),
.Y(n_271)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_146),
.B1(n_148),
.B2(n_174),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_229),
.A2(n_232),
.B1(n_249),
.B2(n_152),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_212),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_230),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_231),
.A2(n_209),
.B(n_193),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_186),
.A2(n_94),
.B1(n_120),
.B2(n_118),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_158),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_234),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_160),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_142),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_243),
.Y(n_281)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_207),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_239),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_242),
.A2(n_219),
.B1(n_182),
.B2(n_198),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_157),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_254),
.B1(n_251),
.B2(n_231),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_143),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_250),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_154),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_247),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_150),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_248),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_195),
.B(n_161),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_183),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_256),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_206),
.A2(n_163),
.B(n_141),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_255),
.B(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_192),
.A2(n_48),
.B1(n_75),
.B2(n_63),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_196),
.B1(n_206),
.B2(n_192),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_199),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_134),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_213),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_205),
.B1(n_200),
.B2(n_204),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_259),
.A2(n_263),
.B1(n_266),
.B2(n_275),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_228),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_257),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_188),
.B1(n_191),
.B2(n_210),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_229),
.A2(n_188),
.B1(n_220),
.B2(n_208),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_264),
.A2(n_265),
.B(n_269),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_220),
.B(n_193),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_283),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_256),
.B1(n_246),
.B2(n_250),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_50),
.B1(n_203),
.B2(n_194),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_243),
.A2(n_221),
.B(n_203),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_285),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_219),
.B(n_221),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_198),
.B(n_176),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_232),
.Y(n_300)
);

NAND2x1_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_155),
.Y(n_287)
);

XOR2x1_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_225),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_288),
.Y(n_317)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_289),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_224),
.Y(n_290)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_290),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_291),
.A2(n_261),
.B(n_273),
.Y(n_338)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_252),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_286),
.B1(n_275),
.B2(n_259),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_245),
.C(n_234),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_236),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_298),
.B(n_301),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_233),
.C(n_227),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_305),
.C(n_307),
.Y(n_335)
);

OA22x2_ASAP7_75t_L g328 ( 
.A1(n_300),
.A2(n_274),
.B1(n_287),
.B2(n_266),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_268),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_302),
.B(n_309),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_230),
.C(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_276),
.Y(n_306)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_247),
.C(n_240),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_310),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_280),
.B(n_248),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_277),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_238),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_262),
.B1(n_282),
.B2(n_264),
.Y(n_315)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_314),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_315),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_284),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_336),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_270),
.B1(n_273),
.B2(n_237),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_318),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_320),
.B(n_338),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_288),
.B(n_258),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_323),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_324),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_334),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_333),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_295),
.A2(n_304),
.B1(n_266),
.B2(n_300),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_292),
.A2(n_266),
.B1(n_269),
.B2(n_265),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_261),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_285),
.B(n_287),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_337),
.A2(n_292),
.B(n_312),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_326),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_319),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_345),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_344),
.A2(n_354),
.B(n_357),
.Y(n_370)
);

NOR3xp33_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_305),
.C(n_291),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_355),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_337),
.B1(n_312),
.B2(n_325),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_349),
.A2(n_356),
.B1(n_333),
.B2(n_328),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_303),
.C(n_296),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_353),
.B(n_330),
.C(n_335),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_307),
.B(n_289),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_321),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_317),
.A2(n_297),
.B1(n_308),
.B2(n_299),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_237),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_239),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_358),
.B(n_322),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_359),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_360),
.A2(n_368),
.B1(n_372),
.B2(n_374),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_364),
.C(n_369),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_335),
.C(n_336),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_316),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_371),
.Y(n_380)
);

BUFx12_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_348),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_350),
.A2(n_319),
.B1(n_328),
.B2(n_338),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_324),
.C(n_332),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_326),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_349),
.A2(n_332),
.B1(n_327),
.B2(n_322),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_272),
.C(n_235),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_373),
.B(n_339),
.C(n_357),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_226),
.B1(n_1),
.B2(n_3),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_363),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_383),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_366),
.A2(n_344),
.B(n_357),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_377),
.B(n_381),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_367),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_361),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_373),
.C(n_369),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_386),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_380),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_346),
.C(n_351),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_372),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_368),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_370),
.B(n_351),
.Y(n_389)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_389),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_392),
.B(n_396),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_394),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_360),
.B1(n_340),
.B2(n_342),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_398),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_367),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_382),
.A2(n_346),
.B(n_342),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_397),
.A2(n_0),
.B(n_3),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_365),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_390),
.A2(n_376),
.B(n_385),
.Y(n_399)
);

AOI21x1_ASAP7_75t_L g409 ( 
.A1(n_399),
.A2(n_400),
.B(n_394),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_386),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_406),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_0),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_401),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_391),
.C(n_397),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_404),
.B(n_388),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_409),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_412),
.C(n_413),
.Y(n_414)
);

AOI21xp33_ASAP7_75t_L g412 ( 
.A1(n_402),
.A2(n_407),
.B(n_406),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_403),
.B(n_0),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_38),
.C(n_5),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_415),
.Y(n_417)
);

OAI21x1_ASAP7_75t_SL g418 ( 
.A1(n_414),
.A2(n_4),
.B(n_5),
.Y(n_418)
);

O2A1O1Ixp33_ASAP7_75t_SL g419 ( 
.A1(n_418),
.A2(n_416),
.B(n_5),
.C(n_6),
.Y(n_419)
);

OAI321xp33_ASAP7_75t_L g420 ( 
.A1(n_419),
.A2(n_417),
.A3(n_8),
.B1(n_10),
.B2(n_4),
.C(n_38),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_10),
.C(n_4),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_8),
.Y(n_422)
);


endmodule