module real_aes_11835_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_1369;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g1102 ( .A(n_0), .Y(n_1102) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_1), .A2(n_447), .B1(n_450), .B2(n_459), .C(n_462), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g517 ( .A1(n_1), .A2(n_518), .B(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g702 ( .A(n_2), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_2), .A2(n_72), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_3), .A2(n_232), .B1(n_285), .B2(n_512), .Y(n_710) );
INVx1_ASAP7_75t_L g742 ( .A(n_3), .Y(n_742) );
INVx1_ASAP7_75t_L g759 ( .A(n_4), .Y(n_759) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_4), .A2(n_31), .B1(n_792), .B2(n_793), .C(n_794), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_5), .A2(n_74), .B1(n_629), .B2(n_630), .Y(n_637) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_5), .Y(n_666) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_6), .Y(n_247) );
AND2x2_ASAP7_75t_L g337 ( .A(n_6), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g392 ( .A(n_6), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_6), .B(n_181), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_7), .A2(n_139), .B1(n_273), .B2(n_593), .C(n_708), .Y(n_1313) );
INVx1_ASAP7_75t_L g1346 ( .A(n_7), .Y(n_1346) );
INVx1_ASAP7_75t_L g374 ( .A(n_8), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g884 ( .A1(n_9), .A2(n_413), .B1(n_885), .B2(n_891), .C(n_897), .Y(n_884) );
INVx1_ASAP7_75t_L g913 ( .A(n_9), .Y(n_913) );
INVx1_ASAP7_75t_L g383 ( .A(n_10), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_11), .A2(n_23), .B1(n_468), .B2(n_471), .C(n_472), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_11), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_12), .A2(n_57), .B1(n_388), .B2(n_473), .C(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g918 ( .A(n_12), .Y(n_918) );
INVx1_ASAP7_75t_L g873 ( .A(n_13), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_13), .A2(n_58), .B1(n_649), .B2(n_659), .Y(n_915) );
AO22x2_ASAP7_75t_L g922 ( .A1(n_14), .A2(n_923), .B1(n_977), .B2(n_978), .Y(n_922) );
CKINVDCx14_ASAP7_75t_R g977 ( .A(n_14), .Y(n_977) );
INVx1_ASAP7_75t_L g1195 ( .A(n_15), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_16), .A2(n_80), .B1(n_699), .B2(n_991), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_16), .A2(n_32), .B1(n_336), .B2(n_397), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_17), .A2(n_207), .B1(n_763), .B2(n_764), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_17), .A2(n_66), .B1(n_505), .B2(n_584), .C(n_802), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_18), .A2(n_40), .B1(n_505), .B2(n_707), .C(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g744 ( .A(n_18), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_19), .A2(n_66), .B1(n_766), .B2(n_768), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_19), .A2(n_207), .B1(n_804), .B2(n_805), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_20), .A2(n_225), .B1(n_802), .B2(n_821), .C(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g844 ( .A(n_20), .Y(n_844) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_21), .A2(n_201), .B1(n_802), .B2(n_961), .C(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1059 ( .A(n_21), .Y(n_1059) );
AO221x2_ASAP7_75t_L g1123 ( .A1(n_22), .A2(n_59), .B1(n_1100), .B2(n_1114), .C(n_1124), .Y(n_1123) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_23), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_24), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g1013 ( .A1(n_25), .A2(n_132), .B1(n_388), .B2(n_1014), .C(n_1015), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_25), .A2(n_200), .B1(n_437), .B2(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g268 ( .A(n_26), .Y(n_268) );
OR2x2_ASAP7_75t_L g427 ( .A(n_26), .B(n_316), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g562 ( .A1(n_27), .A2(n_169), .B1(n_563), .B2(n_564), .C(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g576 ( .A(n_27), .Y(n_576) );
AO22x1_ASAP7_75t_L g868 ( .A1(n_28), .A2(n_869), .B1(n_920), .B2(n_921), .Y(n_868) );
INVx1_ASAP7_75t_L g921 ( .A(n_28), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_29), .A2(n_64), .B1(n_950), .B2(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1010 ( .A(n_29), .Y(n_1010) );
INVx1_ASAP7_75t_L g1142 ( .A(n_30), .Y(n_1142) );
INVx1_ASAP7_75t_L g758 ( .A(n_31), .Y(n_758) );
OAI222xp33_ASAP7_75t_L g1020 ( .A1(n_32), .A2(n_132), .B1(n_138), .B2(n_643), .C1(n_1021), .C2(n_1023), .Y(n_1020) );
BUFx2_ASAP7_75t_L g270 ( .A(n_33), .Y(n_270) );
BUFx2_ASAP7_75t_L g304 ( .A(n_33), .Y(n_304) );
INVx1_ASAP7_75t_L g318 ( .A(n_33), .Y(n_318) );
OR2x2_ASAP7_75t_L g470 ( .A(n_33), .B(n_399), .Y(n_470) );
INVx1_ASAP7_75t_L g1194 ( .A(n_34), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_34), .A2(n_1361), .B1(n_1365), .B2(n_1368), .Y(n_1360) );
INVx1_ASAP7_75t_L g926 ( .A(n_35), .Y(n_926) );
AOI21xp33_ASAP7_75t_L g966 ( .A1(n_35), .A2(n_649), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g542 ( .A(n_36), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_37), .A2(n_144), .B1(n_400), .B2(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g508 ( .A(n_37), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g938 ( .A(n_38), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g1317 ( .A(n_39), .Y(n_1317) );
INVx1_ASAP7_75t_L g737 ( .A(n_40), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_41), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_42), .A2(n_67), .B1(n_827), .B2(n_1039), .Y(n_1038) );
OAI221xp5_ASAP7_75t_L g1061 ( .A1(n_42), .A2(n_67), .B1(n_472), .B2(n_730), .C(n_731), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_43), .A2(n_165), .B1(n_629), .B2(n_630), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_43), .A2(n_219), .B1(n_297), .B2(n_668), .C(n_671), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_44), .A2(n_83), .B1(n_418), .B2(n_464), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_44), .A2(n_83), .B1(n_489), .B2(n_493), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g968 ( .A1(n_45), .A2(n_199), .B1(n_969), .B2(n_970), .C(n_972), .Y(n_968) );
INVx1_ASAP7_75t_L g975 ( .A(n_45), .Y(n_975) );
CKINVDCx16_ASAP7_75t_R g1139 ( .A(n_46), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_47), .A2(n_56), .B1(n_774), .B2(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g809 ( .A(n_47), .Y(n_809) );
INVx1_ASAP7_75t_L g890 ( .A(n_48), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_48), .A2(n_127), .B1(n_273), .B2(n_659), .Y(n_911) );
INVx1_ASAP7_75t_L g1190 ( .A(n_49), .Y(n_1190) );
INVx1_ASAP7_75t_L g552 ( .A(n_50), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_51), .A2(n_140), .B1(n_881), .B2(n_883), .Y(n_880) );
OAI22xp5_ASAP7_75t_SL g904 ( .A1(n_51), .A2(n_140), .B1(n_309), .B2(n_321), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_52), .Y(n_319) );
INVx1_ASAP7_75t_L g998 ( .A(n_53), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_53), .A2(n_81), .B1(n_881), .B2(n_883), .C(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g453 ( .A(n_54), .Y(n_453) );
AOI21xp33_ASAP7_75t_L g504 ( .A1(n_54), .A2(n_505), .B(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_55), .A2(n_87), .B1(n_633), .B2(n_634), .Y(n_636) );
INVxp33_ASAP7_75t_SL g680 ( .A(n_55), .Y(n_680) );
INVx1_ASAP7_75t_L g800 ( .A(n_56), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_57), .A2(n_99), .B1(n_429), .B2(n_437), .Y(n_919) );
INVx1_ASAP7_75t_L g874 ( .A(n_58), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g1324 ( .A(n_60), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_61), .A2(n_179), .B1(n_297), .B2(n_298), .Y(n_296) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_61), .A2(n_231), .B1(n_333), .B2(n_343), .Y(n_332) );
INVx1_ASAP7_75t_L g1153 ( .A(n_62), .Y(n_1153) );
CKINVDCx16_ASAP7_75t_R g1158 ( .A(n_63), .Y(n_1158) );
INVx1_ASAP7_75t_L g1008 ( .A(n_64), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_65), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_68), .A2(n_226), .B1(n_512), .B2(n_804), .Y(n_1048) );
INVx1_ASAP7_75t_L g1064 ( .A(n_68), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_69), .A2(n_114), .B1(n_376), .B2(n_548), .C(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_69), .A2(n_84), .B1(n_587), .B2(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g1103 ( .A(n_70), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_71), .A2(n_212), .B1(n_491), .B2(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g845 ( .A(n_71), .Y(n_845) );
INVx1_ASAP7_75t_L g703 ( .A(n_72), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_73), .Y(n_456) );
INVxp33_ASAP7_75t_L g678 ( .A(n_74), .Y(n_678) );
INVx1_ASAP7_75t_L g551 ( .A(n_75), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_75), .A2(n_114), .B1(n_581), .B2(n_582), .C(n_584), .Y(n_580) );
CKINVDCx16_ASAP7_75t_R g1160 ( .A(n_76), .Y(n_1160) );
AOI22xp5_ASAP7_75t_L g1120 ( .A1(n_77), .A2(n_121), .B1(n_1108), .B2(n_1111), .Y(n_1120) );
INVx1_ASAP7_75t_L g267 ( .A(n_78), .Y(n_267) );
INVx1_ASAP7_75t_L g316 ( .A(n_78), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_79), .A2(n_224), .B1(n_595), .B2(n_991), .Y(n_1314) );
INVx1_ASAP7_75t_L g1351 ( .A(n_79), .Y(n_1351) );
INVx1_ASAP7_75t_L g1016 ( .A(n_80), .Y(n_1016) );
INVx1_ASAP7_75t_L g997 ( .A(n_81), .Y(n_997) );
INVx1_ASAP7_75t_L g567 ( .A(n_82), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_82), .A2(n_169), .B1(n_572), .B2(n_574), .C(n_575), .Y(n_571) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_84), .Y(n_550) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_85), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_85), .A2(n_191), .B1(n_651), .B2(n_653), .Y(n_650) );
NAND2xp33_ASAP7_75t_SL g698 ( .A(n_86), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g725 ( .A(n_86), .Y(n_725) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_87), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_88), .A2(n_133), .B1(n_483), .B2(n_486), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_88), .A2(n_187), .B1(n_274), .B2(n_512), .Y(n_516) );
INVx1_ASAP7_75t_L g559 ( .A(n_89), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_89), .A2(n_125), .B1(n_520), .B2(n_592), .C(n_593), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_90), .A2(n_187), .B1(n_476), .B2(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g514 ( .A(n_90), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_91), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_92), .Y(n_691) );
OAI21xp33_ASAP7_75t_L g533 ( .A1(n_93), .A2(n_534), .B(n_569), .Y(n_533) );
INVx1_ASAP7_75t_L g603 ( .A(n_93), .Y(n_603) );
INVx1_ASAP7_75t_L g1141 ( .A(n_93), .Y(n_1141) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_94), .A2(n_147), .B1(n_670), .B2(n_821), .Y(n_989) );
AOI21xp33_ASAP7_75t_L g1006 ( .A1(n_94), .A2(n_400), .B(n_460), .Y(n_1006) );
INVx1_ASAP7_75t_L g568 ( .A(n_95), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g829 ( .A1(n_96), .A2(n_198), .B1(n_506), .B2(n_802), .C(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g852 ( .A(n_96), .Y(n_852) );
AO221x2_ASAP7_75t_L g1095 ( .A1(n_97), .A2(n_161), .B1(n_1096), .B2(n_1100), .C(n_1101), .Y(n_1095) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_98), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_99), .A2(n_109), .B1(n_563), .B2(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g239 ( .A(n_100), .Y(n_239) );
INVx1_ASAP7_75t_L g718 ( .A(n_101), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_102), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_103), .Y(n_935) );
OA22x2_ASAP7_75t_L g815 ( .A1(n_104), .A2(n_816), .B1(n_863), .B2(n_864), .Y(n_815) );
INVx1_ASAP7_75t_L g864 ( .A(n_104), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_105), .A2(n_172), .B1(n_770), .B2(n_772), .Y(n_769) );
INVx1_ASAP7_75t_L g810 ( .A(n_105), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_106), .Y(n_1051) );
INVx1_ASAP7_75t_L g1076 ( .A(n_107), .Y(n_1076) );
OAI221xp5_ASAP7_75t_SL g555 ( .A1(n_108), .A2(n_211), .B1(n_556), .B2(n_557), .C(n_558), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_108), .A2(n_211), .B1(n_273), .B2(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g917 ( .A(n_109), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_110), .A2(n_174), .B1(n_805), .B2(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1056 ( .A(n_110), .Y(n_1056) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_111), .A2(n_156), .B1(n_1100), .B2(n_1114), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_112), .A2(n_192), .B1(n_278), .B2(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g728 ( .A(n_112), .Y(n_728) );
XOR2xp5_ASAP7_75t_L g443 ( .A(n_113), .B(n_444), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g1329 ( .A(n_115), .Y(n_1329) );
INVx1_ASAP7_75t_L g1125 ( .A(n_116), .Y(n_1125) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_117), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_118), .Y(n_940) );
INVx1_ASAP7_75t_L g813 ( .A(n_119), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_120), .Y(n_836) );
XNOR2xp5_ASAP7_75t_L g982 ( .A(n_121), .B(n_983), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_122), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_123), .A2(n_233), .B1(n_593), .B2(n_961), .C(n_1035), .Y(n_1327) );
INVx1_ASAP7_75t_L g1334 ( .A(n_123), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_124), .A2(n_221), .B1(n_272), .B2(n_277), .Y(n_271) );
INVx1_ASAP7_75t_L g356 ( .A(n_124), .Y(n_356) );
INVx1_ASAP7_75t_L g561 ( .A(n_125), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g1050 ( .A(n_126), .Y(n_1050) );
INVx1_ASAP7_75t_L g888 ( .A(n_127), .Y(n_888) );
INVx1_ASAP7_75t_L g1319 ( .A(n_128), .Y(n_1319) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_128), .A2(n_209), .B1(n_471), .B2(n_1339), .C(n_1341), .Y(n_1338) );
INVx1_ASAP7_75t_L g778 ( .A(n_129), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_129), .A2(n_203), .B1(n_274), .B2(n_300), .Y(n_795) );
INVx1_ASAP7_75t_L g927 ( .A(n_130), .Y(n_927) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_130), .A2(n_177), .B1(n_659), .B2(n_965), .Y(n_964) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_131), .Y(n_1042) );
INVx1_ASAP7_75t_L g522 ( .A(n_133), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g1312 ( .A(n_134), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_135), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g1129 ( .A1(n_136), .A2(n_149), .B1(n_1108), .B2(n_1111), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_137), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_138), .A2(n_200), .B1(n_548), .B2(n_877), .Y(n_1012) );
INVx1_ASAP7_75t_L g1348 ( .A(n_139), .Y(n_1348) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_141), .A2(n_153), .B1(n_278), .B2(n_697), .Y(n_993) );
INVx1_ASAP7_75t_L g1001 ( .A(n_141), .Y(n_1001) );
XOR2x2_ASAP7_75t_L g604 ( .A(n_142), .B(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_143), .A2(n_231), .B1(n_284), .B2(n_290), .Y(n_295) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_143), .A2(n_179), .B1(n_413), .B2(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g503 ( .A(n_144), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_145), .A2(n_167), .B1(n_944), .B2(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g955 ( .A(n_145), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_146), .A2(n_188), .B1(n_483), .B2(n_486), .Y(n_946) );
AOI22xp33_ASAP7_75t_SL g958 ( .A1(n_146), .A2(n_167), .B1(n_649), .B2(n_659), .Y(n_958) );
INVx1_ASAP7_75t_L g1005 ( .A(n_147), .Y(n_1005) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_148), .A2(n_205), .B1(n_1044), .B2(n_1046), .C(n_1047), .Y(n_1043) );
INVx1_ASAP7_75t_L g1071 ( .A(n_148), .Y(n_1071) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_150), .Y(n_936) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_151), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_151), .B(n_239), .Y(n_1084) );
AND3x2_ASAP7_75t_L g1099 ( .A(n_151), .B(n_239), .C(n_1087), .Y(n_1099) );
OA332x1_ASAP7_75t_L g924 ( .A1(n_152), .A2(n_447), .A3(n_459), .B1(n_925), .B2(n_930), .B3(n_933), .C1(n_937), .C2(n_941), .Y(n_924) );
AOI21xp5_ASAP7_75t_L g959 ( .A1(n_152), .A2(n_960), .B(n_961), .Y(n_959) );
INVx1_ASAP7_75t_L g1002 ( .A(n_153), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_154), .A2(n_184), .B1(n_1096), .B2(n_1131), .Y(n_1130) );
INVx2_ASAP7_75t_L g252 ( .A(n_155), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_157), .A2(n_216), .B1(n_821), .B2(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g849 ( .A(n_157), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_158), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_159), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g871 ( .A1(n_160), .A2(n_343), .B(n_872), .C(n_875), .Y(n_871) );
INVx1_ASAP7_75t_L g914 ( .A(n_160), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_162), .A2(n_168), .B1(n_1100), .B2(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g538 ( .A(n_163), .Y(n_538) );
INVxp33_ASAP7_75t_SL g622 ( .A(n_164), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_164), .A2(n_206), .B1(n_656), .B2(n_658), .C(n_660), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_165), .A2(n_186), .B1(n_595), .B2(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g1087 ( .A(n_166), .Y(n_1087) );
CKINVDCx16_ASAP7_75t_R g1137 ( .A(n_170), .Y(n_1137) );
INVx1_ASAP7_75t_L g1192 ( .A(n_171), .Y(n_1192) );
INVx1_ASAP7_75t_L g790 ( .A(n_172), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_173), .A2(n_228), .B1(n_400), .B2(n_458), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_173), .A2(n_228), .B1(n_496), .B2(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g1060 ( .A(n_174), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_175), .A2(n_215), .B1(n_284), .B2(n_290), .Y(n_283) );
INVx1_ASAP7_75t_L g368 ( .A(n_175), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_176), .Y(n_811) );
INVx1_ASAP7_75t_L g931 ( .A(n_177), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_178), .Y(n_1033) );
XNOR2xp5_ASAP7_75t_L g1366 ( .A(n_180), .B(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g254 ( .A(n_181), .Y(n_254) );
INVx2_ASAP7_75t_L g338 ( .A(n_181), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_182), .A2(n_213), .B1(n_1108), .B2(n_1111), .Y(n_1107) );
INVx1_ASAP7_75t_L g900 ( .A(n_183), .Y(n_900) );
INVx1_ASAP7_75t_L g782 ( .A(n_185), .Y(n_782) );
AOI21xp33_ASAP7_75t_L g796 ( .A1(n_185), .A2(n_520), .B(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_186), .A2(n_219), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g973 ( .A(n_188), .Y(n_973) );
CKINVDCx5p33_ASAP7_75t_R g1316 ( .A(n_189), .Y(n_1316) );
INVx1_ASAP7_75t_L g403 ( .A(n_190), .Y(n_403) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_191), .Y(n_612) );
INVx1_ASAP7_75t_L g723 ( .A(n_192), .Y(n_723) );
XOR2xp5_ASAP7_75t_L g259 ( .A(n_193), .B(n_260), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_194), .Y(n_713) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_195), .Y(n_825) );
INVx1_ASAP7_75t_L g617 ( .A(n_196), .Y(n_617) );
INVx1_ASAP7_75t_L g379 ( .A(n_197), .Y(n_379) );
INVx1_ASAP7_75t_L g850 ( .A(n_198), .Y(n_850) );
INVx1_ASAP7_75t_L g976 ( .A(n_199), .Y(n_976) );
INVx1_ASAP7_75t_L g1057 ( .A(n_201), .Y(n_1057) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_202), .A2(n_210), .B1(n_793), .B2(n_827), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g846 ( .A1(n_202), .A2(n_210), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_846) );
INVx1_ASAP7_75t_L g783 ( .A(n_203), .Y(n_783) );
INVx1_ASAP7_75t_L g1154 ( .A(n_204), .Y(n_1154) );
INVx1_ASAP7_75t_L g1067 ( .A(n_205), .Y(n_1067) );
INVxp33_ASAP7_75t_SL g614 ( .A(n_206), .Y(n_614) );
INVx1_ASAP7_75t_L g1088 ( .A(n_208), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_208), .B(n_1086), .Y(n_1105) );
INVx1_ASAP7_75t_L g1320 ( .A(n_209), .Y(n_1320) );
INVx1_ASAP7_75t_L g841 ( .A(n_212), .Y(n_841) );
INVx1_ASAP7_75t_L g1330 ( .A(n_214), .Y(n_1330) );
INVx1_ASAP7_75t_L g364 ( .A(n_215), .Y(n_364) );
INVx1_ASAP7_75t_L g854 ( .A(n_216), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_217), .Y(n_895) );
INVx2_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g1326 ( .A(n_220), .Y(n_1326) );
INVx1_ASAP7_75t_L g350 ( .A(n_221), .Y(n_350) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_222), .A2(n_285), .B(n_520), .Y(n_701) );
INVx1_ASAP7_75t_L g727 ( .A(n_222), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g932 ( .A(n_223), .Y(n_932) );
INVx1_ASAP7_75t_L g1344 ( .A(n_224), .Y(n_1344) );
INVx1_ASAP7_75t_L g842 ( .A(n_225), .Y(n_842) );
INVx1_ASAP7_75t_L g1072 ( .A(n_226), .Y(n_1072) );
INVx1_ASAP7_75t_L g1052 ( .A(n_227), .Y(n_1052) );
BUFx3_ASAP7_75t_L g276 ( .A(n_229), .Y(n_276) );
INVx1_ASAP7_75t_L g282 ( .A(n_229), .Y(n_282) );
INVx1_ASAP7_75t_L g275 ( .A(n_230), .Y(n_275) );
BUFx3_ASAP7_75t_L g281 ( .A(n_230), .Y(n_281) );
INVx1_ASAP7_75t_L g739 ( .A(n_232), .Y(n_739) );
INVx1_ASAP7_75t_L g1336 ( .A(n_233), .Y(n_1336) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_255), .B(n_1080), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_242), .Y(n_236) );
AND2x4_ASAP7_75t_L g1359 ( .A(n_237), .B(n_243), .Y(n_1359) );
NOR2xp33_ASAP7_75t_SL g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx1_ASAP7_75t_SL g1364 ( .A(n_238), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_238), .B(n_240), .Y(n_1369) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_240), .B(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g371 ( .A(n_246), .B(n_254), .Y(n_371) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g460 ( .A(n_247), .B(n_461), .Y(n_460) );
OR2x6_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
BUFx2_ASAP7_75t_L g367 ( .A(n_249), .Y(n_367) );
INVx1_ASAP7_75t_L g385 ( .A(n_249), .Y(n_385) );
OR2x2_ASAP7_75t_L g486 ( .A(n_249), .B(n_470), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_249), .A2(n_381), .B1(n_550), .B2(n_551), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_249), .A2(n_381), .B1(n_567), .B2(n_568), .Y(n_566) );
INVx2_ASAP7_75t_SL g894 ( .A(n_249), .Y(n_894) );
BUFx6f_ASAP7_75t_L g934 ( .A(n_249), .Y(n_934) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x4_ASAP7_75t_L g341 ( .A(n_251), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_251), .Y(n_347) );
INVx2_ASAP7_75t_L g355 ( .A(n_251), .Y(n_355) );
INVx1_ASAP7_75t_L g363 ( .A(n_251), .Y(n_363) );
AND2x2_ASAP7_75t_L g402 ( .A(n_251), .B(n_252), .Y(n_402) );
INVx2_ASAP7_75t_L g342 ( .A(n_252), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_252), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g362 ( .A(n_252), .Y(n_362) );
INVx1_ASAP7_75t_L g409 ( .A(n_252), .Y(n_409) );
INVx1_ASAP7_75t_L g420 ( .A(n_252), .Y(n_420) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_686), .Y(n_255) );
BUFx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
AO22x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_604), .B1(n_684), .B2(n_685), .Y(n_257) );
INVx1_ASAP7_75t_L g684 ( .A(n_258), .Y(n_684) );
XNOR2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_442), .Y(n_258) );
NAND4xp75_ASAP7_75t_L g260 ( .A(n_261), .B(n_331), .C(n_423), .D(n_432), .Y(n_260) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_262), .B(n_307), .Y(n_261) );
AOI33xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_271), .A3(n_283), .B1(n_295), .B2(n_296), .B3(n_301), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_264), .Y(n_263) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
INVx1_ASAP7_75t_L g709 ( .A(n_265), .Y(n_709) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_SL g506 ( .A(n_266), .Y(n_506) );
BUFx3_ASAP7_75t_L g585 ( .A(n_266), .Y(n_585) );
INVx1_ASAP7_75t_L g907 ( .A(n_266), .Y(n_907) );
INVx1_ASAP7_75t_L g967 ( .A(n_266), .Y(n_967) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x4_ASAP7_75t_L g305 ( .A(n_267), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_268), .Y(n_306) );
AND2x2_ASAP7_75t_L g466 ( .A(n_269), .B(n_389), .Y(n_466) );
AND2x4_ASAP7_75t_L g546 ( .A(n_269), .B(n_371), .Y(n_546) );
INVx2_ASAP7_75t_L g599 ( .A(n_269), .Y(n_599) );
AND2x4_ASAP7_75t_L g627 ( .A(n_269), .B(n_371), .Y(n_627) );
BUFx2_ASAP7_75t_L g717 ( .A(n_269), .Y(n_717) );
OR2x2_ASAP7_75t_L g906 ( .A(n_269), .B(n_907), .Y(n_906) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g422 ( .A(n_270), .Y(n_422) );
OR2x6_ASAP7_75t_L g459 ( .A(n_270), .B(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx3_ASAP7_75t_L g297 ( .A(n_273), .Y(n_297) );
INVx1_ASAP7_75t_L g657 ( .A(n_273), .Y(n_657) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_SL g435 ( .A(n_274), .Y(n_435) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_274), .Y(n_491) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_274), .Y(n_505) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_274), .Y(n_649) );
BUFx3_ASAP7_75t_L g697 ( .A(n_274), .Y(n_697) );
BUFx2_ASAP7_75t_L g830 ( .A(n_274), .Y(n_830) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_274), .Y(n_1037) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g441 ( .A(n_275), .Y(n_441) );
INVx2_ASAP7_75t_L g288 ( .A(n_276), .Y(n_288) );
AND2x2_ASAP7_75t_L g294 ( .A(n_276), .B(n_281), .Y(n_294) );
BUFx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x6_ASAP7_75t_L g429 ( .A(n_279), .B(n_426), .Y(n_429) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_279), .B(n_426), .Y(n_1026) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_280), .Y(n_300) );
INVx2_ASAP7_75t_L g494 ( .A(n_280), .Y(n_494) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_280), .Y(n_659) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g289 ( .A(n_281), .Y(n_289) );
INVx1_ASAP7_75t_L g440 ( .A(n_282), .Y(n_440) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g424 ( .A(n_285), .B(n_425), .Y(n_424) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_285), .A2(n_522), .B(n_523), .C(n_529), .Y(n_521) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g674 ( .A(n_286), .Y(n_674) );
INVx1_ASAP7_75t_L g960 ( .A(n_286), .Y(n_960) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g431 ( .A(n_287), .B(n_314), .Y(n_431) );
INVx6_ASAP7_75t_L g519 ( .A(n_287), .Y(n_519) );
BUFx2_ASAP7_75t_L g804 ( .A(n_287), .Y(n_804) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
INVx1_ASAP7_75t_L g324 ( .A(n_289), .Y(n_324) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g675 ( .A(n_292), .B(n_676), .Y(n_675) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g329 ( .A(n_293), .Y(n_329) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_293), .Y(n_593) );
INVx2_ASAP7_75t_L g700 ( .A(n_293), .Y(n_700) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_294), .Y(n_500) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g574 ( .A(n_300), .Y(n_574) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_300), .Y(n_595) );
BUFx6f_ASAP7_75t_L g950 ( .A(n_300), .Y(n_950) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_SL g905 ( .A1(n_302), .A2(n_906), .B1(n_908), .B2(n_912), .Y(n_905) );
INVx4_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x4_ASAP7_75t_L g430 ( .A(n_304), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_L g994 ( .A(n_304), .B(n_305), .Y(n_994) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_305), .Y(n_520) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_305), .Y(n_663) );
INVx1_ASAP7_75t_L g822 ( .A(n_305), .Y(n_822) );
INVx2_ASAP7_75t_SL g961 ( .A(n_305), .Y(n_961) );
AND2x4_ASAP7_75t_L g314 ( .A(n_306), .B(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_319), .B1(n_320), .B2(n_326), .C(n_327), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_308), .A2(n_327), .B1(n_996), .B2(n_997), .C(n_998), .Y(n_995) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x6_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
OR2x2_ASAP7_75t_L g653 ( .A(n_310), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_311), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_525) );
AND2x4_ASAP7_75t_L g578 ( .A(n_311), .B(n_314), .Y(n_578) );
AND2x2_ASAP7_75t_L g971 ( .A(n_311), .B(n_314), .Y(n_971) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_311), .B(n_314), .Y(n_1321) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_SL g325 ( .A(n_313), .Y(n_325) );
INVx1_ASAP7_75t_L g330 ( .A(n_313), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
BUFx2_ASAP7_75t_L g530 ( .A(n_314), .Y(n_530) );
AND2x4_ASAP7_75t_L g577 ( .A(n_314), .B(n_526), .Y(n_577) );
AND2x4_ASAP7_75t_L g652 ( .A(n_314), .B(n_526), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_314), .Y(n_654) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x6_ASAP7_75t_L g639 ( .A(n_317), .B(n_390), .Y(n_639) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g426 ( .A(n_318), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g449 ( .A(n_318), .B(n_337), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_319), .A2(n_326), .B1(n_407), .B2(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g996 ( .A(n_321), .Y(n_996) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g526 ( .A(n_323), .Y(n_526) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR3xp33_ASAP7_75t_L g903 ( .A(n_327), .B(n_904), .C(n_905), .Y(n_903) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI31xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_348), .A3(n_412), .B(n_421), .Y(n_331) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_334), .A2(n_417), .B1(n_873), .B2(n_874), .Y(n_872) );
AOI221x1_ASAP7_75t_L g1000 ( .A1(n_334), .A2(n_417), .B1(n_1001), .B2(n_1002), .C(n_1003), .Y(n_1000) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
AND2x4_ASAP7_75t_L g344 ( .A(n_335), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g414 ( .A(n_337), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g417 ( .A(n_337), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g391 ( .A(n_338), .Y(n_391) );
INVx1_ASAP7_75t_L g461 ( .A(n_338), .Y(n_461) );
INVx1_ASAP7_75t_L g1009 ( .A(n_339), .Y(n_1009) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g464 ( .A(n_340), .Y(n_464) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_341), .Y(n_358) );
INVx3_ASAP7_75t_L g378 ( .A(n_341), .Y(n_378) );
AND2x4_ASAP7_75t_L g346 ( .A(n_342), .B(n_347), .Y(n_346) );
INVx8_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_SL g1011 ( .A1(n_344), .A2(n_1012), .B1(n_1013), .B2(n_1016), .C(n_1017), .Y(n_1011) );
BUFx6f_ASAP7_75t_L g1015 ( .A(n_345), .Y(n_1015) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_346), .Y(n_458) );
BUFx3_ASAP7_75t_L g473 ( .A(n_346), .Y(n_473) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_346), .Y(n_481) );
BUFx2_ASAP7_75t_L g544 ( .A(n_346), .Y(n_544) );
OAI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_359), .B1(n_372), .B2(n_380), .C(n_393), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_356), .B2(n_357), .Y(n_349) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g373 ( .A(n_352), .Y(n_373) );
BUFx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g556 ( .A(n_353), .Y(n_556) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g452 ( .A(n_354), .Y(n_452) );
BUFx2_ASAP7_75t_L g887 ( .A(n_354), .Y(n_887) );
INVx1_ASAP7_75t_L g411 ( .A(n_355), .Y(n_411) );
AND2x4_ASAP7_75t_L g418 ( .A(n_355), .B(n_419), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_357), .A2(n_938), .B1(n_939), .B2(n_940), .Y(n_937) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g635 ( .A(n_358), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .B1(n_365), .B2(n_368), .C(n_369), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g405 ( .A(n_361), .Y(n_405) );
BUFx2_ASAP7_75t_L g750 ( .A(n_361), .Y(n_750) );
INVx2_ASAP7_75t_L g862 ( .A(n_361), .Y(n_862) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_362), .B(n_363), .Y(n_382) );
INVx1_ASAP7_75t_L g541 ( .A(n_363), .Y(n_541) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g741 ( .A(n_366), .Y(n_741) );
INVx2_ASAP7_75t_SL g748 ( .A(n_366), .Y(n_748) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_SL g896 ( .A(n_371), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_375), .B2(n_379), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_374), .A2(n_383), .B1(n_433), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g877 ( .A(n_377), .Y(n_877) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g455 ( .A(n_378), .Y(n_455) );
INVx3_ASAP7_75t_L g485 ( .A(n_378), .Y(n_485) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_379), .A2(n_386), .B1(n_403), .B2(n_424), .C1(n_428), .C2(n_430), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B1(n_384), .B2(n_386), .C(n_387), .Y(n_380) );
BUFx3_ASAP7_75t_L g743 ( .A(n_381), .Y(n_743) );
OAI22xp33_ASAP7_75t_L g933 ( .A1(n_381), .A2(n_934), .B1(n_935), .B2(n_936), .Y(n_933) );
INVx2_ASAP7_75t_L g1066 ( .A(n_381), .Y(n_1066) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_403), .B(n_404), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NOR2xp67_ASAP7_75t_L g902 ( .A(n_395), .B(n_599), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_397), .A2(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g882 ( .A(n_397), .Y(n_882) );
OR2x6_ASAP7_75t_L g883 ( .A(n_397), .B(n_411), .Y(n_883) );
OR2x6_ASAP7_75t_L g897 ( .A(n_397), .B(n_862), .Y(n_897) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g448 ( .A(n_400), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g560 ( .A(n_401), .Y(n_560) );
INVx2_ASAP7_75t_L g763 ( .A(n_401), .Y(n_763) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_402), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_405), .A2(n_892), .B1(n_893), .B2(n_895), .C(n_896), .Y(n_891) );
OAI21xp5_ASAP7_75t_SL g1004 ( .A1(n_405), .A2(n_1005), .B(n_1006), .Y(n_1004) );
NAND2x1_ASAP7_75t_SL g468 ( .A(n_407), .B(n_469), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g881 ( .A(n_407), .B(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_409), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_410), .B(n_469), .Y(n_471) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
CKINVDCx6p67_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_415), .Y(n_879) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_415), .Y(n_1014) );
INVx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_418), .Y(n_478) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_418), .Y(n_548) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_418), .Y(n_563) );
INVx1_ASAP7_75t_L g767 ( .A(n_418), .Y(n_767) );
INVx1_ASAP7_75t_L g771 ( .A(n_418), .Y(n_771) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g531 ( .A(n_421), .Y(n_531) );
BUFx8_ASAP7_75t_SL g898 ( .A(n_421), .Y(n_898) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g683 ( .A(n_422), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g916 ( .A1(n_424), .A2(n_433), .B1(n_917), .B2(n_918), .C(n_919), .Y(n_916) );
AND2x2_ASAP7_75t_L g433 ( .A(n_425), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x6_ASAP7_75t_L g437 ( .A(n_426), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_426), .B(n_1022), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_426), .B(n_1024), .Y(n_1023) );
INVx2_ASAP7_75t_L g492 ( .A(n_427), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_427), .B(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g496 ( .A(n_427), .B(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g948 ( .A1(n_427), .A2(n_949), .B(n_951), .C(n_952), .Y(n_948) );
CKINVDCx6p67_ASAP7_75t_R g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g643 ( .A(n_430), .Y(n_643) );
OR2x6_ASAP7_75t_L g901 ( .A(n_430), .B(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g597 ( .A(n_431), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_431), .B(n_973), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_434), .A2(n_707), .B1(n_936), .B2(n_938), .Y(n_951) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g581 ( .A(n_435), .Y(n_581) );
INVx2_ASAP7_75t_SL g988 ( .A(n_435), .Y(n_988) );
CKINVDCx6p67_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_438), .A2(n_503), .B(n_504), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_438), .A2(n_617), .B1(n_620), .B2(n_661), .C(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g515 ( .A(n_439), .Y(n_515) );
INVx1_ASAP7_75t_L g524 ( .A(n_439), .Y(n_524) );
BUFx4f_ASAP7_75t_L g910 ( .A(n_439), .Y(n_910) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
OR2x2_ASAP7_75t_L g497 ( .A(n_440), .B(n_441), .Y(n_497) );
XNOR2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_532), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_474), .C(n_487), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_467), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g477 ( .A(n_449), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g480 ( .A(n_449), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g484 ( .A(n_449), .B(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_449), .A2(n_466), .B1(n_555), .B2(n_562), .Y(n_554) );
AND2x4_ASAP7_75t_L g616 ( .A(n_449), .B(n_455), .Y(n_616) );
AND2x6_ASAP7_75t_L g618 ( .A(n_449), .B(n_473), .Y(n_618) );
AND2x4_ASAP7_75t_L g621 ( .A(n_449), .B(n_560), .Y(n_621) );
AND2x2_ASAP7_75t_L g623 ( .A(n_449), .B(n_478), .Y(n_623) );
AND2x2_ASAP7_75t_L g784 ( .A(n_449), .B(n_478), .Y(n_784) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_449), .B(n_478), .Y(n_1337) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_454), .B2(n_456), .C(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g736 ( .A(n_452), .Y(n_736) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g557 ( .A(n_455), .Y(n_557) );
BUFx3_ASAP7_75t_L g753 ( .A(n_455), .Y(n_753) );
INVx1_ASAP7_75t_L g889 ( .A(n_455), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_456), .A2(n_508), .B1(n_509), .B2(n_511), .Y(n_507) );
BUFx2_ASAP7_75t_L g776 ( .A(n_458), .Y(n_776) );
OAI33xp33_ASAP7_75t_L g733 ( .A1(n_459), .A2(n_734), .A3(n_740), .B1(n_745), .B2(n_747), .B3(n_751), .Y(n_733) );
OAI33xp33_ASAP7_75t_L g847 ( .A1(n_459), .A2(n_745), .A3(n_848), .B1(n_851), .B2(n_855), .B3(n_859), .Y(n_847) );
OAI33xp33_ASAP7_75t_L g1062 ( .A1(n_459), .A2(n_639), .A3(n_1063), .B1(n_1068), .B2(n_1073), .B3(n_1075), .Y(n_1062) );
OAI33xp33_ASAP7_75t_L g1342 ( .A1(n_459), .A2(n_745), .A3(n_1343), .B1(n_1347), .B2(n_1352), .B3(n_1353), .Y(n_1342) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .C(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g738 ( .A(n_464), .Y(n_738) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_464), .Y(n_768) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_468), .Y(n_730) );
INVx2_ASAP7_75t_L g1340 ( .A(n_468), .Y(n_1340) );
NAND2x1p5_ASAP7_75t_L g472 ( .A(n_469), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g536 ( .A(n_469), .B(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g539 ( .A(n_469), .B(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g543 ( .A(n_469), .B(n_544), .Y(n_543) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx4f_ASAP7_75t_L g731 ( .A(n_471), .Y(n_731) );
BUFx3_ASAP7_75t_L g732 ( .A(n_472), .Y(n_732) );
BUFx2_ASAP7_75t_L g1341 ( .A(n_472), .Y(n_1341) );
NOR2xp33_ASAP7_75t_SL g474 ( .A(n_475), .B(n_482), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_477), .A2(n_621), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g944 ( .A(n_477), .Y(n_944) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g945 ( .A(n_480), .Y(n_945) );
INVx2_ASAP7_75t_SL g631 ( .A(n_481), .Y(n_631) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_481), .Y(n_764) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g565 ( .A(n_485), .Y(n_565) );
INVx2_ASAP7_75t_L g853 ( .A(n_485), .Y(n_853) );
INVx2_ASAP7_75t_L g858 ( .A(n_485), .Y(n_858) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_485), .Y(n_929) );
INVx2_ASAP7_75t_L g553 ( .A(n_486), .Y(n_553) );
AND2x4_ASAP7_75t_L g642 ( .A(n_486), .B(n_643), .Y(n_642) );
OAI31xp33_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_495), .A3(n_501), .B(n_531), .Y(n_487) );
INVx1_ASAP7_75t_L g789 ( .A(n_489), .Y(n_789) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_490), .A2(n_820), .B1(n_823), .B2(n_825), .C(n_826), .Y(n_819) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_491), .A2(n_500), .B1(n_568), .B2(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g1024 ( .A(n_491), .Y(n_1024) );
BUFx4f_ASAP7_75t_L g1046 ( .A(n_491), .Y(n_1046) );
AND2x4_ASAP7_75t_L g499 ( .A(n_492), .B(n_500), .Y(n_499) );
AOI222xp33_ASAP7_75t_L g570 ( .A1(n_492), .A2(n_538), .B1(n_542), .B2(n_571), .C1(n_577), .C2(n_578), .Y(n_570) );
AND2x4_ASAP7_75t_L g648 ( .A(n_492), .B(n_649), .Y(n_648) );
INVx4_ASAP7_75t_L g681 ( .A(n_493), .Y(n_681) );
INVx1_ASAP7_75t_L g512 ( .A(n_494), .Y(n_512) );
INVx2_ASAP7_75t_L g807 ( .A(n_494), .Y(n_807) );
INVx6_ASAP7_75t_L g679 ( .A(n_496), .Y(n_679) );
INVx1_ASAP7_75t_L g510 ( .A(n_497), .Y(n_510) );
INVx1_ASAP7_75t_L g573 ( .A(n_497), .Y(n_573) );
INVx2_ASAP7_75t_L g662 ( .A(n_497), .Y(n_662) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_499), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_499), .A2(n_589), .B1(n_705), .B2(n_706), .C(n_710), .Y(n_704) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_499), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g828 ( .A1(n_499), .A2(n_589), .B1(n_829), .B2(n_831), .C(n_833), .Y(n_828) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_499), .Y(n_1041) );
AOI221xp5_ASAP7_75t_L g1311 ( .A1(n_499), .A2(n_589), .B1(n_1312), .B2(n_1313), .C(n_1314), .Y(n_1311) );
INVx2_ASAP7_75t_SL g583 ( .A(n_500), .Y(n_583) );
AND2x4_ASAP7_75t_L g589 ( .A(n_500), .B(n_530), .Y(n_589) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_500), .Y(n_670) );
BUFx4f_ASAP7_75t_L g707 ( .A(n_500), .Y(n_707) );
INVx1_ASAP7_75t_L g1045 ( .A(n_500), .Y(n_1045) );
OAI211xp5_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_507), .B(n_513), .C(n_521), .Y(n_501) );
INVx1_ASAP7_75t_L g672 ( .A(n_506), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g912 ( .A1(n_509), .A2(n_909), .B1(n_913), .B2(n_914), .C(n_915), .Y(n_912) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI211xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_516), .C(n_517), .Y(n_513) );
OAI211xp5_ASAP7_75t_L g794 ( .A1(n_515), .A2(n_780), .B(n_795), .C(n_796), .Y(n_794) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_518), .Y(n_587) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g592 ( .A(n_519), .Y(n_592) );
INVx2_ASAP7_75t_SL g797 ( .A(n_519), .Y(n_797) );
INVx1_ASAP7_75t_L g821 ( .A(n_519), .Y(n_821) );
INVx1_ASAP7_75t_L g965 ( .A(n_519), .Y(n_965) );
BUFx6f_ASAP7_75t_L g992 ( .A(n_519), .Y(n_992) );
NAND2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g957 ( .A(n_524), .Y(n_957) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_533), .B(n_600), .Y(n_532) );
INVx1_ASAP7_75t_L g602 ( .A(n_534), .Y(n_602) );
NAND3xp33_ASAP7_75t_SL g534 ( .A(n_535), .B(n_545), .C(n_554), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_538), .B1(n_539), .B2(n_542), .C(n_543), .Y(n_535) );
INVx1_ASAP7_75t_L g611 ( .A(n_536), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_536), .A2(n_539), .B1(n_543), .B2(n_758), .C(n_759), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_536), .A2(n_539), .B1(n_543), .B2(n_975), .C(n_976), .Y(n_974) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_539), .Y(n_608) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_543), .A2(n_608), .B1(n_609), .B2(n_610), .C(n_612), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_544), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_552), .B2(n_553), .Y(n_545) );
BUFx2_ASAP7_75t_L g761 ( .A(n_546), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_552), .A2(n_591), .B1(n_594), .B2(n_596), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_556), .A2(n_1008), .B1(n_1009), .B2(n_1010), .Y(n_1007) );
INVx2_ASAP7_75t_L g1070 ( .A(n_556), .Y(n_1070) );
INVx1_ASAP7_75t_L g772 ( .A(n_557), .Y(n_772) );
BUFx3_ASAP7_75t_L g629 ( .A(n_560), .Y(n_629) );
INVx1_ASAP7_75t_L g775 ( .A(n_560), .Y(n_775) );
BUFx3_ASAP7_75t_L g633 ( .A(n_563), .Y(n_633) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
AOI31xp33_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_579), .A3(n_590), .B(n_598), .Y(n_569) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g588 ( .A(n_574), .Y(n_588) );
INVx4_ASAP7_75t_L g792 ( .A(n_577), .Y(n_792) );
INVx2_ASAP7_75t_L g827 ( .A(n_577), .Y(n_827) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_578), .A2(n_652), .A3(n_696), .B1(n_698), .B2(n_701), .C1(n_702), .C2(n_703), .Y(n_695) );
INVx2_ASAP7_75t_SL g793 ( .A(n_578), .Y(n_793) );
INVx2_ASAP7_75t_L g1039 ( .A(n_578), .Y(n_1039) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_586), .B(n_589), .Y(n_579) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVxp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g1047 ( .A(n_585), .Y(n_1047) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_589), .A2(n_799), .B1(n_800), .B2(n_801), .C(n_803), .Y(n_798) );
INVx1_ASAP7_75t_L g952 ( .A(n_589), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g1040 ( .A1(n_589), .A2(n_1041), .B1(n_1042), .B2(n_1043), .C(n_1048), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_592), .A2(n_935), .B1(n_940), .B2(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g1325 ( .A(n_595), .Y(n_1325) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_599), .A2(n_719), .B1(n_818), .B2(n_837), .Y(n_817) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .C(n_603), .Y(n_600) );
INVx2_ASAP7_75t_L g685 ( .A(n_604), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_640), .Y(n_605) );
AND4x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_613), .C(n_619), .D(n_624), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_615), .A2(n_618), .B1(n_1326), .B2(n_1334), .Y(n_1333) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx2_ASAP7_75t_L g724 ( .A(n_616), .Y(n_724) );
BUFx2_ASAP7_75t_L g779 ( .A(n_616), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_616), .A2(n_618), .B1(n_841), .B2(n_842), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_616), .A2(n_618), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_618), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_618), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_621), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_621), .A2(n_623), .B1(n_844), .B2(n_845), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_621), .A2(n_623), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_621), .A2(n_1324), .B1(n_1336), .B2(n_1337), .Y(n_1335) );
AOI33xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_628), .A3(n_632), .B1(n_636), .B2(n_637), .B3(n_638), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI33xp33_ASAP7_75t_L g760 ( .A1(n_638), .A2(n_761), .A3(n_762), .B1(n_765), .B2(n_769), .B3(n_773), .Y(n_760) );
INVx1_ASAP7_75t_L g941 ( .A(n_638), .Y(n_941) );
INVx6_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx5_ASAP7_75t_L g746 ( .A(n_639), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .B(n_645), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_641), .A2(n_786), .B1(n_1310), .B2(n_1330), .Y(n_1309) );
INVx5_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_SL g719 ( .A(n_642), .Y(n_719) );
INVx2_ASAP7_75t_L g812 ( .A(n_642), .Y(n_812) );
AOI31xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_664), .A3(n_677), .B(n_682), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B(n_650), .C(n_655), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_648), .B(n_715), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g1032 ( .A1(n_648), .A2(n_1033), .B1(n_1034), .B2(n_1036), .C(n_1038), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_648), .B(n_1329), .Y(n_1328) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_SL g969 ( .A(n_652), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_652), .A2(n_1319), .B1(n_1320), .B2(n_1321), .Y(n_1318) );
INVx1_ASAP7_75t_SL g676 ( .A(n_654), .Y(n_676) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_659), .Y(n_824) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_661), .A2(n_892), .B1(n_895), .B2(n_909), .C(n_911), .Y(n_908) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g1022 ( .A(n_662), .Y(n_1022) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_667), .B2(n_673), .C(n_675), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_680), .B2(n_681), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_679), .A2(n_681), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_679), .A2(n_681), .B1(n_809), .B2(n_810), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_679), .A2(n_681), .B1(n_835), .B2(n_836), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_679), .A2(n_681), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_679), .A2(n_681), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
INVx1_ASAP7_75t_L g786 ( .A(n_682), .Y(n_786) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI31xp33_ASAP7_75t_L g947 ( .A1(n_683), .A2(n_948), .A3(n_953), .B(n_968), .Y(n_947) );
AOI21x1_ASAP7_75t_L g999 ( .A1(n_683), .A2(n_1000), .B(n_1011), .Y(n_999) );
XNOR2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_865), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_814), .B2(n_815), .Y(n_687) );
INVxp33_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
XNOR2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_754), .Y(n_689) );
XNOR2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_720), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_716), .B1(n_718), .B2(n_719), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_695), .B(n_704), .C(n_711), .D(n_714), .Y(n_694) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx3_ASAP7_75t_L g802 ( .A(n_700), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_705), .A2(n_712), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_713), .A2(n_715), .B1(n_735), .B2(n_752), .Y(n_751) );
CKINVDCx8_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
NOR3xp33_ASAP7_75t_SL g720 ( .A(n_721), .B(n_729), .C(n_733), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_726), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_735), .A2(n_852), .B1(n_853), .B2(n_854), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_735), .A2(n_825), .B1(n_836), .B2(n_856), .Y(n_855) );
BUFx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g939 ( .A(n_736), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_738), .A2(n_1069), .B1(n_1071), .B2(n_1072), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_740) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_743), .A2(n_748), .B1(n_849), .B2(n_850), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_743), .A2(n_893), .B1(n_931), .B2(n_932), .Y(n_930) );
CKINVDCx8_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
OAI22xp33_ASAP7_75t_L g859 ( .A1(n_748), .A2(n_833), .B1(n_835), .B2(n_860), .Y(n_859) );
OAI22xp33_ASAP7_75t_L g1063 ( .A1(n_748), .A2(n_1064), .B1(n_1065), .B2(n_1067), .Y(n_1063) );
OAI22xp33_ASAP7_75t_L g1075 ( .A1(n_748), .A2(n_862), .B1(n_1042), .B2(n_1050), .Y(n_1075) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_748), .A2(n_1344), .B1(n_1345), .B2(n_1346), .Y(n_1343) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g1345 ( .A(n_750), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_752), .A2(n_1033), .B1(n_1051), .B2(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
XNOR2x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_813), .Y(n_754) );
NAND2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_785), .Y(n_755) );
AND4x1_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .C(n_777), .D(n_781), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_763), .B(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B1(n_811), .B2(n_812), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_786), .A2(n_812), .B1(n_1031), .B2(n_1052), .Y(n_1030) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_798), .C(n_808), .Y(n_787) );
AOI21xp5_ASAP7_75t_SL g788 ( .A1(n_789), .A2(n_790), .B(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_SL g832 ( .A(n_806), .Y(n_832) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g863 ( .A(n_816), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_838), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_828), .C(n_834), .Y(n_818) );
NOR3xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_846), .C(n_847), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
INVx2_ASAP7_75t_SL g1350 ( .A(n_853), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_853), .A2(n_1074), .B1(n_1317), .B2(n_1329), .Y(n_1352) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_979), .B1(n_980), .B2(n_1078), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g1079 ( .A(n_867), .Y(n_1079) );
XNOR2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_922), .Y(n_867) );
INVx1_ASAP7_75t_L g920 ( .A(n_869), .Y(n_920) );
NAND4xp25_ASAP7_75t_L g869 ( .A(n_870), .B(n_899), .C(n_903), .D(n_916), .Y(n_869) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_884), .B(n_898), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_878), .B(n_880), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_886), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
BUFx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx3_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
OAI21xp5_ASAP7_75t_L g1003 ( .A1(n_897), .A2(n_1004), .B(n_1007), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
INVx3_ASAP7_75t_L g986 ( .A(n_906), .Y(n_986) );
INVx2_ASAP7_75t_SL g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g963 ( .A(n_910), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_921), .A2(n_1083), .B1(n_1104), .B2(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_SL g978 ( .A(n_923), .Y(n_978) );
NAND4xp75_ASAP7_75t_L g923 ( .A(n_924), .B(n_942), .C(n_947), .D(n_974), .Y(n_923) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g962 ( .A1(n_932), .A2(n_963), .B(n_964), .C(n_966), .Y(n_962) );
INVx1_ASAP7_75t_L g1355 ( .A(n_934), .Y(n_1355) );
NOR2x1_ASAP7_75t_L g942 ( .A(n_943), .B(n_946), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_954), .B(n_962), .Y(n_953) );
OAI211xp5_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_956), .B(n_958), .C(n_959), .Y(n_954) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx3_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
AO22x2_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_1027), .B1(n_1028), .B2(n_1077), .Y(n_980) );
INVxp67_ASAP7_75t_SL g1077 ( .A(n_981), .Y(n_1077) );
INVxp67_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
NOR4xp75_ASAP7_75t_L g983 ( .A(n_984), .B(n_999), .C(n_1020), .D(n_1025), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_995), .Y(n_984) );
AOI33xp33_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_987), .A3(n_989), .B1(n_990), .B2(n_993), .B3(n_994), .Y(n_985) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g1035 ( .A(n_992), .Y(n_1035) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
XOR2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1076), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1053), .Y(n_1029) );
NAND3xp33_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1040), .C(n_1049), .Y(n_1031) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1037), .Y(n_1323) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NOR3xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1061), .C(n_1062), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1058), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1353 ( .A1(n_1065), .A2(n_1312), .B1(n_1316), .B2(n_1354), .Y(n_1353) );
INVx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_1069), .A2(n_1348), .B1(n_1349), .B2(n_1351), .Y(n_1347) );
INVx2_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1070), .Y(n_1074) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1089), .B1(n_1306), .B2(n_1356), .C(n_1360), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_1081), .A2(n_1194), .B1(n_1195), .B2(n_1196), .Y(n_1193) );
BUFx3_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g1101 ( .A1(n_1082), .A2(n_1102), .B1(n_1103), .B2(n_1104), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_1082), .A2(n_1104), .B1(n_1141), .B2(n_1142), .Y(n_1140) );
OAI22xp33_ASAP7_75t_L g1152 ( .A1(n_1082), .A2(n_1153), .B1(n_1154), .B2(n_1155), .Y(n_1152) );
BUFx6f_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1084), .B(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1084), .Y(n_1110) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1085), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1088), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1088), .Y(n_1098) );
NOR2x1_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1243), .Y(n_1089) );
NAND3xp33_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1181), .C(n_1204), .Y(n_1090) );
AOI211xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1115), .B(n_1143), .C(n_1173), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1092), .B(n_1164), .Y(n_1246) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_1093), .A2(n_1106), .B1(n_1284), .B2(n_1285), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1106), .Y(n_1093) );
INVx2_ASAP7_75t_SL g1169 ( .A(n_1094), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1094), .B(n_1128), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1094), .B(n_1106), .Y(n_1252) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_1095), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1148 ( .A(n_1095), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1095), .B(n_1106), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1095), .B(n_1106), .Y(n_1225) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1096), .Y(n_1159) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1096), .Y(n_1191) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1099), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1097), .B(n_1099), .Y(n_1114) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
AND2x4_ASAP7_75t_L g1100 ( .A(n_1098), .B(n_1099), .Y(n_1100) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1100), .Y(n_1132) );
INVx1_ASAP7_75t_SL g1138 ( .A(n_1100), .Y(n_1138) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1104), .Y(n_1156) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1105), .Y(n_1112) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1106), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1106), .B(n_1150), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_1106), .B(n_1150), .Y(n_1201) );
OAI21xp33_ASAP7_75t_L g1205 ( .A1(n_1106), .A2(n_1206), .B(n_1208), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1106), .B(n_1151), .Y(n_1236) );
AND2x4_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1113), .Y(n_1106) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_1109), .B(n_1110), .Y(n_1108) );
OAI21xp33_ASAP7_75t_SL g1368 ( .A1(n_1109), .A2(n_1364), .B(n_1369), .Y(n_1368) );
AND2x4_ASAP7_75t_L g1111 ( .A(n_1110), .B(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1114), .Y(n_1136) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1126), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1117), .B(n_1227), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1237 ( .A(n_1117), .B(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1118), .B(n_1133), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1118), .B(n_1134), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1122), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1119), .B(n_1123), .Y(n_1146) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1119), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1119), .B(n_1134), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1119), .B(n_1123), .Y(n_1265) );
NOR2xp33_ASAP7_75t_SL g1295 ( .A(n_1119), .B(n_1296), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1166 ( .A(n_1122), .B(n_1133), .Y(n_1166) );
NOR3xp33_ASAP7_75t_L g1186 ( .A(n_1122), .B(n_1164), .C(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1122), .B(n_1133), .Y(n_1216) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1123), .B(n_1133), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1123), .B(n_1179), .Y(n_1178) );
OAI322xp33_ASAP7_75t_L g1249 ( .A1(n_1123), .A2(n_1250), .A3(n_1253), .B1(n_1254), .B2(n_1256), .C1(n_1258), .C2(n_1260), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1123), .B(n_1133), .Y(n_1259) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1133), .Y(n_1127) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1128), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1128), .B(n_1133), .Y(n_1180) );
INVx4_ASAP7_75t_L g1185 ( .A(n_1128), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_1128), .B(n_1215), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1128), .B(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1128), .B(n_1255), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1128), .B(n_1151), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1128), .B(n_1169), .Y(n_1296) );
AND2x6_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1130), .Y(n_1128) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_1132), .A2(n_1190), .B1(n_1191), .B2(n_1192), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1133), .B(n_1146), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1133), .B(n_1184), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1133), .B(n_1178), .Y(n_1239) );
CKINVDCx6p67_ASAP7_75t_R g1133 ( .A(n_1134), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1134), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1134), .B(n_1178), .Y(n_1219) );
AOI32xp33_ASAP7_75t_L g1221 ( .A1(n_1134), .A2(n_1200), .A3(n_1222), .B1(n_1226), .B2(n_1228), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1134), .B(n_1146), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1264 ( .A(n_1134), .B(n_1265), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1134), .B(n_1294), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1134), .B(n_1300), .Y(n_1299) );
OR2x6_ASAP7_75t_SL g1134 ( .A(n_1135), .B(n_1140), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_1136), .A2(n_1137), .B1(n_1138), .B2(n_1139), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1157 ( .A1(n_1138), .A2(n_1158), .B1(n_1159), .B2(n_1160), .Y(n_1157) );
OAI221xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1147), .B1(n_1162), .B2(n_1167), .C(n_1170), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1146), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1146), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1148), .Y(n_1278) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1148), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1149), .B(n_1171), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1161), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1150), .B(n_1169), .Y(n_1168) );
INVx3_ASAP7_75t_L g1213 ( .A(n_1150), .Y(n_1213) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1150), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1150), .B(n_1197), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1150), .B(n_1188), .Y(n_1253) );
INVx3_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_1151), .B(n_1225), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1157), .Y(n_1151) );
HB1xp67_ASAP7_75t_L g1196 ( .A(n_1155), .Y(n_1196) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
NOR2x1_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1166), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1164), .B(n_1219), .Y(n_1218) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1164), .B(n_1271), .Y(n_1270) );
NOR2x1_ASAP7_75t_R g1286 ( .A(n_1164), .B(n_1227), .Y(n_1286) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1165), .B(n_1172), .Y(n_1171) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1165), .B(n_1215), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1165), .B(n_1231), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1165), .B(n_1219), .Y(n_1304) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1166), .Y(n_1233) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
AOI322xp5_ASAP7_75t_L g1232 ( .A1(n_1168), .A2(n_1213), .A3(n_1233), .B1(n_1234), .B2(n_1236), .C1(n_1237), .C2(n_1239), .Y(n_1232) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1169), .Y(n_1175) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1169), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1169), .B(n_1236), .Y(n_1257) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1169), .Y(n_1273) );
NOR2xp33_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1177), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1176), .Y(n_1174) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1176), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1180), .Y(n_1177) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1178), .Y(n_1227) );
AOI211xp5_ASAP7_75t_L g1281 ( .A1(n_1179), .A2(n_1282), .B(n_1283), .C(n_1286), .Y(n_1281) );
O2A1O1Ixp33_ASAP7_75t_L g1181 ( .A1(n_1182), .A2(n_1186), .B(n_1197), .C(n_1198), .Y(n_1181) );
INVxp67_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1185), .B(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1185), .Y(n_1210) );
NOR2xp33_ASAP7_75t_L g1300 ( .A(n_1185), .B(n_1265), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1185), .B(n_1224), .Y(n_1302) );
OAI31xp33_ASAP7_75t_L g1204 ( .A1(n_1187), .A2(n_1205), .A3(n_1217), .B(n_1220), .Y(n_1204) );
OAI221xp5_ASAP7_75t_L g1291 ( .A1(n_1187), .A2(n_1225), .B1(n_1292), .B2(n_1297), .C(n_1301), .Y(n_1291) );
CKINVDCx5p33_ASAP7_75t_R g1187 ( .A(n_1188), .Y(n_1187) );
AOI22xp5_ASAP7_75t_L g1266 ( .A1(n_1188), .A2(n_1267), .B1(n_1276), .B2(n_1277), .Y(n_1266) );
OR2x6_ASAP7_75t_SL g1188 ( .A(n_1189), .B(n_1193), .Y(n_1188) );
XNOR2x1_ASAP7_75t_L g1307 ( .A(n_1194), .B(n_1308), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1197), .B(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1202), .Y(n_1199) );
AOI322xp5_ASAP7_75t_L g1292 ( .A1(n_1200), .A2(n_1213), .A3(n_1216), .B1(n_1251), .B2(n_1252), .C1(n_1293), .C2(n_1295), .Y(n_1292) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1202), .B(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1203), .Y(n_1229) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
OAI21xp5_ASAP7_75t_SL g1208 ( .A1(n_1209), .A2(n_1211), .B(n_1216), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1210), .B(n_1231), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1214), .Y(n_1211) );
INVx1_ASAP7_75t_SL g1212 ( .A(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1213), .B(n_1218), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1213), .B(n_1239), .Y(n_1275) );
AOI21xp5_ASAP7_75t_L g1274 ( .A1(n_1214), .A2(n_1227), .B(n_1268), .Y(n_1274) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1214), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1216), .B(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1219), .Y(n_1248) );
NAND3xp33_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1232), .C(n_1240), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1224), .B(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1230), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1229), .B(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1231), .Y(n_1268) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
A2O1A1Ixp33_ASAP7_75t_L g1288 ( .A1(n_1235), .A2(n_1248), .B(n_1264), .C(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1236), .Y(n_1271) );
AOI211xp5_ASAP7_75t_SL g1287 ( .A1(n_1236), .A2(n_1288), .B(n_1291), .C(n_1303), .Y(n_1287) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1238), .Y(n_1290) );
NOR2xp33_ASAP7_75t_L g1258 ( .A(n_1239), .B(n_1259), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1239), .B(n_1273), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1239), .B(n_1290), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1242), .Y(n_1240) );
AOI211xp5_ASAP7_75t_L g1269 ( .A1(n_1241), .A2(n_1270), .B(n_1272), .C(n_1274), .Y(n_1269) );
NAND3xp33_ASAP7_75t_L g1243 ( .A(n_1244), .B(n_1266), .C(n_1287), .Y(n_1243) );
AOI211xp5_ASAP7_75t_SL g1244 ( .A1(n_1245), .A2(n_1247), .B(n_1249), .C(n_1262), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1245 ( .A(n_1246), .Y(n_1245) );
OAI211xp5_ASAP7_75t_L g1277 ( .A1(n_1248), .A2(n_1278), .B(n_1279), .C(n_1281), .Y(n_1277) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1253), .Y(n_1276) );
OAI211xp5_ASAP7_75t_L g1267 ( .A1(n_1256), .A2(n_1268), .B(n_1269), .C(n_1275), .Y(n_1267) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1264), .Y(n_1262) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1265), .Y(n_1294) );
AOI21xp5_ASAP7_75t_L g1303 ( .A1(n_1297), .A2(n_1304), .B(n_1305), .Y(n_1303) );
INVxp67_ASAP7_75t_SL g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx2_ASAP7_75t_SL g1306 ( .A(n_1307), .Y(n_1306) );
HB1xp67_ASAP7_75t_L g1367 ( .A(n_1308), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1331), .Y(n_1308) );
NAND5xp2_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1315), .C(n_1318), .D(n_1322), .E(n_1328), .Y(n_1310) );
OAI221xp5_ASAP7_75t_SL g1322 ( .A1(n_1323), .A2(n_1324), .B1(n_1325), .B2(n_1326), .C(n_1327), .Y(n_1322) );
NOR3xp33_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1338), .C(n_1342), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1335), .Y(n_1332) );
INVx2_ASAP7_75t_SL g1339 ( .A(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx4_ASAP7_75t_SL g1356 ( .A(n_1357), .Y(n_1356) );
BUFx3_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
BUFx2_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
CKINVDCx5p33_ASAP7_75t_R g1362 ( .A(n_1363), .Y(n_1362) );
INVxp33_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
endmodule