module fake_jpeg_143_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_15),
.B(n_32),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_21),
.B(n_27),
.C(n_26),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_36),
.A3(n_32),
.B1(n_35),
.B2(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_16),
.B1(n_27),
.B2(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_48),
.B1(n_62),
.B2(n_0),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_16),
.B1(n_21),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_24),
.B1(n_19),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_57),
.B1(n_45),
.B2(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_24),
.B1(n_19),
.B2(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_15),
.B1(n_25),
.B2(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_42),
.B1(n_39),
.B2(n_30),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_69),
.B1(n_74),
.B2(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_64),
.B(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_29),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_4),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_12),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_12),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_7),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_60),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_78),
.B(n_79),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_0),
.B1(n_1),
.B2(n_9),
.Y(n_77)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_51),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_64),
.B(n_76),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_43),
.B(n_55),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_80),
.B(n_63),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_94),
.B1(n_82),
.B2(n_88),
.Y(n_103)
);

FAx1_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_61),
.CI(n_54),
.CON(n_88),
.SN(n_88)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_85),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_76),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_83),
.B(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_75),
.B1(n_67),
.B2(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_102),
.B(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_101),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_103),
.B1(n_100),
.B2(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_117),
.B(n_120),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_100),
.C(n_98),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_114),
.C(n_111),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_84),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_119),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_127),
.Y(n_130)
);

AOI21x1_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_120),
.B(n_117),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_129),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_121),
.B(n_128),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_131),
.B(n_124),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.Y(n_134)
);


endmodule