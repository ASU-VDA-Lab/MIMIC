module fake_jpeg_25663_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_21),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_41),
.B(n_37),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_29),
.B1(n_16),
.B2(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_16),
.B1(n_29),
.B2(n_20),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_20),
.B1(n_25),
.B2(n_27),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_57),
.Y(n_77)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_62),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_71),
.B1(n_74),
.B2(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_70),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_25),
.B1(n_39),
.B2(n_35),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_25),
.B1(n_39),
.B2(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx2_ASAP7_75t_SL g107 ( 
.A(n_76),
.Y(n_107)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_57),
.B1(n_51),
.B2(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_38),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_39),
.B1(n_17),
.B2(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_54),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_60),
.B1(n_47),
.B2(n_52),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_95),
.B1(n_97),
.B2(n_101),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_60),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_104),
.B(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_52),
.B1(n_58),
.B2(n_46),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_65),
.A2(n_52),
.B1(n_46),
.B2(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_109),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_41),
.C(n_37),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_106),
.C(n_110),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_70),
.A2(n_85),
.B1(n_83),
.B2(n_80),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_88),
.B1(n_98),
.B2(n_103),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_45),
.A3(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_41),
.C(n_54),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_66),
.A3(n_64),
.B1(n_76),
.B2(n_62),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_54),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_54),
.C(n_42),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_57),
.B1(n_51),
.B2(n_17),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_79),
.B1(n_42),
.B2(n_24),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_32),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_82),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_120),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_0),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_78),
.B1(n_72),
.B2(n_67),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_131),
.B1(n_135),
.B2(n_88),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_72),
.B1(n_67),
.B2(n_28),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_124),
.B1(n_133),
.B2(n_134),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_31),
.B(n_28),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_18),
.B(n_19),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_21),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_92),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_24),
.B1(n_23),
.B2(n_17),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_24),
.B1(n_79),
.B2(n_30),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_42),
.B1(n_30),
.B2(n_32),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_114),
.Y(n_160)
);

OAI22x1_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_32),
.B1(n_18),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_138),
.A2(n_106),
.B1(n_102),
.B2(n_110),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_139),
.A2(n_125),
.B1(n_129),
.B2(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_0),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_141),
.A2(n_161),
.B(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_151),
.B1(n_155),
.B2(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_111),
.B1(n_108),
.B2(n_97),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_89),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_156),
.C(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_160),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_111),
.C(n_101),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_2),
.C(n_3),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_113),
.C(n_112),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_103),
.B1(n_98),
.B2(n_105),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_169),
.B1(n_140),
.B2(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_82),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_19),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_18),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_168),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_0),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_1),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_18),
.B1(n_19),
.B2(n_4),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_166),
.B1(n_165),
.B2(n_147),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_114),
.C(n_126),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_116),
.C(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_178),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_122),
.B1(n_124),
.B2(n_131),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_143),
.B1(n_145),
.B2(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_121),
.B1(n_135),
.B2(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_133),
.B1(n_18),
.B2(n_19),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_163),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_189),
.B1(n_193),
.B2(n_11),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_195),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_146),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_198),
.B1(n_14),
.B2(n_12),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_8),
.B(n_9),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_161),
.B(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_202),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_205),
.B1(n_219),
.B2(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_160),
.B1(n_170),
.B2(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_196),
.A2(n_161),
.B1(n_156),
.B2(n_159),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_156),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_206),
.B(n_213),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_191),
.A2(n_147),
.B(n_153),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_142),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_214),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_142),
.B1(n_10),
.B2(n_11),
.Y(n_215)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_215),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_8),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_221),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_11),
.Y(n_221)
);

NAND4xp25_ASAP7_75t_SL g222 ( 
.A(n_190),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_187),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_198),
.B1(n_192),
.B2(n_197),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_176),
.C(n_175),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_229),
.C(n_233),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_184),
.C(n_186),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_184),
.C(n_186),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_180),
.C(n_185),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_240),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_185),
.C(n_182),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_241),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_216),
.B1(n_210),
.B2(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_217),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_255),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_200),
.B1(n_203),
.B2(n_216),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_251),
.A2(n_253),
.B1(n_230),
.B2(n_219),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_205),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_254),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_211),
.B1(n_209),
.B2(n_179),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_212),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_212),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_258),
.A2(n_224),
.B(n_227),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_224),
.B(n_235),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_259),
.A2(n_202),
.B(n_194),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_238),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_177),
.Y(n_281)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_270),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_265),
.B(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_229),
.C(n_236),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_268),
.C(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_228),
.C(n_241),
.Y(n_268)
);

XOR2x2_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_191),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_262),
.C(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_276),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_248),
.B1(n_253),
.B2(n_237),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_282),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_260),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_177),
.C(n_195),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_261),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_288),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_183),
.Y(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_270),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_260),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_280),
.B(n_272),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_292),
.C(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_291),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_274),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_297),
.B(n_287),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_299),
.A2(n_300),
.B(n_301),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_302),
.A2(n_295),
.B(n_296),
.Y(n_303)
);

OAI321xp33_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_298),
.A3(n_294),
.B1(n_223),
.B2(n_193),
.C(n_189),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_222),
.B1(n_199),
.B2(n_14),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_305),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_13),
.B1(n_14),
.B2(n_296),
.Y(n_307)
);


endmodule