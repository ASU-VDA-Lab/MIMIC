module fake_jpeg_28544_n_93 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_31),
.B1(n_33),
.B2(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_38),
.B1(n_37),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_1),
.Y(n_55)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_62),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_13),
.B1(n_29),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_56),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_6),
.B(n_7),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_11),
.B1(n_26),
.B2(n_24),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_5),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_52),
.B1(n_46),
.B2(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_61),
.B1(n_46),
.B2(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_6),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_14),
.C(n_30),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_74),
.B1(n_73),
.B2(n_71),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_77),
.B(n_69),
.C(n_80),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_80),
.C(n_84),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_84),
.A3(n_82),
.B1(n_85),
.B2(n_46),
.C1(n_23),
.C2(n_10),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_9),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_7),
.B(n_8),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);


endmodule