module fake_netlist_5_1279_n_77 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_77);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_77;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_38;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_0),
.A2(n_14),
.B1(n_21),
.B2(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_6),
.B(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_25),
.C(n_31),
.Y(n_43)
);

OAI22x1_ASAP7_75t_R g44 ( 
.A1(n_24),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_26),
.B(n_5),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_36),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AO21x1_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_30),
.B(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_58),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_46),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_SL g67 ( 
.A(n_66),
.B(n_62),
.C(n_61),
.Y(n_67)
);

NOR4xp25_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_39),
.C(n_63),
.D(n_66),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_63),
.B1(n_55),
.B2(n_60),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_64),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_59),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_39),
.C(n_30),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_60),
.B1(n_45),
.B2(n_23),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_60),
.B1(n_65),
.B2(n_26),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_12),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_26),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_27),
.Y(n_77)
);


endmodule