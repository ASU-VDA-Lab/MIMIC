module fake_jpeg_1832_n_93 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_31),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_27),
.Y(n_44)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_37),
.B1(n_34),
.B2(n_35),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_43),
.B1(n_40),
.B2(n_39),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_29),
.B1(n_26),
.B2(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_22),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_27),
.C(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_36),
.B1(n_33),
.B2(n_25),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_38),
.C(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_56),
.B(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_58),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_30),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_1),
.B(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_50),
.B1(n_30),
.B2(n_3),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_65),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_20),
.C(n_17),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_54),
.B(n_7),
.Y(n_76)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_61),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_78),
.B(n_8),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_12),
.C(n_13),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.C(n_84),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_79),
.B(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_86),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_85),
.B(n_14),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_15),
.C(n_10),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_11),
.Y(n_93)
);


endmodule