module fake_jpeg_24853_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_45),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_32),
.B1(n_25),
.B2(n_21),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_58),
.B1(n_61),
.B2(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_51),
.B1(n_67),
.B2(n_71),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_26),
.B1(n_30),
.B2(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_33),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_64),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_21),
.B1(n_24),
.B2(n_22),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_30),
.B1(n_45),
.B2(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_20),
.B1(n_24),
.B2(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_24),
.B1(n_33),
.B2(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_95),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

OR2x4_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_17),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_77),
.A2(n_83),
.B(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_82),
.A2(n_101),
.B1(n_54),
.B2(n_41),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_41),
.C(n_39),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_41),
.Y(n_131)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_19),
.Y(n_91)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_19),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_34),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_58),
.B(n_35),
.C(n_34),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_100),
.Y(n_121)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_102),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_31),
.B(n_23),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_62),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_13),
.Y(n_104)
);

XOR2x2_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_106),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_13),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_27),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_107),
.B(n_88),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_117),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_49),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_131),
.C(n_84),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_59),
.B1(n_47),
.B2(n_49),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_122),
.B1(n_123),
.B2(n_97),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_49),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_113),
.Y(n_142)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_76),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_125),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_47),
.B1(n_52),
.B2(n_22),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_22),
.B1(n_34),
.B2(n_27),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_97),
.B1(n_93),
.B2(n_103),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_83),
.A2(n_31),
.B1(n_29),
.B2(n_39),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_82),
.B1(n_101),
.B2(n_73),
.Y(n_152)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_140),
.B(n_144),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_99),
.B(n_103),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_142),
.B(n_150),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_74),
.C(n_89),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_156),
.C(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_149),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_98),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_87),
.B(n_73),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_160),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_104),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_106),
.C(n_93),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_79),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_78),
.B1(n_72),
.B2(n_92),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_100),
.B1(n_75),
.B2(n_102),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_168),
.B1(n_122),
.B2(n_114),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_14),
.B(n_8),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_9),
.B(n_16),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_133),
.B(n_80),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_9),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_75),
.C(n_108),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_7),
.C(n_15),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_31),
.B1(n_29),
.B2(n_54),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_115),
.A2(n_29),
.B1(n_39),
.B2(n_36),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_119),
.B1(n_120),
.B2(n_114),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_118),
.A3(n_130),
.B1(n_123),
.B2(n_137),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_179),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_113),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_178),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_151),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_133),
.B(n_135),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_190),
.B(n_149),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_189),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_109),
.B1(n_119),
.B2(n_136),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_109),
.B1(n_136),
.B2(n_116),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_116),
.B1(n_120),
.B2(n_41),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_152),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_143),
.A2(n_39),
.B1(n_36),
.B2(n_124),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_124),
.B1(n_36),
.B2(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_36),
.B1(n_124),
.B2(n_2),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_138),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_201),
.C(n_9),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_0),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_200),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_8),
.Y(n_200)
);

OA21x2_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_229),
.B(n_190),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_174),
.A2(n_150),
.B(n_144),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_221),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_140),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_191),
.A2(n_163),
.B1(n_175),
.B2(n_188),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_218),
.B1(n_199),
.B2(n_1),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_138),
.B1(n_146),
.B2(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_186),
.B1(n_185),
.B2(n_179),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_169),
.B1(n_155),
.B2(n_168),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_148),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_220),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_145),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_200),
.C(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_186),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_148),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_7),
.Y(n_229)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_232),
.B(n_13),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_178),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_215),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_245),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_185),
.B1(n_201),
.B2(n_187),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_247),
.B1(n_251),
.B2(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_246),
.C(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_210),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_172),
.C(n_173),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_196),
.B1(n_176),
.B2(n_195),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_220),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_205),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_173),
.C(n_171),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_207),
.B1(n_213),
.B2(n_206),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_252),
.A2(n_267),
.B1(n_268),
.B2(n_251),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_230),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_256),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_204),
.Y(n_256)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_235),
.B(n_229),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_269),
.B(n_242),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_218),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_224),
.C(n_226),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_240),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_237),
.A2(n_208),
.B1(n_203),
.B2(n_212),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_203),
.B1(n_212),
.B2(n_211),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_205),
.B1(n_209),
.B2(n_4),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_235),
.B(n_249),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_231),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_231),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_234),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_276),
.C(n_282),
.Y(n_295)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_278),
.B1(n_281),
.B2(n_233),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_238),
.Y(n_276)
);

AOI21x1_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_266),
.B(n_264),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_277),
.A2(n_253),
.B1(n_233),
.B2(n_243),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_261),
.B1(n_257),
.B2(n_241),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_252),
.B1(n_230),
.B2(n_262),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_271),
.C(n_272),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_267),
.B1(n_14),
.B2(n_11),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_16),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_15),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_15),
.B(n_16),
.Y(n_296)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_304),
.B(n_289),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_295),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_5),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_6),
.B(n_291),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_295),
.B(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.C(n_311),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_286),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_310),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_287),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_288),
.C(n_292),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_290),
.C(n_300),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_300),
.B(n_307),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_312),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_318),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_317),
.Y(n_320)
);


endmodule