module real_jpeg_32689_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_0),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_0),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_100),
.B1(n_104),
.B2(n_109),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_1),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_1),
.A2(n_109),
.B1(n_234),
.B2(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_1),
.A2(n_109),
.B1(n_407),
.B2(n_411),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_2),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_2),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_2),
.A2(n_54),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_2),
.A2(n_54),
.B1(n_177),
.B2(n_181),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_2),
.A2(n_54),
.B1(n_372),
.B2(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_24),
.B1(n_134),
.B2(n_139),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_3),
.B(n_192),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_3),
.A2(n_205),
.B(n_243),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_3),
.B(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_4),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_4),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_76),
.B1(n_80),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_7),
.A2(n_82),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_9),
.A2(n_122),
.B1(n_123),
.B2(n_128),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_9),
.A2(n_122),
.B1(n_219),
.B2(n_223),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_9),
.A2(n_122),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_11),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_12),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_12),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_13),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_14),
.A2(n_337),
.B1(n_338),
.B2(n_340),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_14),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_324),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_226),
.B(n_323),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_171),
.Y(n_18)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_19),
.B(n_171),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_131),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_21),
.B(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_22),
.B(n_46),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_38),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_39),
.C(n_43),
.Y(n_38)
);

NOR2xp67_ASAP7_75t_R g246 ( 
.A(n_24),
.B(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_24),
.B(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_24),
.A2(n_271),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_24),
.B(n_248),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_24),
.B(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_24),
.A2(n_393),
.B(n_397),
.Y(n_392)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_28),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_28),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_31),
.A2(n_146),
.B1(n_154),
.B2(n_157),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_32),
.Y(n_140)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_37),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_37),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_41),
.Y(n_165)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_42),
.Y(n_224)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_43),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_67),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_47),
.A2(n_293),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_61),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_48),
.B(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_58),
.Y(n_341)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_59),
.Y(n_237)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_60),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_60),
.Y(n_268)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_61),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_61),
.A2(n_287),
.B1(n_291),
.B2(n_292),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_61),
.A2(n_68),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_64),
.Y(n_339)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_65),
.Y(n_214)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g245 ( 
.A(n_66),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_75),
.A2(n_205),
.B1(n_206),
.B2(n_213),
.Y(n_204)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_85),
.B(n_132),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_98),
.B1(n_110),
.B2(n_120),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_88),
.Y(n_184)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_94),
.B2(n_96),
.Y(n_88)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_90),
.Y(n_317)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_95),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_113),
.B1(n_115),
.B2(n_117),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_97),
.Y(n_270)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_99),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_103),
.Y(n_402)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_110),
.B(n_275),
.Y(n_274)
);

AO22x1_ASAP7_75t_L g399 ( 
.A1(n_110),
.A2(n_176),
.B1(n_184),
.B2(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_111),
.A2(n_121),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

BUFx4f_ASAP7_75t_SL g259 ( 
.A(n_113),
.Y(n_259)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_119),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_141),
.B(n_160),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_137),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_140),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_140),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_142),
.B(n_162),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_142),
.A2(n_218),
.B1(n_405),
.B2(n_413),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

AOI22x1_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_151),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_188),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_175),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.Y(n_175)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_179),
.Y(n_403)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_185),
.B(n_186),
.C(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_188),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_215),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_203),
.B2(n_204),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_190),
.B(n_204),
.C(n_215),
.Y(n_367)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_192),
.B(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_193),
.B(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_201),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_198),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_198),
.Y(n_365)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_198),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_198),
.Y(n_391)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_233),
.B(n_243),
.Y(n_232)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_206),
.Y(n_335)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_SL g296 ( 
.A(n_212),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B(n_225),
.Y(n_215)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_216),
.Y(n_413)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_282),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_250),
.B(n_281),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_229),
.B(n_231),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.C(n_247),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_247),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_277),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_273),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_252),
.A2(n_273),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

AO221x1_ASAP7_75t_L g319 ( 
.A1(n_252),
.A2(n_273),
.B1(n_286),
.B2(n_299),
.C(n_300),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_257),
.B(n_265),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_269),
.B(n_271),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_283),
.C(n_320),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_301),
.B(n_319),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_298),
.Y(n_285)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_309),
.B(n_318),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_304),
.B(n_305),
.Y(n_318)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_414),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_328),
.B(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_368),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_366),
.B2(n_367),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_342),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI32xp33_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_350),
.A3(n_353),
.B1(n_356),
.B2(n_362),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_355),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_355),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_355),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_356),
.Y(n_397)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_358),
.A2(n_383),
.B1(n_385),
.B2(n_389),
.Y(n_382)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_398),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_380),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_376),
.Y(n_384)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_392),
.Y(n_380)
);

INVx4_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx11_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx12f_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);


endmodule