module fake_jpeg_30993_n_16 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_16);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_16;

wire n_13;
wire n_11;
wire n_14;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx2_ASAP7_75t_SL g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_L g10 ( 
.A1(n_8),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_10)
);

AOI31xp67_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_12),
.A3(n_0),
.B(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

AOI322xp5_ASAP7_75t_L g15 ( 
.A1(n_14),
.A2(n_10),
.A3(n_12),
.B1(n_9),
.B2(n_5),
.C1(n_3),
.C2(n_4),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_13),
.C(n_4),
.Y(n_16)
);


endmodule