module fake_jpeg_21428_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx11_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_2),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx4f_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_0),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_16),
.Y(n_19)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_21),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_6),
.Y(n_26)
);

NOR4xp25_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_12),
.C(n_15),
.D(n_10),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_20),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_30),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_24),
.C(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_7),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_34),
.B1(n_21),
.B2(n_0),
.Y(n_36)
);


endmodule