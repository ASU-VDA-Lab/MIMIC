module fake_netlist_6_1455_n_1932 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1932);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1932;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_8),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_13),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_67),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_25),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_10),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_0),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_26),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_132),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_168),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_90),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_54),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_91),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_114),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_7),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_96),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_73),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_72),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_68),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_115),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_121),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_126),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_80),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_95),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_23),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_61),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_24),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_102),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_99),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_64),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_19),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_41),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_176),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_137),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_37),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_79),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_131),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_112),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_65),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_98),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_15),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_148),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_21),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_13),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_19),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_94),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_42),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_60),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_60),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_70),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_149),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_77),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_46),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_49),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_31),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_173),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_2),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_54),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_134),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_123),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_89),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_106),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_56),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_76),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_16),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_33),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_133),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_30),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_117),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_152),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_17),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_45),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_11),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_71),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_57),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_124),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_66),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_154),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_82),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_50),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_56),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_1),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_129),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_160),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_22),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_44),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_119),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_26),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_100),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_41),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_101),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_30),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_165),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_113),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_103),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_74),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_50),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_35),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_24),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_21),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_88),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_128),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_69),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_97),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_36),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_155),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_164),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_83),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_3),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_143),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_146),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_3),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_10),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_111),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_62),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_2),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_140),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_58),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_105),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_47),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_16),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_178),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_170),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_57),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_180),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_31),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_36),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_84),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_92),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_145),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_120),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_153),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_28),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_45),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_28),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_4),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_37),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_86),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_17),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_35),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_7),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_29),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_118),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_12),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_55),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_33),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_167),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_23),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_174),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_59),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_104),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_43),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_58),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_14),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_15),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_52),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_181),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_144),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_22),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_39),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_330),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_320),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_222),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_196),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_364),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_242),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_334),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_203),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_183),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_223),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_183),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_220),
.B(n_4),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_227),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_254),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_187),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_333),
.B(n_228),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_356),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_5),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_356),
.B(n_5),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_230),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_217),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_316),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_273),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_6),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g397 ( 
.A(n_187),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_273),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_317),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_231),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_232),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_273),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_273),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_204),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_233),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_353),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_234),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_247),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_228),
.B(n_6),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_273),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_283),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_283),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_248),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_283),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_250),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_283),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_257),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_315),
.B(n_8),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_283),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_261),
.B(n_319),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_237),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_314),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_314),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_314),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_314),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_314),
.Y(n_427)
);

BUFx2_ASAP7_75t_SL g428 ( 
.A(n_211),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_261),
.B(n_9),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_260),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_201),
.B(n_9),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_191),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_191),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_194),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_211),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_263),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_267),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_288),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_249),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_278),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_284),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_285),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_201),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_218),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_290),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_218),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_292),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_272),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_229),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_303),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_304),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_190),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_305),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_288),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_249),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_252),
.Y(n_456)
);

CKINVDCx11_ASAP7_75t_R g457 ( 
.A(n_368),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_395),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_404),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_387),
.B(n_184),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_404),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_393),
.B(n_237),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_452),
.B(n_300),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

INVxp33_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

CKINVDCx8_ASAP7_75t_R g468 ( 
.A(n_369),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_404),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_365),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_365),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_389),
.B(n_264),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_421),
.B(n_184),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_403),
.B(n_264),
.Y(n_481)
);

CKINVDCx8_ASAP7_75t_R g482 ( 
.A(n_369),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_367),
.B(n_207),
.Y(n_484)
);

CKINVDCx8_ASAP7_75t_R g485 ( 
.A(n_422),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_410),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_370),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_370),
.Y(n_489)
);

INVx6_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_374),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_435),
.B(n_327),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_412),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_412),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_439),
.B(n_192),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_413),
.B(n_327),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_413),
.B(n_319),
.Y(n_497)
);

BUFx12f_ASAP7_75t_L g498 ( 
.A(n_378),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_455),
.B(n_192),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_415),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_374),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_380),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_417),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_420),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_377),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_377),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_390),
.B(n_195),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_379),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_425),
.B(n_195),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_366),
.A2(n_189),
.B1(n_236),
.B2(n_329),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_379),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_456),
.B(n_252),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_425),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_375),
.A2(n_270),
.B1(n_341),
.B2(n_354),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_426),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_426),
.B(n_357),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_386),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_386),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_388),
.B(n_342),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_388),
.B(n_342),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_391),
.B(n_362),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_443),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_443),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_475),
.B(n_422),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_481),
.B(n_444),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_531),
.A2(n_396),
.B1(n_391),
.B2(n_409),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_528),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_533),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_470),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_528),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_477),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_475),
.B(n_385),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_515),
.B(n_204),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_481),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_533),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_533),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_502),
.B(n_432),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_477),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_484),
.B(n_382),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_477),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_465),
.B(n_392),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_488),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_460),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_488),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_488),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_533),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_531),
.A2(n_396),
.B1(n_429),
.B2(n_371),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_533),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_531),
.B(n_400),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_491),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_531),
.B(n_362),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_515),
.B(n_372),
.C(n_401),
.Y(n_568)
);

AND3x2_ASAP7_75t_L g569 ( 
.A(n_465),
.B(n_272),
.C(n_411),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_533),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_495),
.B(n_405),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_502),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_491),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_480),
.B(n_407),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_460),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

AO21x2_ASAP7_75t_L g578 ( 
.A1(n_495),
.A2(n_500),
.B(n_517),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_500),
.B(n_414),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_479),
.A2(n_419),
.B1(n_431),
.B2(n_381),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_481),
.B(n_444),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_480),
.B(n_416),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_492),
.B(n_430),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_479),
.A2(n_419),
.B1(n_431),
.B2(n_381),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_520),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_474),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_481),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_461),
.B(n_436),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

INVxp33_ASAP7_75t_SL g594 ( 
.A(n_518),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_461),
.B(n_437),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_479),
.A2(n_357),
.B1(n_397),
.B2(n_428),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_514),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_472),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_520),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_460),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_467),
.B(n_440),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_472),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_514),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_516),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_492),
.B(n_441),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_460),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_516),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_516),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_519),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_519),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_496),
.B(n_446),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_464),
.B(n_442),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_492),
.B(n_445),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_519),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_532),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_485),
.B(n_447),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_527),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_527),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_496),
.B(n_450),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_529),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_501),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_476),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_520),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_496),
.B(n_451),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_529),
.A2(n_530),
.B1(n_496),
.B2(n_524),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_529),
.A2(n_428),
.B1(n_287),
.B2(n_251),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_532),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_485),
.B(n_406),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_501),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_476),
.B(n_269),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_478),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_490),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_532),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_524),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_505),
.A2(n_418),
.B1(n_453),
.B2(n_408),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_529),
.A2(n_291),
.B1(n_274),
.B2(n_348),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_490),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_524),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_532),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_478),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_476),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_489),
.Y(n_647)
);

BUFx4f_ASAP7_75t_L g648 ( 
.A(n_530),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_458),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_485),
.B(n_237),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_530),
.A2(n_301),
.B1(n_326),
.B2(n_239),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_457),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_489),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_458),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_459),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_490),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_534),
.B(n_446),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_505),
.B(n_258),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_459),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_466),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_466),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_517),
.B(n_433),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_522),
.A2(n_360),
.B1(n_299),
.B2(n_518),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_468),
.B(n_258),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_530),
.A2(n_244),
.B1(n_262),
.B2(n_266),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_498),
.B(n_490),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_478),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_489),
.B(n_297),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_503),
.B(n_308),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_471),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_471),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_478),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_498),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_503),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_490),
.A2(n_498),
.B1(n_522),
.B2(n_434),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_473),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_497),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_473),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_483),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_478),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_497),
.A2(n_298),
.B1(n_282),
.B2(n_323),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_478),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_468),
.B(n_258),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_503),
.B(n_309),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_503),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_483),
.B(n_312),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_486),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_573),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_649),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_537),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_547),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_592),
.B(n_497),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_588),
.B(n_468),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_586),
.B(n_482),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_595),
.B(n_497),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_537),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_573),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_578),
.B(n_486),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_607),
.B(n_615),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_544),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_537),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_624),
.B(n_482),
.Y(n_703)
);

BUFx4_ASAP7_75t_L g704 ( 
.A(n_652),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_625),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_578),
.B(n_575),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_578),
.B(n_487),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_584),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_585),
.B(n_487),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_674),
.B(n_482),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_R g711 ( 
.A(n_594),
.B(n_373),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_629),
.B(n_494),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_554),
.B(n_494),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_649),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_638),
.B(n_185),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_667),
.B(n_449),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_584),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_584),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_580),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_538),
.B(n_499),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_624),
.B(n_204),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_663),
.A2(n_224),
.B(n_277),
.C(n_279),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_588),
.B(n_383),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_638),
.B(n_186),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_567),
.A2(n_347),
.B1(n_216),
.B2(n_235),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_613),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_565),
.B(n_197),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_613),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_544),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_624),
.B(n_204),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_539),
.B(n_499),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_539),
.B(n_504),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_547),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_648),
.B(n_627),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_654),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_654),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_552),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_655),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_627),
.A2(n_399),
.B1(n_394),
.B2(n_324),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_655),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_601),
.B(n_197),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_552),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_567),
.A2(n_215),
.B1(n_310),
.B2(n_306),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_601),
.B(n_199),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_542),
.B(n_504),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_613),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_542),
.B(n_506),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_659),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_567),
.A2(n_241),
.B1(n_296),
.B2(n_295),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_569),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_621),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_659),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_567),
.A2(n_331),
.B1(n_188),
.B2(n_355),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_678),
.B(n_506),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_678),
.B(n_634),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_571),
.A2(n_313),
.B1(n_321),
.B2(n_325),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_669),
.B(n_507),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_660),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_648),
.A2(n_548),
.B(n_670),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_579),
.A2(n_332),
.B1(n_335),
.B2(n_200),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_628),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_648),
.B(n_204),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_SL g763 ( 
.A(n_650),
.B(n_194),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_660),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_568),
.B(n_199),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_626),
.B(n_507),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_643),
.B(n_200),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_643),
.B(n_509),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_591),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_591),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_623),
.B(n_509),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_661),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_597),
.B(n_202),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_623),
.B(n_510),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_563),
.A2(n_245),
.B1(n_280),
.B2(n_271),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_633),
.Y(n_776)
);

BUFx5_ASAP7_75t_L g777 ( 
.A(n_567),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_625),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_633),
.B(n_510),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_639),
.A2(n_462),
.B(n_463),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_657),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_656),
.B(n_294),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_658),
.B(n_202),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_661),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_671),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_567),
.B(n_288),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_671),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_556),
.B(n_205),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_656),
.B(n_294),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_688),
.B(n_512),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_688),
.B(n_639),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_636),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_646),
.B(n_512),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_625),
.B(n_294),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_646),
.B(n_521),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_625),
.B(n_294),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_657),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_536),
.B(n_449),
.C(n_411),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_647),
.B(n_521),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_647),
.B(n_523),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_672),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_583),
.A2(n_193),
.B(n_351),
.C(n_438),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_625),
.B(n_288),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_653),
.B(n_523),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_653),
.B(n_288),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_636),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_662),
.B(n_675),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_662),
.B(n_525),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_664),
.B(n_219),
.C(n_221),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_603),
.B(n_205),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_587),
.B(n_198),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_567),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_642),
.A2(n_361),
.B1(n_208),
.B2(n_209),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_675),
.B(n_525),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_672),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_686),
.B(n_288),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_686),
.B(n_288),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_546),
.A2(n_289),
.B(n_358),
.C(n_359),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_640),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_642),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_677),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_652),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_580),
.B(n_685),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_679),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_679),
.Y(n_826)
);

CKINVDCx11_ASAP7_75t_R g827 ( 
.A(n_667),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_680),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_614),
.B(n_206),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_630),
.A2(n_687),
.B1(n_641),
.B2(n_651),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_665),
.B(n_286),
.C(n_293),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_680),
.Y(n_832)
);

AO22x2_ASAP7_75t_L g833 ( 
.A1(n_684),
.A2(n_363),
.B1(n_448),
.B2(n_534),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_667),
.B(n_300),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_618),
.B(n_206),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_543),
.Y(n_836)
);

INVxp33_ASAP7_75t_L g837 ( 
.A(n_676),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_619),
.B(n_288),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_546),
.A2(n_462),
.B1(n_463),
.B2(n_469),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_632),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_564),
.B(n_493),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_619),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_594),
.B(n_208),
.Y(n_843)
);

INVx8_ASAP7_75t_L g844 ( 
.A(n_667),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_666),
.B(n_198),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_545),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_564),
.B(n_493),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_543),
.B(n_209),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_564),
.B(n_493),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_545),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_620),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_593),
.B(n_599),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_553),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_553),
.B(n_493),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_555),
.B(n_493),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_545),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_682),
.B(n_300),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_555),
.B(n_557),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_593),
.B(n_535),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_742),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_689),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_699),
.A2(n_559),
.B(n_557),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_706),
.A2(n_589),
.B1(n_559),
.B2(n_560),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_693),
.A2(n_570),
.B(n_576),
.Y(n_864)
);

NAND2x1_ASAP7_75t_L g865 ( 
.A(n_705),
.B(n_856),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_700),
.B(n_560),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_737),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_690),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_700),
.A2(n_598),
.B(n_566),
.C(n_574),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_690),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_696),
.A2(n_570),
.B(n_576),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_755),
.A2(n_570),
.B(n_576),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_824),
.A2(n_582),
.B(n_635),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_R g874 ( 
.A(n_711),
.B(n_210),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_775),
.A2(n_566),
.B(n_574),
.C(n_577),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_577),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_698),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_759),
.A2(n_582),
.B(n_635),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_713),
.B(n_581),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_739),
.B(n_695),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_709),
.B(n_581),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_729),
.B(n_589),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_850),
.A2(n_582),
.B(n_635),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_714),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_712),
.A2(n_600),
.B1(n_596),
.B2(n_598),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_735),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_SL g887 ( 
.A(n_823),
.B(n_210),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_723),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_694),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_734),
.A2(n_551),
.B(n_540),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_734),
.A2(n_551),
.B(n_540),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_705),
.A2(n_551),
.B(n_540),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_810),
.B(n_596),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_810),
.B(n_600),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_707),
.A2(n_551),
.B(n_540),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_711),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_777),
.B(n_545),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_856),
.A2(n_551),
.B(n_540),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_720),
.A2(n_802),
.B(n_722),
.C(n_830),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_780),
.A2(n_605),
.B(n_606),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_695),
.B(n_605),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_719),
.A2(n_561),
.B(n_673),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_735),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_786),
.A2(n_561),
.B(n_673),
.Y(n_904)
);

INVx4_ASAP7_75t_SL g905 ( 
.A(n_812),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_736),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_781),
.A2(n_611),
.B(n_606),
.C(n_609),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_777),
.B(n_545),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_738),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_727),
.B(n_609),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_807),
.A2(n_610),
.B(n_611),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_692),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_757),
.A2(n_561),
.B(n_673),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_727),
.B(n_610),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_740),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_741),
.B(n_535),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_777),
.B(n_558),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_716),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_740),
.Y(n_919)
);

OAI21xp33_ASAP7_75t_L g920 ( 
.A1(n_843),
.A2(n_339),
.B(n_336),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_812),
.B(n_612),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_765),
.A2(n_612),
.B(n_616),
.C(n_337),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_733),
.A2(n_616),
.B1(n_620),
.B2(n_622),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_721),
.A2(n_561),
.B(n_673),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_748),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_751),
.B(n_622),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_761),
.B(n_599),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_730),
.A2(n_561),
.B(n_668),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_797),
.B(n_604),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_716),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_733),
.B(n_604),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_691),
.B(n_645),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_741),
.B(n_448),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_765),
.A2(n_336),
.B(n_337),
.C(n_338),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_776),
.B(n_768),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_837),
.B(n_637),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_744),
.B(n_338),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_777),
.B(n_558),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_792),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_752),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_710),
.B(n_212),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_843),
.B(n_637),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_819),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_840),
.B(n_644),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_744),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_777),
.B(n_558),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_750),
.A2(n_550),
.B(n_541),
.C(n_549),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_730),
.A2(n_668),
.B(n_602),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_752),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_762),
.A2(n_562),
.B(n_590),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_758),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_762),
.A2(n_668),
.B(n_602),
.Y(n_952)
);

O2A1O1Ixp5_ASAP7_75t_L g953 ( 
.A1(n_782),
.A2(n_683),
.B(n_681),
.C(n_645),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_692),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_841),
.A2(n_668),
.B(n_602),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_777),
.B(n_558),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_788),
.A2(n_339),
.B(n_340),
.C(n_341),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_767),
.B(n_644),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_847),
.A2(n_668),
.B(n_602),
.Y(n_959)
);

INVx5_ASAP7_75t_L g960 ( 
.A(n_812),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_758),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_849),
.A2(n_558),
.B(n_602),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_857),
.B(n_340),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_764),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_791),
.A2(n_608),
.B(n_681),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_858),
.A2(n_550),
.B(n_541),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_767),
.B(n_792),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_L g968 ( 
.A(n_835),
.B(n_645),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_806),
.B(n_549),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_692),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_764),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_806),
.B(n_562),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_844),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_821),
.B(n_572),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_772),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_821),
.B(n_715),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_715),
.B(n_572),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_772),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_692),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_846),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_846),
.A2(n_608),
.B(n_683),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_715),
.B(n_590),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_784),
.A2(n_787),
.B(n_785),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_782),
.A2(n_608),
.B(n_683),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_724),
.B(n_608),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_704),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_827),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_811),
.B(n_225),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_724),
.B(n_697),
.Y(n_989)
);

INVx3_ASAP7_75t_SL g990 ( 
.A(n_716),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_784),
.A2(n_617),
.B(n_631),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_724),
.B(n_631),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_702),
.B(n_631),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_708),
.B(n_631),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_812),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_717),
.B(n_631),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_773),
.A2(n_454),
.B(n_463),
.C(n_462),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_718),
.B(n_617),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_777),
.B(n_617),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_783),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_785),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_793),
.A2(n_454),
.B(n_469),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_726),
.B(n_617),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_728),
.B(n_617),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_787),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_835),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_SL g1007 ( 
.A(n_844),
.B(n_213),
.Y(n_1007)
);

AND2x2_ASAP7_75t_SL g1008 ( 
.A(n_788),
.B(n_511),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_763),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_703),
.B(n_226),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_746),
.B(n_214),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_801),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_833),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_801),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_852),
.B(n_275),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_815),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_789),
.A2(n_361),
.B(n_275),
.C(n_511),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_859),
.B(n_511),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_815),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_769),
.B(n_511),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_789),
.A2(n_526),
.B(n_513),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_852),
.B(n_526),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_820),
.A2(n_307),
.B(n_240),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_770),
.B(n_511),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_848),
.B(n_511),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_848),
.B(n_513),
.Y(n_1026)
);

CKINVDCx14_ASAP7_75t_R g1027 ( 
.A(n_834),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_783),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_820),
.Y(n_1029)
);

AO21x1_ASAP7_75t_L g1030 ( 
.A1(n_803),
.A2(n_11),
.B(n_12),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_822),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_825),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_703),
.A2(n_817),
.B(n_816),
.C(n_805),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_852),
.B(n_513),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_798),
.B(n_344),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_766),
.B(n_513),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_822),
.B(n_826),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_826),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_828),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_828),
.B(n_513),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_754),
.A2(n_526),
.B(n_302),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_829),
.A2(n_526),
.B1(n_311),
.B2(n_281),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_829),
.B(n_344),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_832),
.B(n_731),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_845),
.B(n_345),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_864),
.A2(n_778),
.B(n_743),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_880),
.A2(n_831),
.B1(n_833),
.B2(n_756),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_870),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_937),
.B(n_809),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_945),
.B(n_813),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_903),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_973),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_871),
.A2(n_778),
.B(n_725),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_1006),
.A2(n_833),
.B1(n_753),
.B2(n_749),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_988),
.A2(n_760),
.B(n_346),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_877),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_957),
.A2(n_732),
.B(n_745),
.C(n_747),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_866),
.A2(n_855),
.B(n_854),
.Y(n_1058)
);

O2A1O1Ixp5_ASAP7_75t_L g1059 ( 
.A1(n_901),
.A2(n_790),
.B(n_803),
.C(n_796),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_967),
.A2(n_774),
.B(n_771),
.Y(n_1060)
);

BUFx12f_ASAP7_75t_L g1061 ( 
.A(n_987),
.Y(n_1061)
);

CKINVDCx8_ASAP7_75t_R g1062 ( 
.A(n_896),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_903),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1000),
.B(n_844),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_897),
.A2(n_779),
.B(n_794),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1028),
.B(n_832),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_957),
.A2(n_805),
.B(n_816),
.C(n_817),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_943),
.B(n_836),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_860),
.B(n_853),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_889),
.B(n_795),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_886),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_897),
.A2(n_794),
.B(n_796),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_861),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_874),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_889),
.A2(n_799),
.B1(n_804),
.B2(n_808),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1008),
.A2(n_800),
.B1(n_814),
.B2(n_851),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_919),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_867),
.B(n_842),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_SL g1079 ( 
.A1(n_1027),
.A2(n_345),
.B1(n_346),
.B2(n_349),
.Y(n_1079)
);

CKINVDCx10_ASAP7_75t_R g1080 ( 
.A(n_986),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_934),
.A2(n_818),
.B(n_838),
.C(n_842),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_888),
.B(n_851),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_934),
.B(n_354),
.C(n_352),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_908),
.A2(n_838),
.B(n_839),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_958),
.A2(n_526),
.B(n_268),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_908),
.A2(n_526),
.B(n_109),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_940),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_901),
.B(n_352),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_1027),
.B(n_350),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_942),
.B(n_350),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_942),
.B(n_349),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_988),
.A2(n_920),
.B1(n_1043),
.B2(n_1010),
.C(n_963),
.Y(n_1092)
);

AOI21xp33_ASAP7_75t_L g1093 ( 
.A1(n_1010),
.A2(n_899),
.B(n_936),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_916),
.B(n_328),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_861),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_976),
.B(n_322),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_936),
.B(n_318),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_949),
.Y(n_1098)
);

AND2x2_ASAP7_75t_SL g1099 ( 
.A(n_973),
.B(n_14),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_874),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_909),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_995),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_964),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_862),
.A2(n_950),
.B(n_1025),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_995),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_995),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_909),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_917),
.A2(n_87),
.B(n_172),
.Y(n_1108)
);

AOI33xp33_ASAP7_75t_L g1109 ( 
.A1(n_1035),
.A2(n_276),
.A3(n_265),
.B1(n_259),
.B2(n_256),
.B3(n_255),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1008),
.A2(n_253),
.B1(n_246),
.B2(n_243),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_1045),
.B(n_933),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1013),
.A2(n_238),
.B1(n_20),
.B2(n_27),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_876),
.B(n_18),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_917),
.A2(n_63),
.B(n_169),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_876),
.B(n_18),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_989),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1015),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_941),
.B(n_1007),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_922),
.A2(n_34),
.B(n_38),
.C(n_40),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_935),
.B(n_887),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_995),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_879),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1015),
.A2(n_932),
.B1(n_1009),
.B2(n_1011),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_971),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_912),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_918),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_938),
.A2(n_93),
.B(n_163),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_915),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_921),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_930),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_882),
.B(n_85),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1033),
.A2(n_44),
.B(n_46),
.C(n_47),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1005),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_912),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1032),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_960),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_922),
.A2(n_48),
.B(n_49),
.C(n_51),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_915),
.Y(n_1138)
);

OAI21xp33_ASAP7_75t_L g1139 ( 
.A1(n_1023),
.A2(n_882),
.B(n_1042),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_SL g1140 ( 
.A1(n_990),
.A2(n_954),
.B1(n_1032),
.B2(n_944),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_926),
.A2(n_48),
.B(n_51),
.C(n_52),
.Y(n_1141)
);

BUFx4f_ASAP7_75t_L g1142 ( 
.A(n_990),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_881),
.B(n_122),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_938),
.A2(n_116),
.B(n_162),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_939),
.B(n_53),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1016),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1018),
.A2(n_110),
.B(n_159),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_869),
.A2(n_107),
.B(n_158),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_927),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_960),
.B(n_81),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_960),
.B(n_139),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1031),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_932),
.A2(n_78),
.B1(n_156),
.B2(n_151),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_SL g1154 ( 
.A(n_944),
.B(n_53),
.C(n_55),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1038),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_970),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_929),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_893),
.B(n_75),
.Y(n_1158)
);

NAND2x2_ASAP7_75t_L g1159 ( 
.A(n_910),
.B(n_59),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_946),
.A2(n_150),
.B(n_171),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_894),
.B(n_1044),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_914),
.A2(n_968),
.B(n_907),
.C(n_875),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_946),
.A2(n_956),
.B(n_873),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1039),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_977),
.A2(n_982),
.B(n_869),
.C(n_1017),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_954),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_947),
.A2(n_1030),
.B(n_885),
.C(n_923),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_985),
.A2(n_1026),
.B(n_911),
.C(n_1041),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_951),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_970),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_960),
.B(n_998),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_951),
.A2(n_975),
.B1(n_961),
.B2(n_1019),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_961),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_997),
.A2(n_872),
.B(n_1001),
.C(n_868),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_979),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_956),
.A2(n_878),
.B(n_883),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_992),
.A2(n_999),
.B(n_1036),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_975),
.Y(n_1178)
);

BUFx2_ASAP7_75t_SL g1179 ( 
.A(n_979),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_863),
.A2(n_972),
.B(n_974),
.C(n_969),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1014),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1037),
.A2(n_1020),
.B(n_1024),
.C(n_1012),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_900),
.A2(n_965),
.B(n_931),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_980),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_980),
.Y(n_1185)
);

OAI21xp33_ASAP7_75t_SL g1186 ( 
.A1(n_983),
.A2(n_991),
.B(n_1034),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1019),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_998),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_921),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_999),
.A2(n_865),
.B(n_895),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_884),
.A2(n_925),
.B1(n_1029),
.B2(n_978),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_962),
.A2(n_959),
.B(n_955),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_906),
.Y(n_1193)
);

OR2x6_ASAP7_75t_SL g1194 ( 
.A(n_993),
.B(n_996),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_905),
.Y(n_1195)
);

NOR2x1p5_ASAP7_75t_L g1196 ( 
.A(n_994),
.B(n_1004),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_905),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1022),
.A2(n_902),
.B(n_981),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_966),
.A2(n_904),
.B(n_913),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1040),
.Y(n_1200)
);

AO22x1_ASAP7_75t_L g1201 ( 
.A1(n_921),
.A2(n_1003),
.B1(n_905),
.B2(n_953),
.Y(n_1201)
);

OA22x2_ASAP7_75t_L g1202 ( 
.A1(n_1002),
.A2(n_921),
.B1(n_984),
.B2(n_948),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_952),
.A2(n_924),
.B(n_928),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_890),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1197),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1126),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1094),
.B(n_1021),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1168),
.A2(n_891),
.A3(n_892),
.B(n_898),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1093),
.A2(n_1199),
.B(n_1183),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1093),
.A2(n_1139),
.B(n_1162),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1092),
.A2(n_1055),
.B(n_1113),
.C(n_1115),
.Y(n_1211)
);

AO32x2_ASAP7_75t_L g1212 ( 
.A1(n_1122),
.A2(n_1112),
.A3(n_1140),
.B1(n_1054),
.B2(n_1076),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1176),
.A2(n_1190),
.B(n_1192),
.Y(n_1213)
);

O2A1O1Ixp5_ASAP7_75t_L g1214 ( 
.A1(n_1118),
.A2(n_1120),
.B(n_1088),
.C(n_1131),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1165),
.A2(n_1183),
.A3(n_1174),
.B(n_1076),
.Y(n_1215)
);

OAI22x1_ASAP7_75t_L g1216 ( 
.A1(n_1047),
.A2(n_1145),
.B1(n_1123),
.B2(n_1049),
.Y(n_1216)
);

AO21x1_ASAP7_75t_L g1217 ( 
.A1(n_1158),
.A2(n_1167),
.B(n_1137),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1203),
.A2(n_1202),
.B(n_1163),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1056),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1092),
.A2(n_1100),
.B1(n_1050),
.B2(n_1068),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1057),
.A2(n_1088),
.B(n_1161),
.C(n_1158),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1059),
.A2(n_1186),
.B(n_1161),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1169),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1046),
.A2(n_1053),
.B(n_1060),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1111),
.A2(n_1157),
.B1(n_1070),
.B2(n_1091),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1132),
.A2(n_1177),
.A3(n_1172),
.B(n_1198),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1069),
.B(n_1095),
.Y(n_1227)
);

NAND3xp33_ASAP7_75t_L g1228 ( 
.A(n_1083),
.B(n_1154),
.C(n_1117),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1090),
.A2(n_1091),
.B(n_1112),
.C(n_1122),
.Y(n_1229)
);

OR2x6_ASAP7_75t_L g1230 ( 
.A(n_1052),
.B(n_1195),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1150),
.A2(n_1151),
.B(n_1143),
.C(n_1054),
.Y(n_1231)
);

O2A1O1Ixp5_ASAP7_75t_SL g1232 ( 
.A1(n_1204),
.A2(n_1097),
.B(n_1096),
.C(n_1110),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1090),
.B(n_1073),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1109),
.B(n_1116),
.C(n_1110),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1060),
.A2(n_1058),
.B(n_1180),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1051),
.Y(n_1236)
);

NAND3x1_ASAP7_75t_L g1237 ( 
.A(n_1064),
.B(n_1078),
.C(n_1066),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1135),
.B(n_1149),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1067),
.A2(n_1081),
.B(n_1143),
.C(n_1119),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1075),
.B(n_1200),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1052),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_1130),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1104),
.A2(n_1204),
.B(n_1072),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1061),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1172),
.A2(n_1085),
.A3(n_1065),
.B(n_1084),
.Y(n_1245)
);

O2A1O1Ixp5_ASAP7_75t_L g1246 ( 
.A1(n_1201),
.A2(n_1085),
.B(n_1086),
.C(n_1147),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1129),
.A2(n_1136),
.B(n_1182),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1188),
.B(n_1185),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1129),
.A2(n_1136),
.B(n_1171),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1141),
.A2(n_1082),
.B(n_1152),
.C(n_1071),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1173),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1178),
.A2(n_1181),
.A3(n_1146),
.B(n_1155),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1129),
.A2(n_1194),
.B1(n_1164),
.B2(n_1133),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1129),
.A2(n_1103),
.B1(n_1124),
.B2(n_1087),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1189),
.A2(n_1196),
.B(n_1063),
.Y(n_1255)
);

NAND3x1_ASAP7_75t_L g1256 ( 
.A(n_1153),
.B(n_1099),
.C(n_1080),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1077),
.B(n_1098),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1074),
.A2(n_1079),
.B1(n_1159),
.B2(n_1142),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1191),
.A2(n_1193),
.B(n_1127),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1108),
.A2(n_1160),
.B(n_1144),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1101),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1114),
.A2(n_1184),
.B(n_1187),
.C(n_1128),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1107),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1138),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1166),
.A2(n_1148),
.B(n_1184),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1142),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1195),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1148),
.A2(n_1106),
.B(n_1102),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1102),
.A2(n_1105),
.B(n_1106),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1156),
.B(n_1170),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1105),
.A2(n_1121),
.B(n_1125),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_SL g1272 ( 
.A1(n_1179),
.A2(n_1125),
.B(n_1134),
.C(n_1175),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1089),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1125),
.A2(n_1134),
.B(n_1062),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1134),
.A2(n_1092),
.B(n_1139),
.C(n_1055),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1168),
.A2(n_869),
.A3(n_1162),
.B(n_1165),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1048),
.Y(n_1278)
);

AO32x2_ASAP7_75t_L g1279 ( 
.A1(n_1122),
.A2(n_1013),
.A3(n_1112),
.B1(n_775),
.B2(n_1140),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1169),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1061),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1111),
.B(n_1006),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1169),
.Y(n_1284)
);

AO32x2_ASAP7_75t_L g1285 ( 
.A1(n_1122),
.A2(n_1013),
.A3(n_1112),
.B1(n_775),
.B2(n_1140),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1183),
.A2(n_1168),
.B(n_869),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1169),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1094),
.B(n_937),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1168),
.A2(n_869),
.A3(n_1162),
.B(n_1165),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1094),
.B(n_937),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1197),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1168),
.A2(n_869),
.A3(n_1162),
.B(n_1165),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1088),
.B(n_700),
.Y(n_1295)
);

OAI22x1_ASAP7_75t_L g1296 ( 
.A1(n_1113),
.A2(n_1006),
.B1(n_1115),
.B2(n_1047),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1168),
.A2(n_869),
.A3(n_1162),
.B(n_1165),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1093),
.A2(n_1139),
.B(n_700),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1056),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1051),
.Y(n_1300)
);

AOI221x1_ASAP7_75t_L g1301 ( 
.A1(n_1093),
.A2(n_1139),
.B1(n_1132),
.B2(n_1113),
.C(n_1115),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1168),
.A2(n_869),
.A3(n_1162),
.B(n_1165),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1113),
.A2(n_1115),
.B(n_1000),
.C(n_1028),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1197),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1122),
.A2(n_1013),
.A3(n_1112),
.B1(n_775),
.B2(n_1140),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1183),
.A2(n_1168),
.B(n_869),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1093),
.A2(n_1139),
.B(n_700),
.Y(n_1309)
);

AO32x2_ASAP7_75t_L g1310 ( 
.A1(n_1122),
.A2(n_1013),
.A3(n_1112),
.B1(n_775),
.B2(n_1140),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1176),
.A2(n_1002),
.B(n_1190),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1168),
.A2(n_869),
.A3(n_1162),
.B(n_1165),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1094),
.B(n_937),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1052),
.B(n_1188),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1111),
.B(n_742),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1088),
.B(n_700),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1126),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1176),
.A2(n_1002),
.B(n_1190),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1093),
.A2(n_1139),
.B(n_700),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1126),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1176),
.A2(n_1002),
.B(n_1190),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1162),
.A2(n_1161),
.B(n_1168),
.Y(n_1323)
);

AOI221xp5_ASAP7_75t_L g1324 ( 
.A1(n_1092),
.A2(n_664),
.B1(n_988),
.B2(n_843),
.C(n_1006),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1176),
.A2(n_1002),
.B(n_1190),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1176),
.A2(n_1002),
.B(n_1190),
.Y(n_1326)
);

NAND2x1p5_ASAP7_75t_L g1327 ( 
.A(n_1195),
.B(n_1129),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1048),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1055),
.A2(n_957),
.B1(n_934),
.B2(n_664),
.C(n_1113),
.Y(n_1329)
);

O2A1O1Ixp5_ASAP7_75t_SL g1330 ( 
.A1(n_1093),
.A2(n_1122),
.B(n_775),
.C(n_1204),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1088),
.B(n_700),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1093),
.A2(n_1199),
.B(n_1183),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1052),
.B(n_1188),
.Y(n_1333)
);

INVx3_ASAP7_75t_SL g1334 ( 
.A(n_1074),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1169),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1092),
.A2(n_1006),
.B1(n_711),
.B2(n_373),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1092),
.A2(n_1139),
.B(n_1055),
.C(n_1093),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1113),
.A2(n_1115),
.B(n_1000),
.C(n_1028),
.Y(n_1339)
);

NOR2xp67_ASAP7_75t_L g1340 ( 
.A(n_1111),
.B(n_751),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1341)
);

AOI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1092),
.A2(n_664),
.B1(n_988),
.B2(n_843),
.C(n_1006),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1113),
.A2(n_1115),
.B(n_1000),
.C(n_1028),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1093),
.A2(n_1139),
.B(n_700),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1161),
.A2(n_1006),
.B1(n_945),
.B2(n_1092),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1093),
.A2(n_1139),
.B(n_700),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1093),
.A2(n_1199),
.B(n_1183),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1073),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1176),
.A2(n_1002),
.B(n_1190),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_SL g1351 ( 
.A(n_1129),
.B(n_485),
.Y(n_1351)
);

INVx8_ASAP7_75t_L g1352 ( 
.A(n_1052),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1094),
.B(n_937),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1048),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1183),
.A2(n_1168),
.B(n_869),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1088),
.B(n_700),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1111),
.B(n_751),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1051),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1051),
.Y(n_1359)
);

AOI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1104),
.A2(n_862),
.B(n_1163),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1055),
.A2(n_1092),
.B1(n_843),
.B2(n_810),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1168),
.A2(n_1176),
.B(n_648),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1073),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_SL g1364 ( 
.A(n_1062),
.B(n_823),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1257),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1219),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1244),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1361),
.A2(n_1342),
.B1(n_1324),
.B2(n_1211),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1334),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1282),
.Y(n_1370)
);

BUFx4f_ASAP7_75t_L g1371 ( 
.A(n_1352),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1273),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1267),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1336),
.A2(n_1220),
.B1(n_1283),
.B2(n_1237),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1295),
.B(n_1316),
.Y(n_1375)
);

INVx6_ASAP7_75t_L g1376 ( 
.A(n_1241),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1206),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1331),
.B(n_1356),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1278),
.Y(n_1379)
);

BUFx2_ASAP7_75t_SL g1380 ( 
.A(n_1241),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1296),
.A2(n_1216),
.B1(n_1228),
.B2(n_1234),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1345),
.A2(n_1210),
.B1(n_1298),
.B2(n_1346),
.Y(n_1382)
);

INVx6_ASAP7_75t_L g1383 ( 
.A(n_1352),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1328),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1299),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1267),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1354),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1317),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1315),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1261),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1309),
.A2(n_1344),
.B1(n_1320),
.B2(n_1225),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1364),
.A2(n_1222),
.B1(n_1353),
.B2(n_1291),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1263),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1264),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1351),
.B(n_1255),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1321),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1288),
.A2(n_1313),
.B1(n_1217),
.B2(n_1207),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1223),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1240),
.A2(n_1233),
.B1(n_1227),
.B2(n_1209),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1276),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1223),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1251),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1256),
.A2(n_1357),
.B1(n_1340),
.B2(n_1329),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1242),
.Y(n_1404)
);

BUFx10_ASAP7_75t_L g1405 ( 
.A(n_1205),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1258),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1280),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1301),
.A2(n_1238),
.B1(n_1349),
.B2(n_1363),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1303),
.A2(n_1343),
.B(n_1339),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1253),
.A2(n_1259),
.B1(n_1332),
.B2(n_1348),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1254),
.A2(n_1266),
.B1(n_1358),
.B2(n_1359),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1300),
.A2(n_1280),
.B1(n_1284),
.B2(n_1335),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1230),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1284),
.A2(n_1335),
.B1(n_1287),
.B2(n_1333),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1314),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1205),
.A2(n_1292),
.B1(n_1304),
.B2(n_1212),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1230),
.Y(n_1417)
);

BUFx10_ASAP7_75t_L g1418 ( 
.A(n_1205),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1286),
.A2(n_1308),
.B1(n_1355),
.B2(n_1235),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1287),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1252),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1252),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1292),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1286),
.A2(n_1355),
.B1(n_1308),
.B2(n_1224),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1337),
.A2(n_1275),
.B1(n_1239),
.B2(n_1221),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1229),
.A2(n_1212),
.B1(n_1292),
.B2(n_1304),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1212),
.A2(n_1304),
.B1(n_1260),
.B2(n_1285),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1323),
.A2(n_1310),
.B1(n_1306),
.B2(n_1285),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1248),
.A2(n_1270),
.B1(n_1310),
.B2(n_1306),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1314),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1333),
.A2(n_1250),
.B1(n_1327),
.B2(n_1262),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1272),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1279),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1231),
.B(n_1312),
.Y(n_1434)
);

BUFx4f_ASAP7_75t_SL g1435 ( 
.A(n_1274),
.Y(n_1435)
);

INVx5_ASAP7_75t_L g1436 ( 
.A(n_1246),
.Y(n_1436)
);

BUFx4f_ASAP7_75t_L g1437 ( 
.A(n_1214),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1279),
.A2(n_1310),
.B1(n_1306),
.B2(n_1285),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1290),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1290),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1232),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_1271),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1247),
.A2(n_1249),
.B1(n_1265),
.B2(n_1362),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1277),
.A2(n_1347),
.B1(n_1319),
.B2(n_1341),
.Y(n_1444)
);

INVxp67_ASAP7_75t_SL g1445 ( 
.A(n_1218),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1294),
.Y(n_1446)
);

BUFx8_ASAP7_75t_SL g1447 ( 
.A(n_1360),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1269),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1294),
.Y(n_1449)
);

OAI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1281),
.A2(n_1307),
.B1(n_1338),
.B2(n_1305),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1297),
.Y(n_1451)
);

CKINVDCx6p67_ASAP7_75t_R g1452 ( 
.A(n_1330),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1289),
.A2(n_1293),
.B1(n_1302),
.B2(n_1297),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1268),
.A2(n_1243),
.B1(n_1213),
.B2(n_1312),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_1297),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1245),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1245),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1302),
.B(n_1312),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1226),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1245),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1350),
.A2(n_1318),
.B1(n_1325),
.B2(n_1322),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_SL g1462 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_1208),
.B2(n_1311),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1326),
.B(n_1215),
.Y(n_1463)
);

BUFx4_ASAP7_75t_SL g1464 ( 
.A(n_1226),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1208),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1215),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1295),
.B(n_1316),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1336),
.A2(n_1006),
.B1(n_1342),
.B2(n_1324),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1219),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1324),
.B(n_1006),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1211),
.A2(n_1361),
.B(n_810),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1324),
.A2(n_1342),
.B1(n_1296),
.B2(n_1361),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1241),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1257),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1288),
.B(n_1291),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1276),
.Y(n_1476)
);

INVx6_ASAP7_75t_L g1477 ( 
.A(n_1241),
.Y(n_1477)
);

BUFx10_ASAP7_75t_L g1478 ( 
.A(n_1205),
.Y(n_1478)
);

INVx6_ASAP7_75t_L g1479 ( 
.A(n_1241),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1244),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1324),
.A2(n_1342),
.B1(n_1006),
.B2(n_1296),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1351),
.B(n_1129),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1236),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1257),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1345),
.A2(n_465),
.B1(n_475),
.B2(n_1099),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1257),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1219),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1244),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1257),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1295),
.B(n_1316),
.Y(n_1490)
);

CKINVDCx11_ASAP7_75t_R g1491 ( 
.A(n_1244),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1257),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1324),
.A2(n_1342),
.B1(n_1296),
.B2(n_1361),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1324),
.A2(n_1342),
.B1(n_1296),
.B2(n_1361),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1295),
.B(n_1316),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1236),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1257),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1324),
.A2(n_1342),
.B1(n_1361),
.B2(n_1296),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1447),
.Y(n_1499)
);

BUFx4f_ASAP7_75t_SL g1500 ( 
.A(n_1488),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1465),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1457),
.B(n_1466),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1421),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1481),
.A2(n_1368),
.B1(n_1374),
.B2(n_1468),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1422),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1458),
.B(n_1439),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1400),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1400),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1470),
.B(n_1475),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1365),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1476),
.B(n_1427),
.Y(n_1511)
);

BUFx4f_ASAP7_75t_SL g1512 ( 
.A(n_1369),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1476),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1461),
.A2(n_1443),
.B(n_1454),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1389),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1440),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1433),
.B(n_1455),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1377),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1446),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1449),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1451),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1461),
.A2(n_1454),
.B(n_1444),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1459),
.Y(n_1523)
);

CKINVDCx16_ASAP7_75t_R g1524 ( 
.A(n_1480),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1458),
.B(n_1428),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1398),
.Y(n_1526)
);

AOI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1463),
.A2(n_1425),
.B(n_1431),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1388),
.B(n_1404),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1401),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1456),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1375),
.B(n_1378),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1428),
.B(n_1438),
.Y(n_1532)
);

AOI211xp5_ASAP7_75t_L g1533 ( 
.A1(n_1468),
.A2(n_1409),
.B(n_1471),
.C(n_1408),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1467),
.B(n_1490),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1402),
.Y(n_1535)
);

BUFx2_ASAP7_75t_SL g1536 ( 
.A(n_1448),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1407),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1420),
.Y(n_1538)
);

AO21x2_ASAP7_75t_L g1539 ( 
.A1(n_1450),
.A2(n_1434),
.B(n_1445),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1436),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1395),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1464),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1396),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1438),
.B(n_1416),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1424),
.A2(n_1419),
.B(n_1395),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1464),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1437),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1474),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1436),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1416),
.B(n_1391),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1436),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1385),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1419),
.A2(n_1424),
.B(n_1410),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1445),
.A2(n_1482),
.B(n_1412),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1498),
.A2(n_1472),
.B1(n_1493),
.B2(n_1494),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1436),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1379),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1384),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1498),
.A2(n_1391),
.B(n_1382),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1495),
.B(n_1484),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1387),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1390),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1393),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1394),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1372),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1462),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1485),
.A2(n_1381),
.B1(n_1403),
.B2(n_1426),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1397),
.A2(n_1399),
.B(n_1426),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1482),
.A2(n_1432),
.B(n_1414),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1460),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1452),
.Y(n_1571)
);

AO21x2_ASAP7_75t_L g1572 ( 
.A1(n_1450),
.A2(n_1429),
.B(n_1408),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1429),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1417),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1437),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1453),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1453),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1382),
.B(n_1399),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1483),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1485),
.A2(n_1392),
.B(n_1411),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1486),
.B(n_1497),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1496),
.Y(n_1582)
);

OAI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1406),
.A2(n_1435),
.B1(n_1417),
.B2(n_1492),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1441),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1489),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1442),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1373),
.A2(n_1442),
.B(n_1392),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1413),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1435),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1415),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1430),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1430),
.A2(n_1386),
.B(n_1380),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1376),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1386),
.B(n_1477),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1371),
.A2(n_1366),
.B(n_1469),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1376),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1376),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1473),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1473),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1473),
.A2(n_1477),
.B(n_1479),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1477),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1515),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1555),
.A2(n_1371),
.B1(n_1479),
.B2(n_1383),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1527),
.B(n_1383),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1510),
.B(n_1487),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1517),
.B(n_1405),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_SL g1607 ( 
.A(n_1547),
.B(n_1491),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1533),
.A2(n_1479),
.B1(n_1383),
.B2(n_1423),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1548),
.B(n_1405),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1501),
.B(n_1367),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1517),
.B(n_1418),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1526),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1529),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1570),
.B(n_1418),
.Y(n_1614)
);

INVx11_ASAP7_75t_L g1615 ( 
.A(n_1512),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1559),
.A2(n_1370),
.B(n_1478),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1535),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1524),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1514),
.A2(n_1522),
.B(n_1566),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1501),
.B(n_1506),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1531),
.B(n_1534),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1504),
.A2(n_1567),
.B1(n_1533),
.B2(n_1580),
.C(n_1578),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_SL g1623 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1578),
.A2(n_1550),
.B1(n_1576),
.B2(n_1577),
.C(n_1509),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1502),
.B(n_1511),
.Y(n_1625)
);

NOR2xp67_ASAP7_75t_SL g1626 ( 
.A(n_1499),
.B(n_1589),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1560),
.B(n_1581),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1585),
.B(n_1518),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1550),
.A2(n_1576),
.B(n_1577),
.C(n_1587),
.Y(n_1629)
);

OAI21x1_ASAP7_75t_L g1630 ( 
.A1(n_1522),
.A2(n_1545),
.B(n_1587),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1535),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1499),
.A2(n_1586),
.B(n_1547),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1518),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1573),
.A2(n_1584),
.B1(n_1572),
.B2(n_1544),
.C(n_1566),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1525),
.B(n_1542),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1572),
.A2(n_1539),
.B(n_1553),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1536),
.A2(n_1583),
.B1(n_1575),
.B2(n_1547),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1572),
.A2(n_1539),
.B(n_1553),
.Y(n_1638)
);

AOI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1573),
.A2(n_1584),
.B1(n_1572),
.B2(n_1544),
.C(n_1532),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1584),
.A2(n_1571),
.B(n_1499),
.C(n_1590),
.Y(n_1640)
);

OA21x2_ASAP7_75t_L g1641 ( 
.A1(n_1545),
.A2(n_1551),
.B(n_1549),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1525),
.B(n_1542),
.Y(n_1642)
);

AO32x2_ASAP7_75t_L g1643 ( 
.A1(n_1532),
.A2(n_1502),
.A3(n_1511),
.B1(n_1513),
.B2(n_1508),
.Y(n_1643)
);

AO21x2_ASAP7_75t_L g1644 ( 
.A1(n_1540),
.A2(n_1556),
.B(n_1551),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1575),
.A2(n_1547),
.B(n_1589),
.C(n_1571),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1541),
.B(n_1600),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1546),
.B(n_1530),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1589),
.A2(n_1571),
.B(n_1569),
.C(n_1554),
.Y(n_1648)
);

A2O1A1Ixp33_ASAP7_75t_L g1649 ( 
.A1(n_1589),
.A2(n_1569),
.B(n_1554),
.C(n_1600),
.Y(n_1649)
);

AO32x2_ASAP7_75t_L g1650 ( 
.A1(n_1507),
.A2(n_1513),
.A3(n_1508),
.B1(n_1503),
.B2(n_1505),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1562),
.B(n_1563),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1552),
.A2(n_1595),
.B(n_1592),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1574),
.A2(n_1568),
.B(n_1599),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1523),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1568),
.A2(n_1553),
.B1(n_1574),
.B2(n_1539),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1538),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1564),
.B(n_1537),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1538),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1591),
.B(n_1568),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1557),
.Y(n_1660)
);

AND4x1_ASAP7_75t_L g1661 ( 
.A(n_1622),
.B(n_1528),
.C(n_1601),
.D(n_1599),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1539),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1654),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1650),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1609),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1619),
.B(n_1553),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1619),
.B(n_1523),
.Y(n_1667)
);

NOR2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1618),
.B(n_1588),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1616),
.A2(n_1543),
.B1(n_1565),
.B2(n_1561),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1643),
.B(n_1659),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1659),
.B(n_1520),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1646),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1641),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1624),
.A2(n_1557),
.B1(n_1558),
.B2(n_1579),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1643),
.B(n_1521),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1643),
.B(n_1521),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1621),
.B(n_1652),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1643),
.B(n_1521),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1650),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1641),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1655),
.B(n_1519),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1630),
.B(n_1519),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1650),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1640),
.B(n_1588),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1639),
.A2(n_1579),
.B1(n_1582),
.B2(n_1591),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1634),
.B(n_1541),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1644),
.B(n_1516),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1629),
.A2(n_1588),
.B1(n_1598),
.B2(n_1597),
.Y(n_1689)
);

INVx4_ASAP7_75t_L g1690 ( 
.A(n_1604),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1670),
.B(n_1636),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1670),
.B(n_1638),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1670),
.B(n_1635),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1677),
.A2(n_1602),
.B1(n_1608),
.B2(n_1637),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1677),
.A2(n_1611),
.B1(n_1606),
.B2(n_1618),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1662),
.B(n_1664),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_SL g1697 ( 
.A(n_1661),
.B(n_1640),
.C(n_1629),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1667),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1642),
.Y(n_1699)
);

NAND4xp25_ASAP7_75t_L g1700 ( 
.A(n_1686),
.B(n_1623),
.C(n_1605),
.D(n_1653),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1662),
.B(n_1664),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1663),
.Y(n_1702)
);

AO21x2_ASAP7_75t_L g1703 ( 
.A1(n_1666),
.A2(n_1648),
.B(n_1649),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1690),
.Y(n_1704)
);

AO21x2_ASAP7_75t_L g1705 ( 
.A1(n_1666),
.A2(n_1648),
.B(n_1649),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1663),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1688),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1686),
.A2(n_1603),
.B1(n_1610),
.B2(n_1614),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1679),
.B(n_1651),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1671),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1688),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1679),
.B(n_1657),
.Y(n_1712)
);

OAI33xp33_ASAP7_75t_L g1713 ( 
.A1(n_1687),
.A2(n_1628),
.A3(n_1633),
.B1(n_1627),
.B2(n_1660),
.B3(n_1656),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1688),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1672),
.Y(n_1715)
);

AOI33xp33_ASAP7_75t_L g1716 ( 
.A1(n_1674),
.A2(n_1647),
.A3(n_1617),
.B1(n_1658),
.B2(n_1631),
.B3(n_1612),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1680),
.B(n_1613),
.Y(n_1717)
);

NAND2x1_ASAP7_75t_SL g1718 ( 
.A(n_1682),
.B(n_1620),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1681),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1694),
.B(n_1661),
.C(n_1674),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1719),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1702),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_SL g1723 ( 
.A1(n_1697),
.A2(n_1689),
.B1(n_1607),
.B2(n_1682),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1717),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1691),
.B(n_1676),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1717),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1717),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1691),
.B(n_1676),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1706),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1698),
.Y(n_1731)
);

NOR4xp25_ASAP7_75t_SL g1732 ( 
.A(n_1697),
.B(n_1687),
.C(n_1645),
.D(n_1673),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1691),
.B(n_1678),
.Y(n_1733)
);

AND2x4_ASAP7_75t_SL g1734 ( 
.A(n_1704),
.B(n_1604),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1706),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1715),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1692),
.B(n_1678),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1702),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1709),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1710),
.B(n_1684),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1704),
.B(n_1715),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1715),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1709),
.Y(n_1743)
);

AND2x4_ASAP7_75t_SL g1744 ( 
.A(n_1704),
.B(n_1604),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1709),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1712),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1718),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1692),
.B(n_1711),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1710),
.B(n_1711),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1722),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1731),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1736),
.Y(n_1754)
);

NOR2x1_ASAP7_75t_L g1755 ( 
.A(n_1720),
.B(n_1700),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1736),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1723),
.B(n_1665),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1739),
.B(n_1696),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1731),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1721),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1729),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1741),
.B(n_1736),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1729),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1735),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1735),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1723),
.B(n_1665),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1722),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1747),
.B(n_1693),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1747),
.B(n_1693),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1724),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1724),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1748),
.B(n_1693),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1726),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1726),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1748),
.B(n_1692),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1727),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1721),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1731),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1738),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1748),
.B(n_1741),
.Y(n_1780)
);

AOI21xp33_ASAP7_75t_L g1781 ( 
.A1(n_1720),
.A2(n_1685),
.B(n_1694),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1736),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1727),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1742),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1742),
.Y(n_1785)
);

INVxp67_ASAP7_75t_SL g1786 ( 
.A(n_1742),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1699),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1738),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1739),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1741),
.B(n_1699),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1743),
.B(n_1701),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1743),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1741),
.B(n_1610),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1742),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_1745),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1779),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1761),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1780),
.Y(n_1798)
);

XOR2xp5_ASAP7_75t_L g1799 ( 
.A(n_1755),
.B(n_1610),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1755),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1780),
.B(n_1732),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1761),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1781),
.B(n_1732),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1793),
.B(n_1615),
.Y(n_1804)
);

NOR2x1p5_ASAP7_75t_L g1805 ( 
.A(n_1757),
.B(n_1766),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1785),
.B(n_1716),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1787),
.B(n_1725),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1762),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1794),
.B(n_1716),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1786),
.B(n_1745),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1754),
.B(n_1746),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1784),
.B(n_1746),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1767),
.B(n_1789),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1789),
.A2(n_1700),
.B1(n_1713),
.B2(n_1689),
.C(n_1705),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1763),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1782),
.B(n_1750),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1763),
.Y(n_1817)
);

NAND4xp25_ASAP7_75t_L g1818 ( 
.A(n_1782),
.B(n_1708),
.C(n_1669),
.D(n_1695),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1787),
.B(n_1790),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1756),
.B(n_1750),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1767),
.B(n_1792),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1725),
.Y(n_1822)
);

NAND4xp25_ASAP7_75t_L g1823 ( 
.A(n_1762),
.B(n_1708),
.C(n_1669),
.D(n_1695),
.Y(n_1823)
);

NOR3xp33_ASAP7_75t_L g1824 ( 
.A(n_1756),
.B(n_1713),
.C(n_1685),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1772),
.B(n_1749),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1762),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1762),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1772),
.B(n_1725),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1775),
.B(n_1728),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1768),
.B(n_1730),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1813),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1813),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1821),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1821),
.Y(n_1834)
);

AOI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1800),
.A2(n_1803),
.B1(n_1814),
.B2(n_1796),
.C(n_1824),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1797),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1805),
.B(n_1768),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1802),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1815),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1806),
.A2(n_1788),
.B(n_1792),
.C(n_1765),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1808),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1808),
.Y(n_1842)
);

AOI322xp5_ASAP7_75t_L g1843 ( 
.A1(n_1809),
.A2(n_1775),
.A3(n_1737),
.B1(n_1728),
.B2(n_1733),
.C1(n_1769),
.C2(n_1707),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1808),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1795),
.B(n_1788),
.Y(n_1845)
);

AOI222xp33_ASAP7_75t_L g1846 ( 
.A1(n_1801),
.A2(n_1769),
.B1(n_1749),
.B2(n_1682),
.C1(n_1783),
.C2(n_1771),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1799),
.A2(n_1632),
.B(n_1703),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1801),
.A2(n_1668),
.B1(n_1744),
.B2(n_1734),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1826),
.Y(n_1850)
);

INVxp67_ASAP7_75t_SL g1851 ( 
.A(n_1826),
.Y(n_1851)
);

AOI322xp5_ASAP7_75t_L g1852 ( 
.A1(n_1828),
.A2(n_1733),
.A3(n_1737),
.B1(n_1728),
.B2(n_1714),
.C1(n_1707),
.C2(n_1699),
.Y(n_1852)
);

OAI21xp33_ASAP7_75t_L g1853 ( 
.A1(n_1823),
.A2(n_1818),
.B(n_1827),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1795),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1798),
.B(n_1770),
.Y(n_1855)
);

CKINVDCx16_ASAP7_75t_R g1856 ( 
.A(n_1804),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_L g1857 ( 
.A(n_1810),
.B(n_1771),
.C(n_1770),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1841),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1854),
.B(n_1798),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1851),
.Y(n_1860)
);

AOI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1835),
.A2(n_1816),
.B1(n_1820),
.B2(n_1812),
.C(n_1811),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1853),
.A2(n_1830),
.B1(n_1819),
.B2(n_1826),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1856),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1837),
.B(n_1804),
.Y(n_1864)
);

OAI222xp33_ASAP7_75t_L g1865 ( 
.A1(n_1848),
.A2(n_1825),
.B1(n_1829),
.B2(n_1819),
.C1(n_1830),
.C2(n_1822),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1841),
.Y(n_1866)
);

OAI21xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1846),
.A2(n_1822),
.B(n_1807),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1851),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1831),
.Y(n_1869)
);

BUFx2_ASAP7_75t_SL g1870 ( 
.A(n_1842),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1857),
.A2(n_1705),
.B1(n_1703),
.B2(n_1830),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1842),
.B(n_1807),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1831),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1832),
.B(n_1828),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1845),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1833),
.B(n_1773),
.Y(n_1877)
);

AOI222xp33_ASAP7_75t_L g1878 ( 
.A1(n_1834),
.A2(n_1773),
.B1(n_1783),
.B2(n_1774),
.C1(n_1776),
.C2(n_1765),
.Y(n_1878)
);

XNOR2x2_ASAP7_75t_L g1879 ( 
.A(n_1863),
.B(n_1844),
.Y(n_1879)
);

NOR2x1_ASAP7_75t_L g1880 ( 
.A(n_1860),
.B(n_1844),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1849),
.Y(n_1881)
);

NAND2x1_ASAP7_75t_L g1882 ( 
.A(n_1868),
.B(n_1850),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1862),
.A2(n_1850),
.B1(n_1855),
.B2(n_1838),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1870),
.B(n_1840),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1858),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1872),
.B(n_1843),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1858),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1866),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1871),
.A2(n_1847),
.B1(n_1839),
.B2(n_1836),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1866),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1861),
.A2(n_1705),
.B1(n_1703),
.B2(n_1626),
.Y(n_1891)
);

NAND4xp75_ASAP7_75t_L g1892 ( 
.A(n_1880),
.B(n_1867),
.C(n_1869),
.D(n_1873),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1879),
.Y(n_1893)
);

NAND2xp33_ASAP7_75t_SL g1894 ( 
.A(n_1882),
.B(n_1872),
.Y(n_1894)
);

AOI211xp5_ASAP7_75t_L g1895 ( 
.A1(n_1889),
.A2(n_1865),
.B(n_1864),
.C(n_1859),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1885),
.Y(n_1896)
);

NAND3xp33_ASAP7_75t_L g1897 ( 
.A(n_1884),
.B(n_1889),
.C(n_1883),
.Y(n_1897)
);

OAI321xp33_ASAP7_75t_L g1898 ( 
.A1(n_1886),
.A2(n_1871),
.A3(n_1874),
.B1(n_1876),
.B2(n_1875),
.C(n_1877),
.Y(n_1898)
);

AOI211xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1881),
.A2(n_1877),
.B(n_1774),
.C(n_1776),
.Y(n_1899)
);

A2O1A1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1891),
.A2(n_1852),
.B(n_1718),
.C(n_1764),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1893),
.A2(n_1888),
.B(n_1887),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1894),
.Y(n_1902)
);

AOI322xp5_ASAP7_75t_L g1903 ( 
.A1(n_1898),
.A2(n_1890),
.A3(n_1737),
.B1(n_1733),
.B2(n_1878),
.C1(n_1764),
.C2(n_1714),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1895),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1896),
.Y(n_1905)
);

AOI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1904),
.A2(n_1897),
.B1(n_1900),
.B2(n_1892),
.C(n_1899),
.Y(n_1906)
);

XNOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1905),
.B(n_1668),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1902),
.A2(n_1751),
.B1(n_1730),
.B2(n_1703),
.Y(n_1908)
);

NOR4xp75_ASAP7_75t_L g1909 ( 
.A(n_1903),
.B(n_1718),
.C(n_1760),
.D(n_1777),
.Y(n_1909)
);

OAI221xp5_ASAP7_75t_SL g1910 ( 
.A1(n_1901),
.A2(n_1791),
.B1(n_1758),
.B2(n_1645),
.C(n_1753),
.Y(n_1910)
);

OAI311xp33_ASAP7_75t_L g1911 ( 
.A1(n_1902),
.A2(n_1758),
.A3(n_1791),
.B1(n_1760),
.C1(n_1777),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1907),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1906),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1910),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1908),
.B(n_1753),
.Y(n_1915)
);

XNOR2xp5_ASAP7_75t_L g1916 ( 
.A(n_1909),
.B(n_1593),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1913),
.B(n_1911),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_SL g1918 ( 
.A(n_1912),
.B(n_1740),
.C(n_1597),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1914),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1917),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1920),
.A2(n_1919),
.B1(n_1916),
.B2(n_1915),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1921),
.Y(n_1922)
);

OA21x2_ASAP7_75t_L g1923 ( 
.A1(n_1921),
.A2(n_1918),
.B(n_1759),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1923),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1923),
.Y(n_1925)
);

AO22x2_ASAP7_75t_SL g1926 ( 
.A1(n_1925),
.A2(n_1922),
.B1(n_1923),
.B2(n_1753),
.Y(n_1926)
);

OAI22xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1924),
.A2(n_1778),
.B1(n_1759),
.B2(n_1760),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1927),
.A2(n_1778),
.B1(n_1759),
.B2(n_1760),
.Y(n_1928)
);

AO21x2_ASAP7_75t_L g1929 ( 
.A1(n_1928),
.A2(n_1926),
.B(n_1778),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1929),
.Y(n_1930)
);

AOI221xp5_ASAP7_75t_L g1931 ( 
.A1(n_1930),
.A2(n_1777),
.B1(n_1730),
.B2(n_1751),
.C(n_1721),
.Y(n_1931)
);

AOI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1931),
.A2(n_1594),
.B(n_1596),
.C(n_1598),
.Y(n_1932)
);


endmodule