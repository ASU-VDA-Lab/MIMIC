module fake_ariane_3265_n_2078 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2078);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2078;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_279;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_1083;
wire n_274;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1856;
wire n_1733;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1865;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_246;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_88),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_60),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_106),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_15),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_60),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_97),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_12),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_174),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_39),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_16),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_61),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_104),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_150),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_75),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_26),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_149),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_71),
.Y(n_238)
);

BUFx8_ASAP7_75t_SL g239 ( 
.A(n_191),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_12),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_46),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_21),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_199),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_82),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_69),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_186),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_61),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_25),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_107),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_156),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_105),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_167),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_76),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_133),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_79),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_44),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_54),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_17),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_102),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_42),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_52),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_41),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_101),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_163),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_98),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_74),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_36),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_201),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_99),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_65),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_1),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_94),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_100),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_33),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_36),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_130),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_24),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_111),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_69),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_165),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_152),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_119),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_128),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_49),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_29),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_49),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_154),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_20),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_41),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_67),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_103),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_40),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_202),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_143),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_38),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_146),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_62),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_51),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_200),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_6),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_67),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_141),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_2),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_136),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_66),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_27),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_11),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_0),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_157),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_147),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_175),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_4),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_112),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_29),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_52),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_179),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_56),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_137),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_159),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_46),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_145),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_114),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_18),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_166),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_24),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_110),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_160),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_9),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_162),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_161),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_93),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_124),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_126),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_50),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_108),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_85),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_113),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_38),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_42),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_169),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_72),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_81),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_53),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_171),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_54),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_187),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_51),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_80),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_28),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_144),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_39),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_115),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_28),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_95),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_31),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_71),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_125),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_194),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_172),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_20),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_34),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_33),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_203),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_91),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_11),
.Y(n_373)
);

BUFx2_ASAP7_75t_SL g374 ( 
.A(n_48),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_178),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_62),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_183),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_122),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_30),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_37),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_6),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_185),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_65),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_89),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_9),
.Y(n_385)
);

BUFx8_ASAP7_75t_SL g386 ( 
.A(n_48),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_120),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_53),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_138),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_37),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_27),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_35),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_139),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_196),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_47),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_208),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_109),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_116),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_204),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_127),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_181),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_140),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_182),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_3),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_64),
.Y(n_405)
);

BUFx10_ASAP7_75t_L g406 ( 
.A(n_58),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_193),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_189),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_45),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_129),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_55),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_177),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_7),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_21),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_56),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_155),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_50),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_210),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_267),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_386),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_248),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_272),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_267),
.B(n_0),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_267),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_356),
.B(n_3),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_297),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_226),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_297),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_348),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_243),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_220),
.B(n_4),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_220),
.B(n_241),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_369),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_263),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_217),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_241),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_343),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_238),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_238),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_225),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_238),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_238),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_238),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_269),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_261),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_405),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_240),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_269),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_269),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_250),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_276),
.B(n_5),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_326),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_261),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_213),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_214),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_326),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_326),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_277),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_352),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_216),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_217),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_414),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_352),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_221),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_239),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_352),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_212),
.B(n_7),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_250),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_255),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_211),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_235),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_261),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_276),
.B(n_8),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_368),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_344),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_242),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_368),
.B(n_8),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_261),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_273),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_411),
.B(n_10),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_211),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_215),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_393),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_300),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_308),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_215),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_221),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_367),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_311),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_367),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_250),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_322),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_323),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_382),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_336),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_257),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_342),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_353),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_219),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_285),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_382),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_219),
.Y(n_509)
);

INVxp33_ASAP7_75t_SL g510 ( 
.A(n_223),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_223),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_355),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_218),
.B(n_10),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_363),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_222),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_285),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_261),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_325),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_222),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_394),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_228),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_394),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_224),
.B(n_230),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_285),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_251),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_503),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

BUFx12f_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_459),
.B(n_249),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_475),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_427),
.B(n_252),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_450),
.B(n_406),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_444),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_444),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_422),
.B(n_253),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_503),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_419),
.B(n_227),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_447),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_503),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_445),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_448),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_419),
.B(n_227),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_445),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_511),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_448),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_449),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_449),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_451),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_424),
.B(n_233),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_452),
.B(n_233),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_523),
.B(n_258),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_426),
.B(n_259),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_478),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_478),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_484),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_484),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_517),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_517),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_518),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_429),
.B(n_315),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_473),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_422),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_525),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_438),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_438),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_431),
.B(n_315),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_460),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_471),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_461),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_433),
.B(n_390),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_466),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_436),
.B(n_265),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_477),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_482),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_485),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_425),
.B(n_268),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_490),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_434),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_476),
.B(n_325),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_496),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_437),
.B(n_284),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_441),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_428),
.B(n_390),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_500),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_502),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_504),
.B(n_325),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_430),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_512),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_457),
.B(n_229),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_430),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_479),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_432),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_486),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_421),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_450),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_435),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_442),
.B(n_312),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_440),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_599),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_568),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_571),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_534),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_603),
.B(n_432),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_554),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_531),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_603),
.B(n_476),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_534),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_603),
.B(n_487),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_571),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_568),
.B(n_454),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_601),
.B(n_487),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_567),
.B(n_488),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_568),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_554),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_567),
.B(n_488),
.Y(n_628)
);

AO22x1_ASAP7_75t_L g629 ( 
.A1(n_601),
.A2(n_494),
.B1(n_510),
.B2(n_470),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_607),
.B(n_493),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_568),
.B(n_454),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_535),
.Y(n_632)
);

INVx4_ASAP7_75t_SL g633 ( 
.A(n_601),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_554),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_535),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_539),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_539),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_599),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_541),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_571),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_541),
.Y(n_641)
);

BUFx8_ASAP7_75t_SL g642 ( 
.A(n_528),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_607),
.B(n_493),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_571),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_599),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_571),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_570),
.B(n_455),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_571),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_601),
.A2(n_483),
.B1(n_467),
.B2(n_495),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_572),
.Y(n_650)
);

OAI21xp33_ASAP7_75t_SL g651 ( 
.A1(n_557),
.A2(n_492),
.B(n_480),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_544),
.Y(n_652)
);

AND2x4_ASAP7_75t_SL g653 ( 
.A(n_607),
.B(n_481),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_544),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_533),
.A2(n_509),
.B1(n_515),
.B2(n_506),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_554),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_572),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_549),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_587),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_607),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_548),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_570),
.B(n_455),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_549),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_550),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_607),
.B(n_506),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_531),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_550),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_572),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_593),
.A2(n_509),
.B1(n_519),
.B2(n_515),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_562),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_607),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_572),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_562),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_572),
.Y(n_674)
);

NAND2xp33_ASAP7_75t_R g675 ( 
.A(n_597),
.B(n_458),
.Y(n_675)
);

NAND2x1p5_ASAP7_75t_L g676 ( 
.A(n_546),
.B(n_324),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_593),
.B(n_507),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_538),
.B(n_456),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_548),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_572),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_607),
.B(n_519),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_551),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_605),
.B(n_458),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_572),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_538),
.B(n_545),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_605),
.B(n_462),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_599),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_562),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_563),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_599),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_552),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_563),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_551),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_605),
.B(n_521),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_606),
.B(n_423),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_558),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_563),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_601),
.A2(n_501),
.B1(n_508),
.B2(n_497),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_605),
.B(n_462),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_558),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_605),
.B(n_463),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_577),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_SL g705 ( 
.A(n_597),
.B(n_521),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_543),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_559),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_543),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_559),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_599),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_560),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_552),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_543),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_533),
.B(n_463),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_547),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_599),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_547),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_547),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_605),
.B(n_465),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_605),
.B(n_465),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_600),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_601),
.A2(n_522),
.B1(n_520),
.B2(n_381),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_557),
.B(n_469),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_560),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_546),
.B(n_469),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_552),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_552),
.Y(n_727)
);

BUFx4f_ASAP7_75t_L g728 ( 
.A(n_601),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_593),
.B(n_262),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_552),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_608),
.B(n_472),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_584),
.B(n_472),
.C(n_260),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_564),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_608),
.B(n_474),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_600),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_610),
.B(n_580),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_546),
.B(n_498),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_593),
.B(n_364),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_606),
.B(n_516),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_552),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_577),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_546),
.B(n_489),
.Y(n_742)
);

AND3x1_ASAP7_75t_L g743 ( 
.A(n_530),
.B(n_392),
.C(n_383),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_569),
.B(n_553),
.Y(n_744)
);

INVx5_ASAP7_75t_L g745 ( 
.A(n_526),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_610),
.B(n_580),
.Y(n_746)
);

XNOR2xp5_ASAP7_75t_L g747 ( 
.A(n_576),
.B(n_446),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_552),
.Y(n_748)
);

XOR2xp5_ASAP7_75t_L g749 ( 
.A(n_602),
.B(n_439),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_561),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_564),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_528),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_565),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_561),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_601),
.A2(n_395),
.B1(n_404),
.B2(n_413),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_565),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_546),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_561),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_593),
.B(n_409),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_546),
.B(n_282),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_561),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_556),
.B(n_335),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_569),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_615),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_677),
.B(n_555),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_728),
.B(n_602),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_619),
.B(n_593),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_683),
.B(n_601),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_642),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_755),
.A2(n_556),
.B1(n_582),
.B2(n_577),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_621),
.B(n_555),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_728),
.B(n_604),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_723),
.A2(n_588),
.B1(n_530),
.B2(n_574),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_706),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_615),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_L g776 ( 
.A(n_686),
.B(n_574),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_620),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_728),
.B(n_604),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_736),
.A2(n_579),
.B(n_581),
.C(n_575),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_647),
.B(n_529),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_695),
.B(n_600),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_620),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_662),
.B(n_746),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_625),
.A2(n_592),
.B1(n_536),
.B2(n_555),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_762),
.B(n_529),
.Y(n_785)
);

AND2x6_ASAP7_75t_L g786 ( 
.A(n_738),
.B(n_538),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_628),
.B(n_592),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_632),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_616),
.B(n_592),
.Y(n_789)
);

BUFx8_ASAP7_75t_L g790 ( 
.A(n_661),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_618),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_666),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_708),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_701),
.B(n_600),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_632),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_635),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_703),
.B(n_536),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_635),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_719),
.B(n_600),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_720),
.B(n_600),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_617),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_661),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_677),
.B(n_575),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_636),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_685),
.B(n_700),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_677),
.B(n_579),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_685),
.B(n_738),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_636),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_700),
.B(n_600),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_660),
.B(n_725),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_700),
.B(n_596),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_708),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_623),
.B(n_596),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_637),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_763),
.B(n_553),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_637),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_639),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_763),
.B(n_553),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_631),
.B(n_596),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_639),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_655),
.A2(n_251),
.B1(n_331),
.B2(n_260),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_624),
.A2(n_582),
.B(n_590),
.C(n_585),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_624),
.A2(n_581),
.B(n_586),
.C(n_583),
.Y(n_823)
);

OAI221xp5_ASAP7_75t_L g824 ( 
.A1(n_649),
.A2(n_609),
.B1(n_351),
.B2(n_388),
.C(n_245),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_629),
.B(n_738),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_659),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_729),
.A2(n_759),
.B1(n_744),
.B2(n_609),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_713),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_713),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_629),
.B(n_737),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_SL g831 ( 
.A(n_752),
.B(n_528),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_641),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_641),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_715),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_652),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_626),
.B(n_583),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_715),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_714),
.B(n_586),
.Y(n_838)
);

AO22x2_ASAP7_75t_L g839 ( 
.A1(n_749),
.A2(n_722),
.B1(n_669),
.B2(n_744),
.Y(n_839)
);

OAI22xp33_ASAP7_75t_L g840 ( 
.A1(n_729),
.A2(n_532),
.B1(n_585),
.B2(n_582),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_652),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_671),
.B(n_228),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_617),
.Y(n_843)
);

AOI22x1_ASAP7_75t_L g844 ( 
.A1(n_627),
.A2(n_634),
.B1(n_656),
.B2(n_654),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_704),
.B(n_589),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_633),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_654),
.Y(n_847)
);

INVx8_ASAP7_75t_L g848 ( 
.A(n_752),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_749),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_717),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_658),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_684),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_684),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_705),
.B(n_420),
.C(n_333),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_741),
.B(n_613),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_611),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_718),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_759),
.A2(n_585),
.B1(n_594),
.B2(n_590),
.Y(n_858)
);

NOR2x1p5_ASAP7_75t_L g859 ( 
.A(n_739),
.B(n_589),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_613),
.B(n_678),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_718),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_658),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_671),
.B(n_232),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_670),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_663),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_633),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_678),
.B(n_759),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_659),
.Y(n_868)
);

CKINVDCx11_ASAP7_75t_R g869 ( 
.A(n_679),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_SL g870 ( 
.A(n_696),
.B(n_443),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_673),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_651),
.A2(n_590),
.B(n_594),
.C(n_532),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_653),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_663),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_664),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_759),
.B(n_595),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_627),
.B(n_595),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_664),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_667),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_634),
.B(n_598),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_732),
.B(n_598),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_673),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_667),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_729),
.A2(n_594),
.B1(n_578),
.B2(n_573),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_671),
.B(n_232),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_675),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_742),
.B(n_591),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_729),
.B(n_591),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_731),
.B(n_566),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_653),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_688),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_SL g892 ( 
.A1(n_679),
.A2(n_464),
.B1(n_468),
.B2(n_453),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_656),
.B(n_630),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_643),
.B(n_545),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_665),
.A2(n_545),
.B1(n_345),
.B2(n_237),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_633),
.B(n_234),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_682),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_681),
.B(n_566),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_633),
.B(n_234),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_696),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_682),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_SL g902 ( 
.A1(n_699),
.A2(n_524),
.B1(n_379),
.B2(n_415),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_694),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_694),
.B(n_566),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_611),
.B(n_236),
.Y(n_905)
);

NAND3xp33_ASAP7_75t_L g906 ( 
.A(n_739),
.B(n_333),
.C(n_331),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_734),
.B(n_573),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_697),
.B(n_573),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_611),
.B(n_236),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_697),
.B(n_578),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_611),
.B(n_638),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_747),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_702),
.B(n_707),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_743),
.A2(n_349),
.B1(n_346),
.B2(n_347),
.C(n_357),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_702),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_707),
.B(n_578),
.Y(n_916)
);

OAI22xp33_ASAP7_75t_L g917 ( 
.A1(n_709),
.A2(n_349),
.B1(n_346),
.B2(n_347),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_688),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_709),
.B(n_573),
.Y(n_919)
);

BUFx8_ASAP7_75t_L g920 ( 
.A(n_747),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_711),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_690),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_611),
.B(n_237),
.Y(n_923)
);

BUFx6f_ASAP7_75t_SL g924 ( 
.A(n_711),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_760),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_724),
.B(n_573),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_638),
.B(n_244),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_660),
.A2(n_357),
.B1(n_359),
.B2(n_361),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_690),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_724),
.B(n_578),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_687),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_733),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_638),
.B(n_244),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_783),
.B(n_733),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_783),
.B(n_751),
.Y(n_935)
);

INVx3_ASAP7_75t_SL g936 ( 
.A(n_769),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_799),
.A2(n_644),
.B(n_640),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_768),
.A2(n_800),
.B(n_794),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_846),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_780),
.B(n_751),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_791),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_780),
.B(n_753),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_794),
.A2(n_800),
.B(n_913),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_781),
.A2(n_668),
.B(n_657),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_805),
.B(n_753),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_793),
.Y(n_946)
);

BUFx8_ASAP7_75t_L g947 ( 
.A(n_924),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_781),
.A2(n_672),
.B(n_689),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_765),
.B(n_578),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_822),
.A2(n_756),
.B(n_676),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_815),
.B(n_406),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_868),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_787),
.A2(n_756),
.B1(n_676),
.B2(n_689),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_793),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_787),
.B(n_693),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_837),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_771),
.B(n_693),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_785),
.B(n_698),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_887),
.B(n_698),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_869),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_904),
.A2(n_779),
.B(n_767),
.C(n_908),
.Y(n_961)
);

BUFx4f_ASAP7_75t_L g962 ( 
.A(n_848),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_887),
.B(n_676),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_797),
.A2(n_757),
.B(n_689),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_888),
.A2(n_881),
.B(n_838),
.C(n_823),
.Y(n_965)
);

NAND2x1_ASAP7_75t_L g966 ( 
.A(n_846),
.B(n_692),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_911),
.A2(n_757),
.B(n_646),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_802),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_852),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_911),
.A2(n_757),
.B(n_646),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_764),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_810),
.A2(n_646),
.B(n_622),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_837),
.Y(n_973)
);

NOR2x1p5_ASAP7_75t_L g974 ( 
.A(n_867),
.B(n_359),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_888),
.B(n_687),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_809),
.A2(n_648),
.B(n_622),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_813),
.A2(n_819),
.B(n_855),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_827),
.B(n_638),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_886),
.B(n_692),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_807),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_822),
.A2(n_789),
.B(n_836),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_893),
.A2(n_863),
.B(n_842),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_827),
.A2(n_716),
.B1(n_721),
.B2(n_691),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_910),
.A2(n_761),
.B(n_692),
.C(n_712),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_818),
.B(n_406),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_784),
.B(n_716),
.Y(n_986)
);

OAI22x1_ASAP7_75t_L g987 ( 
.A1(n_859),
.A2(n_361),
.B1(n_373),
.B2(n_376),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_906),
.B(n_266),
.C(n_264),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_807),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_842),
.A2(n_648),
.B(n_622),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_811),
.B(n_721),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_803),
.B(n_638),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_792),
.B(n_712),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_860),
.B(n_773),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_775),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_765),
.B(n_761),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_900),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_866),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_863),
.A2(n_674),
.B(n_648),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_830),
.B(n_825),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_852),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_881),
.A2(n_761),
.B(n_730),
.C(n_712),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_916),
.A2(n_730),
.B(n_748),
.C(n_750),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_803),
.B(n_645),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_866),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_786),
.B(n_730),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_885),
.A2(n_880),
.B(n_877),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_838),
.A2(n_748),
.B(n_750),
.C(n_754),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_919),
.A2(n_750),
.B(n_748),
.C(n_674),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_824),
.B(n_612),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_777),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_786),
.B(n_674),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_924),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_900),
.B(n_373),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_782),
.A2(n_612),
.B1(n_650),
.B2(n_614),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_885),
.A2(n_680),
.B(n_614),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_806),
.B(n_884),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_840),
.B(n_645),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_872),
.A2(n_727),
.B(n_726),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_845),
.A2(n_680),
.B(n_614),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_806),
.B(n_884),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_788),
.A2(n_612),
.B1(n_650),
.B2(n_680),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_786),
.B(n_645),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_786),
.B(n_645),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_801),
.Y(n_1025)
);

AOI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_839),
.A2(n_727),
.B(n_726),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_801),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_930),
.A2(n_758),
.B(n_754),
.C(n_740),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_843),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_795),
.A2(n_650),
.B1(n_735),
.B2(n_710),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_852),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_SL g1032 ( 
.A1(n_796),
.A2(n_758),
.B(n_740),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_786),
.B(n_645),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_896),
.A2(n_537),
.B(n_527),
.Y(n_1034)
);

AOI22x1_ASAP7_75t_L g1035 ( 
.A1(n_798),
.A2(n_691),
.B1(n_735),
.B2(n_710),
.Y(n_1035)
);

AOI22x1_ASAP7_75t_L g1036 ( 
.A1(n_804),
.A2(n_691),
.B1(n_735),
.B2(n_710),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_926),
.B(n_691),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_872),
.A2(n_745),
.B(n_334),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_808),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_365),
.B(n_396),
.C(n_377),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_843),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_SL g1042 ( 
.A1(n_814),
.A2(n_330),
.B(n_338),
.C(n_339),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_889),
.B(n_691),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_816),
.A2(n_735),
.B(n_710),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_817),
.A2(n_735),
.B(n_710),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_SL g1046 ( 
.A(n_856),
.B(n_376),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_820),
.A2(n_745),
.B(n_254),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_832),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_844),
.A2(n_745),
.B(n_358),
.Y(n_1049)
);

NAND2xp33_ASAP7_75t_L g1050 ( 
.A(n_856),
.B(n_745),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_870),
.B(n_379),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_833),
.A2(n_745),
.B(n_254),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_835),
.A2(n_256),
.B(n_247),
.Y(n_1053)
);

BUFx5_ASAP7_75t_L g1054 ( 
.A(n_841),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_914),
.B(n_281),
.C(n_280),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_826),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_889),
.B(n_380),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_766),
.B(n_247),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_873),
.B(n_340),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_847),
.A2(n_329),
.B(n_256),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_851),
.A2(n_332),
.B(n_329),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_862),
.A2(n_341),
.B(n_332),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_766),
.B(n_341),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_852),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_865),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_874),
.B(n_380),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_875),
.Y(n_1067)
);

NAND2x1_ASAP7_75t_L g1068 ( 
.A(n_856),
.B(n_561),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_772),
.B(n_366),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_772),
.B(n_778),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_778),
.B(n_391),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_774),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_812),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_878),
.B(n_391),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_876),
.B(n_415),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_907),
.B(n_283),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_879),
.B(n_287),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_883),
.B(n_292),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_790),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_897),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_901),
.B(n_293),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_790),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_903),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_920),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_SL g1085 ( 
.A(n_831),
.B(n_362),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_915),
.A2(n_372),
.B(n_384),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_SL g1087 ( 
.A1(n_921),
.A2(n_403),
.B(n_401),
.C(n_416),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_932),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_776),
.A2(n_931),
.B(n_909),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_840),
.B(n_345),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_907),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_917),
.B(n_306),
.C(n_305),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_828),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_931),
.A2(n_354),
.B(n_375),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_853),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_925),
.B(n_294),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_858),
.A2(n_309),
.B1(n_316),
.B2(n_328),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_848),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_890),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_896),
.A2(n_527),
.B(n_542),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_898),
.B(n_296),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_853),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_853),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_894),
.B(n_770),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_858),
.B(n_229),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_905),
.A2(n_354),
.B(n_375),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_895),
.A2(n_246),
.B(n_278),
.C(n_371),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_905),
.A2(n_360),
.B(n_384),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_853),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_899),
.A2(n_527),
.B(n_542),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_909),
.A2(n_360),
.B(n_387),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_770),
.B(n_298),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_856),
.B(n_848),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_929),
.B(n_303),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_899),
.A2(n_537),
.B(n_542),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_912),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_917),
.B(n_313),
.Y(n_1117)
);

AOI21x1_ASAP7_75t_L g1118 ( 
.A1(n_864),
.A2(n_540),
.B(n_537),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_839),
.A2(n_320),
.B1(n_314),
.B2(n_385),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_923),
.A2(n_372),
.B(n_397),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_902),
.B(n_378),
.Y(n_1121)
);

NOR2xp67_ASAP7_75t_SL g1122 ( 
.A(n_923),
.B(n_325),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_968),
.B(n_849),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_934),
.B(n_839),
.Y(n_1124)
);

AO21x2_ASAP7_75t_L g1125 ( 
.A1(n_1000),
.A2(n_933),
.B(n_927),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_938),
.A2(n_891),
.B(n_871),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_971),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_936),
.Y(n_1128)
);

AND2x2_ASAP7_75t_SL g1129 ( 
.A(n_1092),
.B(n_854),
.Y(n_1129)
);

AO21x1_ASAP7_75t_L g1130 ( 
.A1(n_963),
.A2(n_933),
.B(n_927),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_935),
.B(n_882),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1121),
.A2(n_1092),
.B1(n_1076),
.B2(n_1119),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_940),
.A2(n_918),
.B(n_922),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_SL g1134 ( 
.A(n_939),
.B(n_920),
.Y(n_1134)
);

CKINVDCx16_ASAP7_75t_R g1135 ( 
.A(n_960),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_942),
.A2(n_928),
.B1(n_821),
.B2(n_325),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_968),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_969),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_946),
.Y(n_1139)
);

CKINVDCx14_ASAP7_75t_R g1140 ( 
.A(n_952),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_949),
.B(n_829),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_959),
.A2(n_834),
.B(n_861),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_962),
.B(n_892),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_995),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_962),
.B(n_849),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_965),
.A2(n_945),
.B1(n_1091),
.B2(n_994),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_994),
.B(n_850),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1091),
.B(n_378),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_945),
.A2(n_385),
.B1(n_417),
.B2(n_857),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_939),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1011),
.Y(n_1151)
);

AO22x1_ASAP7_75t_L g1152 ( 
.A1(n_1121),
.A2(n_407),
.B1(n_389),
.B2(n_397),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_SL g1153 ( 
.A1(n_1046),
.A2(n_1009),
.B(n_1003),
.C(n_984),
.Y(n_1153)
);

AOI22x1_ASAP7_75t_L g1154 ( 
.A1(n_977),
.A2(n_981),
.B1(n_1052),
.B2(n_1047),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1084),
.B(n_231),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1076),
.A2(n_231),
.B(n_246),
.C(n_278),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_955),
.A2(n_371),
.B(n_275),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_958),
.B(n_561),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1055),
.A2(n_387),
.B1(n_389),
.B2(n_398),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_961),
.A2(n_410),
.B(n_400),
.C(n_402),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_949),
.B(n_561),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1039),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1104),
.B(n_398),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_953),
.A2(n_950),
.B(n_964),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_969),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_R g1166 ( 
.A(n_936),
.B(n_399),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_947),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_957),
.B(n_399),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1048),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1065),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_954),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_SL g1172 ( 
.A(n_1079),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_969),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_947),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1075),
.B(n_400),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1056),
.A2(n_402),
.B1(n_407),
.B2(n_408),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1013),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_956),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_969),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_997),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1067),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1037),
.A2(n_307),
.B(n_270),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_943),
.A2(n_310),
.B(n_271),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1080),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_997),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_951),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_980),
.B(n_540),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1117),
.A2(n_540),
.B(n_14),
.C(n_15),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1083),
.B(n_408),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_998),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_941),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1088),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_980),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_973),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_961),
.A2(n_304),
.B(n_418),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1075),
.B(n_410),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1055),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1013),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_985),
.B(n_412),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1072),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1073),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1007),
.A2(n_301),
.B(n_274),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1057),
.A2(n_417),
.B1(n_385),
.B2(n_412),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1014),
.B(n_385),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_989),
.B(n_279),
.Y(n_1205)
);

INVx8_ASAP7_75t_L g1206 ( 
.A(n_1059),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1051),
.B(n_989),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1085),
.B(n_286),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_941),
.Y(n_1209)
);

OA22x2_ASAP7_75t_L g1210 ( 
.A1(n_987),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1082),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1116),
.B(n_291),
.Y(n_1212)
);

OA22x2_ASAP7_75t_L g1213 ( 
.A1(n_1017),
.A2(n_295),
.B1(n_299),
.B2(n_302),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_976),
.A2(n_321),
.B(n_317),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1059),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1044),
.A2(n_327),
.B(n_318),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_SL g1217 ( 
.A1(n_1082),
.A2(n_385),
.B1(n_417),
.B2(n_319),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1116),
.B(n_13),
.Y(n_1218)
);

AO32x2_ASAP7_75t_L g1219 ( 
.A1(n_1030),
.A2(n_417),
.A3(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1070),
.A2(n_417),
.B(n_350),
.C(n_257),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1021),
.B(n_17),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1071),
.B(n_19),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1045),
.A2(n_350),
.B(n_257),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1093),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1098),
.B(n_22),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1071),
.B(n_23),
.Y(n_1226)
);

CKINVDCx8_ASAP7_75t_R g1227 ( 
.A(n_1001),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1105),
.A2(n_257),
.B1(n_350),
.B2(n_32),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_974),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1025),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1105),
.A2(n_257),
.B1(n_350),
.B2(n_32),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1070),
.A2(n_350),
.B1(n_526),
.B2(n_34),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1027),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1029),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1099),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1041),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1020),
.A2(n_526),
.B(n_86),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1099),
.Y(n_1238)
);

OR2x6_ASAP7_75t_SL g1239 ( 
.A(n_1097),
.B(n_25),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1040),
.B(n_526),
.C(n_35),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_1122),
.A2(n_31),
.B(n_40),
.C(n_43),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1101),
.B(n_43),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1054),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1096),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_979),
.B(n_44),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_998),
.Y(n_1246)
);

AO21x1_ASAP7_75t_L g1247 ( 
.A1(n_1038),
.A2(n_92),
.B(n_207),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_979),
.B(n_45),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1001),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1066),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1074),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1001),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1077),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1009),
.A2(n_47),
.B(n_55),
.C(n_57),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1031),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_996),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_988),
.A2(n_526),
.B1(n_58),
.B2(n_59),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1054),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1112),
.A2(n_57),
.B1(n_59),
.B2(n_63),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1023),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_988),
.A2(n_63),
.B(n_64),
.C(n_66),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1078),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1113),
.Y(n_1263)
);

OAI211xp5_ASAP7_75t_L g1264 ( 
.A1(n_1081),
.A2(n_68),
.B(n_70),
.C(n_72),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1114),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_982),
.A2(n_526),
.B(n_132),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1054),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_972),
.A2(n_526),
.B(n_134),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1090),
.A2(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1001),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_992),
.A2(n_77),
.B1(n_78),
.B2(n_83),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_967),
.A2(n_84),
.B(n_87),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_970),
.A2(n_90),
.B(n_96),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1042),
.A2(n_117),
.B1(n_123),
.B2(n_131),
.C(n_135),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1107),
.A2(n_1002),
.B(n_1008),
.C(n_1087),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1054),
.B(n_142),
.Y(n_1276)
);

OR2x6_ASAP7_75t_L g1277 ( 
.A(n_1024),
.B(n_1033),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1010),
.A2(n_151),
.B(n_153),
.C(n_158),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_991),
.A2(n_164),
.B(n_180),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1010),
.B(n_184),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1004),
.B(n_190),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_984),
.A2(n_192),
.B(n_195),
.C(n_1003),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_948),
.A2(n_1050),
.B(n_1016),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1089),
.A2(n_1028),
.B(n_1094),
.C(n_1061),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1031),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1128),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1227),
.Y(n_1287)
);

AO21x1_ASAP7_75t_L g1288 ( 
.A1(n_1146),
.A2(n_978),
.B(n_1018),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1130),
.A2(n_1022),
.A3(n_1015),
.B(n_937),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1211),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_1147),
.B(n_1102),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1138),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1206),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1244),
.B(n_1063),
.Y(n_1294)
);

AO21x1_ASAP7_75t_L g1295 ( 
.A1(n_1146),
.A2(n_1018),
.B(n_1000),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1164),
.A2(n_1028),
.B(n_1043),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1132),
.B(n_1054),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1136),
.A2(n_1032),
.B(n_1019),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1221),
.A2(n_986),
.B1(n_975),
.B2(n_1054),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1283),
.A2(n_1036),
.B(n_1035),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1135),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1127),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1139),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1144),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1126),
.A2(n_1034),
.B(n_1100),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1228),
.A2(n_1012),
.B(n_1103),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1131),
.B(n_1109),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1185),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1222),
.A2(n_1058),
.B(n_1062),
.C(n_1060),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1247),
.A2(n_1282),
.A3(n_1149),
.B(n_1220),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1190),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1280),
.A2(n_1276),
.B(n_1131),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1167),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1226),
.A2(n_1086),
.B(n_1053),
.C(n_1006),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1276),
.A2(n_1049),
.B(n_990),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1180),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1266),
.A2(n_1110),
.B(n_1115),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1151),
.Y(n_1318)
);

OR2x6_ASAP7_75t_L g1319 ( 
.A(n_1206),
.B(n_993),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1137),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1136),
.A2(n_944),
.B(n_999),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1149),
.A2(n_1124),
.A3(n_1142),
.B(n_1231),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1245),
.A2(n_1069),
.B(n_1111),
.C(n_1120),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1237),
.A2(n_1068),
.B(n_1103),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1123),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1154),
.A2(n_1118),
.B(n_1109),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1206),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1207),
.B(n_1108),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_SL g1329 ( 
.A1(n_1153),
.A2(n_966),
.B(n_1106),
.C(n_1026),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1249),
.B(n_1064),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1223),
.A2(n_983),
.B(n_1064),
.Y(n_1331)
);

AO32x2_ASAP7_75t_L g1332 ( 
.A1(n_1228),
.A2(n_1064),
.A3(n_1095),
.B1(n_1103),
.B2(n_1005),
.Y(n_1332)
);

NOR2xp67_ASAP7_75t_L g1333 ( 
.A(n_1270),
.B(n_1150),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1162),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1248),
.A2(n_1005),
.B(n_1064),
.C(n_1095),
.Y(n_1335)
);

INVx3_ASAP7_75t_SL g1336 ( 
.A(n_1198),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1169),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1231),
.A2(n_1095),
.A3(n_1103),
.B(n_1156),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1268),
.A2(n_1095),
.B(n_1275),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1203),
.A2(n_1195),
.B(n_1158),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1191),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1197),
.B(n_1257),
.C(n_1261),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1159),
.A2(n_1129),
.B1(n_1175),
.B2(n_1196),
.Y(n_1343)
);

OA21x2_ASAP7_75t_L g1344 ( 
.A1(n_1133),
.A2(n_1158),
.B(n_1278),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1140),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1284),
.A2(n_1267),
.B(n_1243),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1242),
.A2(n_1262),
.B(n_1253),
.C(n_1232),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1174),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1260),
.B(n_1256),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1260),
.B(n_1256),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1215),
.B(n_1193),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1272),
.A2(n_1273),
.B(n_1258),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1279),
.A2(n_1157),
.B(n_1188),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1190),
.B(n_1177),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1163),
.B(n_1170),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1181),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1163),
.A2(n_1168),
.B(n_1125),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1239),
.A2(n_1250),
.B1(n_1251),
.B2(n_1160),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1171),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1143),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_SL g1361 ( 
.A1(n_1254),
.A2(n_1148),
.B(n_1189),
.C(n_1168),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1184),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1138),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1192),
.B(n_1193),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1138),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1235),
.Y(n_1366)
);

NOR2xp67_ASAP7_75t_L g1367 ( 
.A(n_1150),
.B(n_1246),
.Y(n_1367)
);

AOI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1203),
.A2(n_1240),
.B(n_1213),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1240),
.A2(n_1265),
.B(n_1269),
.C(n_1281),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1178),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1259),
.A2(n_1186),
.B1(n_1152),
.B2(n_1134),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1194),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1202),
.A2(n_1241),
.B(n_1183),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_SL g1374 ( 
.A(n_1134),
.B(n_1172),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1204),
.B(n_1209),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1145),
.B(n_1205),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1125),
.A2(n_1189),
.B(n_1182),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1200),
.A2(n_1201),
.A3(n_1224),
.B(n_1236),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1274),
.A2(n_1214),
.B(n_1246),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1218),
.A2(n_1264),
.B(n_1212),
.C(n_1263),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1277),
.A2(n_1216),
.B(n_1285),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1233),
.A2(n_1234),
.B(n_1271),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1230),
.A2(n_1199),
.B(n_1208),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1172),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1238),
.A2(n_1225),
.B(n_1229),
.C(n_1155),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1213),
.A2(n_1210),
.B(n_1277),
.Y(n_1386)
);

INVx8_ASAP7_75t_L g1387 ( 
.A(n_1161),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1210),
.A2(n_1277),
.B(n_1179),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1165),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1255),
.A2(n_1252),
.B(n_1165),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1165),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1155),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1217),
.A2(n_1225),
.B1(n_1176),
.B2(n_1155),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1141),
.B(n_1252),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1187),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1141),
.B(n_1166),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1161),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1173),
.A2(n_1179),
.B(n_1252),
.Y(n_1398)
);

NOR4xp25_ASAP7_75t_L g1399 ( 
.A(n_1219),
.B(n_1132),
.C(n_1146),
.D(n_1197),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1219),
.A2(n_1130),
.A3(n_1164),
.B(n_1247),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1173),
.B(n_1179),
.Y(n_1401)
);

AO31x2_ASAP7_75t_L g1402 ( 
.A1(n_1219),
.A2(n_1130),
.A3(n_1164),
.B(n_1247),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1173),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1164),
.A2(n_942),
.B(n_940),
.Y(n_1404)
);

AO31x2_ASAP7_75t_L g1405 ( 
.A1(n_1130),
.A2(n_1164),
.A3(n_1247),
.B(n_1282),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1128),
.Y(n_1406)
);

BUFx4f_ASAP7_75t_L g1407 ( 
.A(n_1206),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1211),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1164),
.A2(n_942),
.B(n_940),
.Y(n_1409)
);

AO31x2_ASAP7_75t_L g1410 ( 
.A1(n_1130),
.A2(n_1164),
.A3(n_1247),
.B(n_1282),
.Y(n_1410)
);

INVx5_ASAP7_75t_L g1411 ( 
.A(n_1138),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1244),
.B(n_659),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1164),
.A2(n_1130),
.B(n_1000),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1130),
.A2(n_1164),
.A3(n_1247),
.B(n_1282),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1139),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1211),
.Y(n_1416)
);

NAND3xp33_ASAP7_75t_L g1417 ( 
.A(n_1132),
.B(n_1146),
.C(n_1245),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1146),
.B(n_940),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1146),
.A2(n_783),
.B(n_1092),
.C(n_1222),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1164),
.A2(n_942),
.B(n_940),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1164),
.A2(n_942),
.B(n_940),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1139),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1139),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1239),
.A2(n_533),
.B1(n_1085),
.B2(n_870),
.Y(n_1424)
);

AO32x2_ASAP7_75t_L g1425 ( 
.A1(n_1146),
.A2(n_1119),
.A3(n_1231),
.B1(n_1228),
.B2(n_1136),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1185),
.Y(n_1426)
);

AOI22x1_ASAP7_75t_L g1427 ( 
.A1(n_1195),
.A2(n_605),
.B1(n_603),
.B2(n_607),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1283),
.A2(n_1126),
.B(n_1164),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1164),
.A2(n_1283),
.B(n_1130),
.Y(n_1429)
);

NAND2x1_ASAP7_75t_L g1430 ( 
.A(n_1150),
.B(n_1246),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1283),
.A2(n_1126),
.B(n_1164),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1127),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1180),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1146),
.A2(n_965),
.B(n_963),
.Y(n_1434)
);

AO32x2_ASAP7_75t_L g1435 ( 
.A1(n_1146),
.A2(n_1119),
.A3(n_1231),
.B1(n_1228),
.B2(n_1136),
.Y(n_1435)
);

AO31x2_ASAP7_75t_L g1436 ( 
.A1(n_1130),
.A2(n_1164),
.A3(n_1247),
.B(n_1282),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1146),
.B(n_940),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1227),
.Y(n_1438)
);

AOI31xp67_ASAP7_75t_L g1439 ( 
.A1(n_1280),
.A2(n_1018),
.A3(n_781),
.B(n_800),
.Y(n_1439)
);

CKINVDCx11_ASAP7_75t_R g1440 ( 
.A(n_1128),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1185),
.B(n_783),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1132),
.A2(n_743),
.B1(n_783),
.B2(n_736),
.C(n_746),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1132),
.B(n_1146),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1164),
.A2(n_942),
.B(n_940),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1227),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1283),
.A2(n_1126),
.B(n_1164),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1146),
.A2(n_783),
.B(n_1092),
.C(n_1222),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1128),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1139),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1146),
.A2(n_965),
.B(n_963),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1146),
.A2(n_965),
.B(n_963),
.Y(n_1451)
);

AO31x2_ASAP7_75t_L g1452 ( 
.A1(n_1130),
.A2(n_1164),
.A3(n_1247),
.B(n_1282),
.Y(n_1452)
);

AO31x2_ASAP7_75t_L g1453 ( 
.A1(n_1130),
.A2(n_1164),
.A3(n_1247),
.B(n_1282),
.Y(n_1453)
);

AO31x2_ASAP7_75t_L g1454 ( 
.A1(n_1130),
.A2(n_1164),
.A3(n_1247),
.B(n_1282),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1180),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1139),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1442),
.A2(n_1417),
.B(n_1443),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1417),
.A2(n_1447),
.B(n_1419),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1358),
.A2(n_1343),
.B1(n_1342),
.B2(n_1437),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1358),
.A2(n_1343),
.B1(n_1342),
.B2(n_1437),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1418),
.B(n_1434),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1424),
.A2(n_1368),
.B1(n_1328),
.B2(n_1375),
.Y(n_1462)
);

BUFx2_ASAP7_75t_SL g1463 ( 
.A(n_1345),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1374),
.A2(n_1392),
.B1(n_1418),
.B2(n_1298),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1301),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1368),
.A2(n_1383),
.B1(n_1371),
.B2(n_1396),
.Y(n_1466)
);

CKINVDCx6p67_ASAP7_75t_R g1467 ( 
.A(n_1336),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1290),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1286),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1445),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1434),
.A2(n_1450),
.B1(n_1451),
.B2(n_1441),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1308),
.B(n_1426),
.Y(n_1472)
);

CKINVDCx11_ASAP7_75t_R g1473 ( 
.A(n_1440),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1298),
.A2(n_1450),
.B1(n_1451),
.B2(n_1374),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1294),
.A2(n_1412),
.B1(n_1376),
.B2(n_1384),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1371),
.A2(n_1393),
.B1(n_1325),
.B2(n_1392),
.Y(n_1476)
);

INVx6_ASAP7_75t_L g1477 ( 
.A(n_1445),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1416),
.Y(n_1478)
);

INVx6_ASAP7_75t_L g1479 ( 
.A(n_1445),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1383),
.A2(n_1393),
.B1(n_1359),
.B2(n_1370),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1320),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1308),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1303),
.A2(n_1456),
.B1(n_1372),
.B2(n_1415),
.Y(n_1483)
);

BUFx8_ASAP7_75t_L g1484 ( 
.A(n_1360),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1302),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1422),
.A2(n_1423),
.B1(n_1449),
.B2(n_1349),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1304),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1355),
.A2(n_1407),
.B1(n_1426),
.B2(n_1299),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1348),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1380),
.A2(n_1369),
.B(n_1297),
.Y(n_1490)
);

INVx5_ASAP7_75t_L g1491 ( 
.A(n_1319),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1366),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1407),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1349),
.A2(n_1350),
.B1(n_1288),
.B2(n_1355),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1287),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1318),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1334),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1404),
.A2(n_1421),
.B1(n_1444),
.B2(n_1420),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1409),
.A2(n_1347),
.B1(n_1299),
.B2(n_1433),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1455),
.A2(n_1316),
.B1(n_1323),
.B2(n_1341),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1387),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1313),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1408),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1337),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1356),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1387),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1406),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1362),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1432),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1399),
.A2(n_1327),
.B1(n_1293),
.B2(n_1438),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1319),
.Y(n_1511)
);

OAI21xp33_ASAP7_75t_L g1512 ( 
.A1(n_1399),
.A2(n_1357),
.B(n_1309),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1395),
.Y(n_1513)
);

BUFx10_ASAP7_75t_L g1514 ( 
.A(n_1401),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1386),
.A2(n_1425),
.B1(n_1435),
.B2(n_1388),
.Y(n_1515)
);

BUFx8_ASAP7_75t_L g1516 ( 
.A(n_1448),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1425),
.A2(n_1435),
.B1(n_1350),
.B2(n_1427),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_SL g1518 ( 
.A1(n_1425),
.A2(n_1435),
.B1(n_1312),
.B2(n_1351),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1384),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1307),
.B(n_1295),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1335),
.A2(n_1296),
.B(n_1379),
.Y(n_1521)
);

BUFx4f_ASAP7_75t_L g1522 ( 
.A(n_1354),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1397),
.A2(n_1291),
.B1(n_1382),
.B2(n_1319),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1291),
.A2(n_1382),
.B1(n_1307),
.B2(n_1377),
.Y(n_1524)
);

BUFx10_ASAP7_75t_L g1525 ( 
.A(n_1292),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1394),
.A2(n_1287),
.B1(n_1438),
.B2(n_1413),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1413),
.B(n_1322),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1322),
.B(n_1394),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1403),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1322),
.B(n_1402),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1391),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1391),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1363),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1311),
.A2(n_1367),
.B1(n_1385),
.B2(n_1321),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1381),
.A2(n_1321),
.B1(n_1330),
.B2(n_1344),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1430),
.A2(n_1311),
.B1(n_1429),
.B2(n_1365),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1365),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1332),
.Y(n_1538)
);

OAI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1333),
.A2(n_1367),
.B1(n_1332),
.B2(n_1340),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1332),
.A2(n_1390),
.B1(n_1389),
.B2(n_1398),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1389),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1333),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1338),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1439),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1338),
.B(n_1400),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1338),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1315),
.A2(n_1344),
.B1(n_1331),
.B2(n_1429),
.Y(n_1547)
);

INVx4_ASAP7_75t_SL g1548 ( 
.A(n_1400),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1331),
.Y(n_1549)
);

BUFx10_ASAP7_75t_L g1550 ( 
.A(n_1361),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1400),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1353),
.A2(n_1346),
.B1(n_1373),
.B2(n_1339),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1306),
.A2(n_1314),
.B1(n_1300),
.B2(n_1324),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1402),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1352),
.A2(n_1317),
.B1(n_1305),
.B2(n_1326),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1310),
.A2(n_1454),
.B1(n_1436),
.B2(n_1405),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1310),
.A2(n_1454),
.B1(n_1436),
.B2(n_1405),
.Y(n_1557)
);

BUFx5_ASAP7_75t_L g1558 ( 
.A(n_1428),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1329),
.Y(n_1559)
);

CKINVDCx6p67_ASAP7_75t_R g1560 ( 
.A(n_1405),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1410),
.A2(n_1414),
.B1(n_1436),
.B2(n_1452),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1410),
.A2(n_1414),
.B1(n_1452),
.B2(n_1453),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1289),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1289),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1414),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1453),
.A2(n_1289),
.B1(n_1431),
.B2(n_1446),
.Y(n_1566)
);

INVx6_ASAP7_75t_L g1567 ( 
.A(n_1453),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1424),
.A2(n_839),
.B1(n_1132),
.B2(n_1417),
.Y(n_1568)
);

BUFx8_ASAP7_75t_SL g1569 ( 
.A(n_1301),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1424),
.A2(n_839),
.B1(n_1132),
.B2(n_1417),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1424),
.A2(n_1132),
.B1(n_533),
.B2(n_1442),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1320),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1308),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1417),
.A2(n_839),
.B1(n_1231),
.B2(n_1228),
.Y(n_1574)
);

BUFx4f_ASAP7_75t_SL g1575 ( 
.A(n_1313),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1301),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1417),
.A2(n_1418),
.B1(n_1437),
.B2(n_1442),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1364),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1286),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1411),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1424),
.A2(n_839),
.B1(n_1132),
.B2(n_1417),
.Y(n_1581)
);

OAI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1393),
.A2(n_533),
.B1(n_1239),
.B2(n_1417),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1308),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1424),
.A2(n_839),
.B1(n_1132),
.B2(n_1417),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1393),
.A2(n_533),
.B1(n_1239),
.B2(n_1417),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1301),
.Y(n_1586)
);

BUFx10_ASAP7_75t_L g1587 ( 
.A(n_1412),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1364),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1393),
.A2(n_533),
.B1(n_1239),
.B2(n_1417),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1417),
.A2(n_839),
.B1(n_1231),
.B2(n_1228),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1424),
.A2(n_839),
.B1(n_1132),
.B2(n_1417),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1364),
.Y(n_1592)
);

INVx6_ASAP7_75t_L g1593 ( 
.A(n_1445),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1417),
.A2(n_839),
.B1(n_1231),
.B2(n_1228),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_SL g1595 ( 
.A1(n_1371),
.A2(n_1132),
.B1(n_659),
.B2(n_826),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1364),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1308),
.B(n_997),
.Y(n_1597)
);

NAND2x1p5_ASAP7_75t_L g1598 ( 
.A(n_1407),
.B(n_1445),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1424),
.A2(n_839),
.B1(n_1132),
.B2(n_1417),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1378),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1424),
.A2(n_839),
.B1(n_1132),
.B2(n_1417),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1343),
.A2(n_1239),
.B1(n_1119),
.B2(n_533),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1597),
.B(n_1472),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1528),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1512),
.A2(n_1521),
.B(n_1527),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1602),
.A2(n_1577),
.B1(n_1595),
.B2(n_1471),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1540),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1553),
.A2(n_1566),
.B(n_1561),
.Y(n_1608)
);

INVx4_ASAP7_75t_SL g1609 ( 
.A(n_1565),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1520),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1520),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1459),
.B(n_1460),
.Y(n_1612)
);

CKINVDCx6p67_ASAP7_75t_R g1613 ( 
.A(n_1465),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1569),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1551),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1530),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1530),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1548),
.B(n_1461),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1527),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1538),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1482),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1485),
.B(n_1487),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1565),
.Y(n_1625)
);

INVx2_ASAP7_75t_SL g1626 ( 
.A(n_1573),
.Y(n_1626)
);

INVx4_ASAP7_75t_SL g1627 ( 
.A(n_1565),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1457),
.A2(n_1577),
.B(n_1460),
.Y(n_1629)
);

AO31x2_ASAP7_75t_L g1630 ( 
.A1(n_1561),
.A2(n_1546),
.A3(n_1566),
.B(n_1554),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1491),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1468),
.Y(n_1632)
);

OAI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1521),
.A2(n_1553),
.B(n_1498),
.Y(n_1633)
);

AO21x2_ASAP7_75t_L g1634 ( 
.A1(n_1547),
.A2(n_1557),
.B(n_1539),
.Y(n_1634)
);

AO31x2_ASAP7_75t_L g1635 ( 
.A1(n_1498),
.A2(n_1544),
.A3(n_1600),
.B(n_1563),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1504),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1505),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1567),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1471),
.B(n_1583),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1640)
);

AOI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1499),
.A2(n_1534),
.B(n_1500),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1560),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1545),
.Y(n_1643)
);

AO21x2_ASAP7_75t_L g1644 ( 
.A1(n_1458),
.A2(n_1564),
.B(n_1488),
.Y(n_1644)
);

BUFx2_ASAP7_75t_SL g1645 ( 
.A(n_1491),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1549),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1548),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1457),
.A2(n_1589),
.B(n_1585),
.C(n_1582),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1548),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1549),
.Y(n_1650)
);

AO21x1_ASAP7_75t_SL g1651 ( 
.A1(n_1458),
.A2(n_1535),
.B(n_1571),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1552),
.A2(n_1555),
.B(n_1524),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1543),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1567),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1499),
.A2(n_1534),
.B(n_1500),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1523),
.A2(n_1526),
.B(n_1466),
.Y(n_1656)
);

AOI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1542),
.A2(n_1531),
.B(n_1532),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1556),
.B(n_1515),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1475),
.B(n_1576),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1477),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1494),
.A2(n_1480),
.B(n_1490),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1490),
.A2(n_1462),
.B(n_1510),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1478),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1578),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1588),
.A2(n_1596),
.B(n_1592),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1562),
.B(n_1517),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1459),
.B(n_1517),
.Y(n_1667)
);

AO21x2_ASAP7_75t_L g1668 ( 
.A1(n_1529),
.A2(n_1476),
.B(n_1513),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1559),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1558),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1536),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1514),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1558),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1550),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1558),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1481),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1492),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1574),
.A2(n_1590),
.B1(n_1594),
.B2(n_1599),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1558),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1558),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1486),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1489),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1464),
.B(n_1601),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1550),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1483),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1568),
.A2(n_1584),
.B1(n_1581),
.B2(n_1591),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1491),
.B(n_1511),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1537),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1537),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1570),
.B(n_1572),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1495),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1495),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1503),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1580),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1574),
.B(n_1594),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1586),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_SL g1697 ( 
.A1(n_1590),
.A2(n_1479),
.B1(n_1593),
.B2(n_1477),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1541),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1514),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1507),
.A2(n_1519),
.B1(n_1463),
.B2(n_1493),
.C(n_1470),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1533),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1525),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1501),
.B(n_1598),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1593),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1629),
.A2(n_1522),
.B1(n_1469),
.B2(n_1501),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1603),
.B(n_1587),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1696),
.B(n_1587),
.Y(n_1707)
);

NAND4xp25_ASAP7_75t_L g1708 ( 
.A(n_1612),
.B(n_1606),
.C(n_1648),
.D(n_1667),
.Y(n_1708)
);

AO32x2_ASAP7_75t_L g1709 ( 
.A1(n_1622),
.A2(n_1516),
.A3(n_1484),
.B1(n_1473),
.B2(n_1467),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1632),
.B(n_1579),
.Y(n_1710)
);

O2A1O1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1667),
.A2(n_1598),
.B(n_1484),
.C(n_1522),
.Y(n_1711)
);

OAI211xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1639),
.A2(n_1516),
.B(n_1575),
.C(n_1502),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1662),
.A2(n_1620),
.B(n_1623),
.C(n_1661),
.Y(n_1713)
);

CKINVDCx20_ASAP7_75t_R g1714 ( 
.A(n_1614),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1626),
.B(n_1663),
.Y(n_1715)
);

NAND4xp25_ASAP7_75t_L g1716 ( 
.A(n_1684),
.B(n_1493),
.C(n_1501),
.D(n_1506),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1636),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1620),
.A2(n_1506),
.B1(n_1623),
.B2(n_1695),
.C(n_1678),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1695),
.A2(n_1686),
.B1(n_1666),
.B2(n_1683),
.C(n_1658),
.Y(n_1719)
);

AO21x2_ASAP7_75t_L g1720 ( 
.A1(n_1657),
.A2(n_1661),
.B(n_1652),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1683),
.A2(n_1641),
.B1(n_1697),
.B2(n_1666),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1626),
.B(n_1636),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_SL g1723 ( 
.A1(n_1684),
.A2(n_1669),
.B(n_1674),
.C(n_1700),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1724)
);

OAI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1641),
.A2(n_1659),
.B1(n_1671),
.B2(n_1658),
.C(n_1605),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1677),
.Y(n_1726)
);

OAI21xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1655),
.A2(n_1662),
.B(n_1674),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1633),
.A2(n_1655),
.B(n_1605),
.Y(n_1728)
);

BUFx12f_ASAP7_75t_L g1729 ( 
.A(n_1614),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1637),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1624),
.B(n_1628),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1628),
.B(n_1640),
.Y(n_1732)
);

CKINVDCx20_ASAP7_75t_R g1733 ( 
.A(n_1613),
.Y(n_1733)
);

AND2x6_ASAP7_75t_L g1734 ( 
.A(n_1687),
.B(n_1631),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_SL g1735 ( 
.A1(n_1669),
.A2(n_1674),
.B(n_1672),
.C(n_1693),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1640),
.B(n_1664),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1633),
.A2(n_1608),
.B(n_1605),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1699),
.B(n_1698),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1670),
.A2(n_1675),
.B(n_1679),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1609),
.B(n_1627),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1696),
.B(n_1682),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1664),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1610),
.B(n_1611),
.C(n_1694),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1656),
.A2(n_1690),
.B(n_1618),
.C(n_1652),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1610),
.B(n_1611),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1618),
.A2(n_1642),
.B(n_1669),
.C(n_1651),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1675),
.A2(n_1679),
.B(n_1608),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1618),
.B(n_1672),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1670),
.A2(n_1634),
.B(n_1680),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1691),
.B(n_1692),
.Y(n_1751)
);

A2O1A1Ixp33_ASAP7_75t_L g1752 ( 
.A1(n_1642),
.A2(n_1651),
.B(n_1681),
.C(n_1649),
.Y(n_1752)
);

O2A1O1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1644),
.A2(n_1634),
.B(n_1702),
.C(n_1701),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1616),
.A2(n_1617),
.B1(n_1681),
.B2(n_1703),
.C(n_1604),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1616),
.A2(n_1617),
.B(n_1604),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1613),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1665),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1644),
.A2(n_1634),
.B1(n_1685),
.B2(n_1668),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1647),
.A2(n_1649),
.B(n_1685),
.C(n_1643),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1665),
.B(n_1644),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1660),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1621),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1619),
.B(n_1615),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1673),
.A2(n_1680),
.B(n_1653),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1621),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1615),
.B(n_1694),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1751),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1765),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1731),
.B(n_1635),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1707),
.B(n_1712),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1763),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1765),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1732),
.B(n_1650),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1749),
.B(n_1646),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1763),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1715),
.B(n_1673),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1739),
.B(n_1635),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1724),
.B(n_1737),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1717),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1730),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1736),
.B(n_1627),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1762),
.B(n_1635),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1762),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1722),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1726),
.B(n_1630),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_1734),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1766),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1746),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1764),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1743),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1744),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1755),
.B(n_1688),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1734),
.B(n_1638),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1755),
.B(n_1630),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1757),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1706),
.B(n_1689),
.Y(n_1796)
);

NOR2xp67_ASAP7_75t_L g1797 ( 
.A(n_1750),
.B(n_1704),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1719),
.A2(n_1668),
.B1(n_1647),
.B2(n_1654),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1760),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1738),
.B(n_1625),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1713),
.B(n_1689),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1745),
.B(n_1653),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1760),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1798),
.A2(n_1708),
.B1(n_1719),
.B2(n_1718),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1769),
.B(n_1725),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1769),
.B(n_1725),
.Y(n_1806)
);

NAND2xp33_ASAP7_75t_L g1807 ( 
.A(n_1791),
.B(n_1756),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1786),
.B(n_1734),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1789),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1785),
.B(n_1738),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1771),
.B(n_1753),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1772),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1801),
.A2(n_1718),
.B1(n_1721),
.B2(n_1705),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1795),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1785),
.B(n_1728),
.Y(n_1815)
);

NAND4xp25_ASAP7_75t_L g1816 ( 
.A(n_1770),
.B(n_1728),
.C(n_1783),
.D(n_1742),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1771),
.B(n_1753),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1795),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1775),
.B(n_1727),
.Y(n_1819)
);

NOR3xp33_ASAP7_75t_L g1820 ( 
.A(n_1794),
.B(n_1705),
.C(n_1721),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1773),
.B(n_1748),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1778),
.B(n_1758),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1779),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1773),
.B(n_1748),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1779),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1794),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1788),
.B(n_1740),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1776),
.B(n_1740),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1802),
.A2(n_1758),
.B1(n_1754),
.B2(n_1720),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1768),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1793),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1788),
.B(n_1759),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1780),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1768),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1796),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1793),
.Y(n_1836)
);

INVx5_ASAP7_75t_L g1837 ( 
.A(n_1781),
.Y(n_1837)
);

AOI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1782),
.A2(n_1723),
.B1(n_1711),
.B2(n_1752),
.C(n_1747),
.Y(n_1838)
);

NOR3xp33_ASAP7_75t_L g1839 ( 
.A(n_1792),
.B(n_1712),
.C(n_1702),
.Y(n_1839)
);

AO21x2_ASAP7_75t_L g1840 ( 
.A1(n_1799),
.A2(n_1657),
.B(n_1654),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1777),
.B(n_1709),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1828),
.B(n_1783),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1828),
.B(n_1767),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1808),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1814),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1814),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1828),
.B(n_1821),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1837),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1840),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1827),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1827),
.B(n_1787),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1811),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1821),
.B(n_1767),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1840),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1818),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1818),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1822),
.B(n_1784),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1822),
.B(n_1784),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1823),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1819),
.B(n_1787),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1840),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1823),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1837),
.B(n_1797),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1825),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1811),
.B(n_1790),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1837),
.B(n_1793),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1825),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1833),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1808),
.Y(n_1869)
);

OAI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1816),
.A2(n_1735),
.B(n_1802),
.C(n_1711),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1833),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1819),
.B(n_1803),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1837),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1840),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1824),
.B(n_1800),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1817),
.B(n_1790),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1824),
.B(n_1800),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1809),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1841),
.B(n_1774),
.Y(n_1879)
);

NAND2x1p5_ASAP7_75t_L g1880 ( 
.A(n_1837),
.B(n_1741),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1845),
.Y(n_1881)
);

AND2x4_ASAP7_75t_SL g1882 ( 
.A(n_1844),
.B(n_1808),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1845),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1846),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1846),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1860),
.B(n_1817),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1855),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_L g1888 ( 
.A(n_1852),
.B(n_1816),
.C(n_1820),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1880),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1869),
.B(n_1837),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1869),
.B(n_1831),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1855),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1878),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1852),
.B(n_1841),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1850),
.B(n_1832),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1856),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_SL g1897 ( 
.A(n_1880),
.B(n_1733),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1843),
.B(n_1831),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1856),
.Y(n_1899)
);

NOR5xp2_ASAP7_75t_L g1900 ( 
.A(n_1870),
.B(n_1850),
.C(n_1812),
.D(n_1848),
.E(n_1873),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1880),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1865),
.B(n_1832),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1865),
.B(n_1810),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1859),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1859),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1860),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1862),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1862),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1876),
.B(n_1810),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1864),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1860),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1864),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1867),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1878),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1872),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1872),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1872),
.B(n_1834),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1876),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1878),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1843),
.B(n_1831),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1867),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1868),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1843),
.B(n_1831),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1868),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1880),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1871),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1921),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1886),
.B(n_1851),
.Y(n_1928)
);

OR2x6_ASAP7_75t_L g1929 ( 
.A(n_1888),
.B(n_1848),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1882),
.B(n_1847),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1895),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1882),
.B(n_1844),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1882),
.B(n_1847),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1893),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1902),
.B(n_1810),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1890),
.B(n_1847),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1906),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1926),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1890),
.B(n_1844),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1881),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1890),
.B(n_1844),
.Y(n_1941)
);

NAND2x1p5_ASAP7_75t_L g1942 ( 
.A(n_1890),
.B(n_1837),
.Y(n_1942)
);

NAND2x1_ASAP7_75t_SL g1943 ( 
.A(n_1911),
.B(n_1863),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1888),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1881),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1891),
.B(n_1842),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1883),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1886),
.B(n_1842),
.Y(n_1948)
);

NOR3xp33_ASAP7_75t_L g1949 ( 
.A(n_1918),
.B(n_1870),
.C(n_1820),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1893),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1891),
.B(n_1842),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1883),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1897),
.B(n_1875),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1901),
.B(n_1848),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1884),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1915),
.B(n_1916),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1903),
.B(n_1879),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1884),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1894),
.B(n_1851),
.Y(n_1959)
);

NOR2x1_ASAP7_75t_L g1960 ( 
.A(n_1901),
.B(n_1807),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1885),
.Y(n_1961)
);

AOI221xp5_ASAP7_75t_L g1962 ( 
.A1(n_1909),
.A2(n_1815),
.B1(n_1854),
.B2(n_1861),
.C(n_1874),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1885),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1949),
.B(n_1917),
.Y(n_1964)
);

O2A1O1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1944),
.A2(n_1900),
.B(n_1917),
.C(n_1839),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1929),
.A2(n_1813),
.B1(n_1804),
.B2(n_1953),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1953),
.B(n_1898),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1931),
.B(n_1879),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1940),
.Y(n_1969)
);

INVx1_ASAP7_75t_SL g1970 ( 
.A(n_1943),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1940),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1958),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1930),
.B(n_1901),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1937),
.Y(n_1974)
);

AOI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1929),
.A2(n_1813),
.B1(n_1804),
.B2(n_1806),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1956),
.B(n_1879),
.Y(n_1976)
);

OAI211xp5_ASAP7_75t_L g1977 ( 
.A1(n_1943),
.A2(n_1925),
.B(n_1889),
.C(n_1839),
.Y(n_1977)
);

INVxp67_ASAP7_75t_SL g1978 ( 
.A(n_1960),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1958),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1928),
.B(n_1887),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1936),
.B(n_1898),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1961),
.Y(n_1982)
);

OAI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1929),
.A2(n_1962),
.B(n_1935),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1961),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1963),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1936),
.B(n_1920),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1929),
.A2(n_1873),
.B(n_1866),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1930),
.Y(n_1988)
);

NAND2xp33_ASAP7_75t_L g1989 ( 
.A(n_1927),
.B(n_1714),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1933),
.A2(n_1806),
.B1(n_1805),
.B2(n_1829),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1933),
.Y(n_1991)
);

AOI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1965),
.A2(n_1938),
.B1(n_1927),
.B2(n_1963),
.C(n_1959),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1978),
.A2(n_1948),
.B(n_1938),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1975),
.B(n_1966),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1964),
.B(n_1968),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1976),
.B(n_1928),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1988),
.B(n_1946),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1970),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1974),
.B(n_1957),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1967),
.Y(n_2000)
);

AOI221xp5_ASAP7_75t_L g2001 ( 
.A1(n_1983),
.A2(n_1959),
.B1(n_1955),
.B2(n_1945),
.C(n_1952),
.Y(n_2001)
);

OAI32xp33_ASAP7_75t_L g2002 ( 
.A1(n_1988),
.A2(n_1942),
.A3(n_1889),
.B1(n_1925),
.B2(n_1951),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1991),
.B(n_1947),
.Y(n_2003)
);

AOI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_1990),
.A2(n_1861),
.B1(n_1874),
.B2(n_1854),
.C(n_1849),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1989),
.B(n_1729),
.Y(n_2005)
);

INVx1_ASAP7_75t_SL g2006 ( 
.A(n_1989),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1991),
.B(n_1946),
.Y(n_2007)
);

OAI322xp33_ASAP7_75t_L g2008 ( 
.A1(n_1980),
.A2(n_1942),
.A3(n_1934),
.B1(n_1950),
.B2(n_1904),
.C1(n_1908),
.C2(n_1899),
.Y(n_2008)
);

O2A1O1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1977),
.A2(n_1950),
.B(n_1934),
.C(n_1942),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1969),
.Y(n_2010)
);

AOI221xp5_ASAP7_75t_L g2011 ( 
.A1(n_1971),
.A2(n_1972),
.B1(n_1979),
.B2(n_1985),
.C(n_1984),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1982),
.Y(n_2012)
);

OAI21xp5_ASAP7_75t_SL g2013 ( 
.A1(n_1967),
.A2(n_1932),
.B(n_1954),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_R g2014 ( 
.A(n_2006),
.B(n_1710),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2000),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_2003),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1997),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_2008),
.A2(n_1987),
.B(n_1973),
.Y(n_2018)
);

NAND4xp75_ASAP7_75t_L g2019 ( 
.A(n_1992),
.B(n_1994),
.C(n_2001),
.D(n_1993),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1998),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_2009),
.B(n_1973),
.Y(n_2021)
);

XNOR2x2_ASAP7_75t_L g2022 ( 
.A(n_2011),
.B(n_1980),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2007),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1995),
.A2(n_1973),
.B1(n_1981),
.B2(n_1986),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1996),
.B(n_1981),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_2013),
.A2(n_1986),
.B1(n_1954),
.B2(n_1815),
.Y(n_2026)
);

OAI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_2004),
.A2(n_1805),
.B1(n_1861),
.B2(n_1874),
.C(n_1854),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_2020),
.B(n_1999),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2024),
.B(n_2005),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_2022),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_2024),
.B(n_2008),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2025),
.Y(n_2032)
);

NAND4xp75_ASAP7_75t_L g2033 ( 
.A(n_2021),
.B(n_2012),
.C(n_2010),
.D(n_1939),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_2025),
.B(n_2016),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_2019),
.B(n_2002),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2018),
.A2(n_2015),
.B(n_2027),
.Y(n_2036)
);

AOI211xp5_ASAP7_75t_L g2037 ( 
.A1(n_2017),
.A2(n_2023),
.B(n_2014),
.C(n_2026),
.Y(n_2037)
);

NOR3xp33_ASAP7_75t_L g2038 ( 
.A(n_2020),
.B(n_1954),
.C(n_1925),
.Y(n_2038)
);

NAND3xp33_ASAP7_75t_SL g2039 ( 
.A(n_2018),
.B(n_1951),
.C(n_1941),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2020),
.B(n_1932),
.Y(n_2040)
);

OAI21xp33_ASAP7_75t_L g2041 ( 
.A1(n_2030),
.A2(n_1941),
.B(n_1939),
.Y(n_2041)
);

AOI211xp5_ASAP7_75t_SL g2042 ( 
.A1(n_2031),
.A2(n_1932),
.B(n_1925),
.C(n_1889),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2040),
.B(n_2029),
.Y(n_2043)
);

NAND3xp33_ASAP7_75t_SL g2044 ( 
.A(n_2035),
.B(n_1838),
.C(n_1761),
.Y(n_2044)
);

AOI221xp5_ASAP7_75t_L g2045 ( 
.A1(n_2036),
.A2(n_1849),
.B1(n_1914),
.B2(n_1919),
.C(n_1896),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_2033),
.A2(n_1889),
.B(n_1873),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_2028),
.B(n_1887),
.Y(n_2047)
);

OAI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_2039),
.A2(n_1849),
.B1(n_1914),
.B2(n_1919),
.C(n_1829),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2043),
.B(n_2032),
.Y(n_2049)
);

AOI221xp5_ASAP7_75t_L g2050 ( 
.A1(n_2045),
.A2(n_2048),
.B1(n_2047),
.B2(n_2041),
.C(n_2034),
.Y(n_2050)
);

AOI322xp5_ASAP7_75t_L g2051 ( 
.A1(n_2044),
.A2(n_2038),
.A3(n_2037),
.B1(n_1815),
.B2(n_1875),
.C1(n_1877),
.C2(n_1826),
.Y(n_2051)
);

INVx1_ASAP7_75t_SL g2052 ( 
.A(n_2046),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_2042),
.B(n_2037),
.C(n_1838),
.Y(n_2053)
);

NOR3xp33_ASAP7_75t_L g2054 ( 
.A(n_2043),
.B(n_1709),
.C(n_1863),
.Y(n_2054)
);

OAI211xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2042),
.A2(n_1924),
.B(n_1892),
.C(n_1922),
.Y(n_2055)
);

NOR4xp25_ASAP7_75t_L g2056 ( 
.A(n_2043),
.B(n_1924),
.C(n_1892),
.D(n_1922),
.Y(n_2056)
);

NOR2x1_ASAP7_75t_L g2057 ( 
.A(n_2049),
.B(n_1896),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_2052),
.B(n_1920),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_2053),
.B(n_1923),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2056),
.B(n_1899),
.Y(n_2060)
);

NAND4xp75_ASAP7_75t_L g2061 ( 
.A(n_2050),
.B(n_1709),
.C(n_1923),
.D(n_1912),
.Y(n_2061)
);

NAND4xp75_ASAP7_75t_L g2062 ( 
.A(n_2051),
.B(n_1912),
.C(n_1910),
.D(n_1908),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_L g2063 ( 
.A(n_2057),
.B(n_2061),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2059),
.B(n_2054),
.Y(n_2064)
);

AOI221xp5_ASAP7_75t_SL g2065 ( 
.A1(n_2060),
.A2(n_2055),
.B1(n_1913),
.B2(n_1910),
.C(n_1907),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_2063),
.B(n_2058),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2066),
.Y(n_2067)
);

OAI21xp33_ASAP7_75t_L g2068 ( 
.A1(n_2067),
.A2(n_2064),
.B(n_2062),
.Y(n_2068)
);

AOI21xp33_ASAP7_75t_L g2069 ( 
.A1(n_2067),
.A2(n_2065),
.B(n_1905),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2068),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2069),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_1905),
.B(n_1904),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2070),
.A2(n_1913),
.B1(n_1907),
.B2(n_1877),
.Y(n_2073)
);

NAND3xp33_ASAP7_75t_L g2074 ( 
.A(n_2072),
.B(n_1858),
.C(n_1857),
.Y(n_2074)
);

AOI211xp5_ASAP7_75t_SL g2075 ( 
.A1(n_2074),
.A2(n_2073),
.B(n_1863),
.C(n_1836),
.Y(n_2075)
);

OAI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_2075),
.A2(n_1877),
.B1(n_1875),
.B2(n_1858),
.Y(n_2076)
);

OAI221xp5_ASAP7_75t_R g2077 ( 
.A1(n_2076),
.A2(n_1834),
.B1(n_1830),
.B2(n_1835),
.C(n_1853),
.Y(n_2077)
);

AOI211xp5_ASAP7_75t_L g2078 ( 
.A1(n_2077),
.A2(n_1863),
.B(n_1716),
.C(n_1857),
.Y(n_2078)
);


endmodule