module real_jpeg_12538_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_3),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_52),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_5),
.B(n_30),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_5),
.B(n_44),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_61),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_5),
.B(n_26),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_6),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_6),
.B(n_44),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_6),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_6),
.B(n_26),
.Y(n_105)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_6),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_6),
.B(n_50),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_8),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_8),
.B(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_8),
.B(n_61),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_8),
.B(n_50),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_8),
.B(n_52),
.Y(n_280)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_9),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_9),
.B(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_9),
.B(n_61),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_9),
.B(n_71),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_9),
.B(n_50),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_10),
.B(n_26),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_10),
.B(n_52),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_10),
.B(n_30),
.Y(n_147)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_13),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_13),
.B(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_13),
.B(n_44),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_13),
.B(n_61),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_13),
.B(n_26),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_13),
.B(n_71),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_13),
.B(n_50),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_13),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_14),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_14),
.Y(n_120)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_167),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_165),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_19),
.B(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_83),
.C(n_98),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_20),
.B(n_83),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_63),
.B2(n_64),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_21),
.B(n_65),
.C(n_76),
.Y(n_164)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_23),
.B(n_40),
.C(n_57),
.Y(n_132)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_25),
.B(n_29),
.C(n_32),
.Y(n_163)
);

INVx5_ASAP7_75t_SL g185 ( 
.A(n_26),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_33),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_33),
.B(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_36),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_36),
.B(n_119),
.Y(n_256)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_55),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_43),
.B(n_51),
.C(n_53),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_44),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_47),
.A2(n_53),
.B1(n_105),
.B2(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_49),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_49),
.B(n_107),
.Y(n_288)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_67),
.C(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_51),
.A2(n_54),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_51),
.B(n_258),
.Y(n_268)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_105),
.C(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_60),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_62),
.B(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_76),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_74),
.C(n_75),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_69),
.A2(n_70),
.B1(n_179),
.B2(n_180),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_70),
.B(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_72),
.B(n_123),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_72),
.B(n_107),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_75),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_77),
.B(n_79),
.C(n_81),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_80),
.A2(n_81),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_80),
.A2(n_81),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_80),
.A2(n_81),
.B1(n_95),
.B2(n_115),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_81),
.B(n_95),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.C(n_93),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_84),
.B(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_88),
.B(n_93),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.C(n_92),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_91),
.A2(n_157),
.B1(n_158),
.B2(n_161),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_91),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_91),
.A2(n_161),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_92),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.C(n_96),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_98),
.B(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_112),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_103),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_110),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_104),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_106),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_122),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_112),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_124),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_113),
.B(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_116),
.A2(n_117),
.B1(n_124),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_117),
.A2(n_118),
.B(n_121),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_119),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_123),
.B(n_185),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_124),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.C(n_127),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_125),
.B(n_126),
.CI(n_127),
.CON(n_177),
.SN(n_177)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_164),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_142),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_153),
.B2(n_154),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_147),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_162),
.B2(n_163),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_159),
.A2(n_160),
.B1(n_182),
.B2(n_183),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_182),
.C(n_184),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_195),
.B(n_326),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_193),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_169),
.B(n_193),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_172),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_186),
.C(n_189),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_181),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_176),
.A2(n_177),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_177),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_178),
.B(n_181),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_184),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_243),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_220),
.B(n_242),
.Y(n_197)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_198),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_218),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.C(n_206),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.C(n_217),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_207),
.B(n_210),
.CI(n_217),
.CON(n_226),
.SN(n_226)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_211),
.A2(n_212),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_221),
.B(n_224),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.C(n_231),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_225),
.A2(n_226),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_226),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_227),
.A2(n_228),
.B1(n_231),
.B2(n_232),
.Y(n_322)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.C(n_236),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_233),
.B(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_236),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.C(n_240),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_324),
.C(n_325),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_318),
.B(n_323),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_303),
.B(n_317),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_273),
.B(n_302),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_260),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_248),
.B(n_260),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.C(n_257),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_249),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_249),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_299),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.CI(n_252),
.CON(n_249),
.SN(n_249)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_300),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_267),
.B2(n_272),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_266),
.C(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_270),
.C(n_271),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_296),
.B(n_301),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_286),
.B(n_295),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_276),
.B(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_290),
.B(n_294),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_289),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_305),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_311),
.C(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_315),
.B2(n_316),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);


endmodule