module fake_jpeg_17002_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_27),
.C(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_40),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_29),
.B1(n_27),
.B2(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_35),
.B1(n_20),
.B2(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_58),
.B1(n_64),
.B2(n_21),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_35),
.B1(n_20),
.B2(n_24),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_30),
.B1(n_28),
.B2(n_26),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_30),
.B1(n_28),
.B2(n_26),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_67),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_31),
.B1(n_21),
.B2(n_34),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_87),
.B1(n_99),
.B2(n_100),
.Y(n_114)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_76),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_37),
.B(n_43),
.C(n_34),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_89),
.B(n_22),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_37),
.B(n_39),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_22),
.B(n_38),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_74),
.A2(n_82),
.B(n_93),
.Y(n_126)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_86),
.Y(n_127)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_27),
.B1(n_40),
.B2(n_18),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_38),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_38),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_39),
.B(n_32),
.C(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_25),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_50),
.B(n_25),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_42),
.C(n_17),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_102),
.Y(n_123)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_47),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_104),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_46),
.A2(n_39),
.B1(n_17),
.B2(n_32),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_38),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_98),
.C(n_65),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_9),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_120),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_86),
.B1(n_77),
.B2(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_38),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_0),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_73),
.B(n_1),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_9),
.B(n_12),
.C(n_16),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_71),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_138),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_154),
.B(n_117),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_143),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_118),
.B(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_72),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_150),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_74),
.C(n_78),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_152),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_74),
.B1(n_73),
.B2(n_96),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_162),
.B1(n_114),
.B2(n_14),
.Y(n_173)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_75),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_99),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_153),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_42),
.C(n_95),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_122),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_76),
.B1(n_81),
.B2(n_87),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_161),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_68),
.B1(n_85),
.B2(n_80),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_100),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_159),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_0),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_128),
.B1(n_127),
.B2(n_126),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_111),
.B(n_107),
.C(n_123),
.D(n_118),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_169),
.B(n_180),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_164),
.B(n_186),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_174),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_121),
.B(n_110),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_110),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_183),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_158),
.B(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_105),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_105),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_121),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_121),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_117),
.B(n_119),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_131),
.B(n_129),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_22),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_210),
.B1(n_211),
.B2(n_192),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_135),
.B1(n_146),
.B2(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_198),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_152),
.B1(n_136),
.B2(n_140),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_191),
.A2(n_153),
.B1(n_144),
.B2(n_159),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_144),
.B1(n_142),
.B2(n_138),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_213),
.B1(n_167),
.B2(n_190),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_188),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_215),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_131),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_119),
.Y(n_214)
);

NOR4xp25_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_129),
.C(n_108),
.D(n_7),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_170),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_219),
.C(n_221),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_217),
.A2(n_213),
.B(n_200),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_170),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_178),
.B1(n_168),
.B2(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_171),
.C(n_172),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_187),
.B(n_178),
.C(n_164),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVxp33_ASAP7_75t_SL g225 ( 
.A(n_206),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_175),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_171),
.C(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_231),
.C(n_232),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_169),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_194),
.A2(n_186),
.B1(n_189),
.B2(n_176),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_202),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_193),
.C(n_197),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_251),
.C(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_242),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_195),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_231),
.C(n_222),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_204),
.C(n_197),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_254),
.C(n_255),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_232),
.C(n_228),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_222),
.C(n_234),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_257),
.C(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_249),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_212),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_252),
.C(n_254),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_267),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_163),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_247),
.C(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_259),
.B(n_204),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_1),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_269),
.A2(n_250),
.B1(n_263),
.B2(n_205),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_279),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_210),
.C(n_188),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_277),
.C(n_268),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_273),
.A2(n_213),
.B1(n_108),
.B2(n_7),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_1),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_283),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_SL g284 ( 
.A(n_275),
.B(n_266),
.Y(n_284)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_285),
.A3(n_276),
.B1(n_278),
.B2(n_277),
.C1(n_8),
.C2(n_5),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_6),
.CI(n_13),
.CON(n_285),
.SN(n_285)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_287),
.A3(n_10),
.B1(n_14),
.B2(n_3),
.C1(n_4),
.C2(n_1),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_5),
.B(n_10),
.Y(n_287)
);

A2O1A1O1Ixp25_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_281),
.B(n_285),
.C(n_6),
.D(n_10),
.Y(n_290)
);

AOI321xp33_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_291),
.A3(n_2),
.B1(n_3),
.B2(n_288),
.C(n_56),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_2),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_2),
.Y(n_294)
);


endmodule