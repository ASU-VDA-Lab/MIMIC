module fake_jpeg_12952_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_44),
.B(n_70),
.Y(n_102)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_3),
.C(n_4),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_62),
.Y(n_96)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_50),
.Y(n_107)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_3),
.CON(n_52),
.SN(n_52)
);

OR2x4_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_5),
.Y(n_85)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_67),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_20),
.B(n_12),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_68),
.Y(n_98)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_4),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_10),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_37),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_75),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_78),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_74),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_37),
.B(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_5),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_89),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_93),
.B1(n_113),
.B2(n_91),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_85),
.A2(n_91),
.B(n_106),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_47),
.B1(n_51),
.B2(n_72),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_110),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_29),
.B1(n_31),
.B2(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_31),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_55),
.A2(n_25),
.B1(n_29),
.B2(n_19),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_43),
.B1(n_73),
.B2(n_58),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_26),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_124),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_76),
.A2(n_26),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_118),
.A2(n_108),
.B1(n_95),
.B2(n_92),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_45),
.B(n_6),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_112),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_43),
.A2(n_9),
.B1(n_64),
.B2(n_56),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_121),
.B1(n_96),
.B2(n_118),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_126),
.A2(n_139),
.B(n_157),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_85),
.A2(n_79),
.B1(n_62),
.B2(n_9),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_9),
.B1(n_112),
.B2(n_115),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_121),
.A2(n_117),
.B1(n_109),
.B2(n_86),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_157),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_138),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_109),
.B1(n_86),
.B2(n_94),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_151),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_99),
.B(n_88),
.C(n_92),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_88),
.A2(n_84),
.B(n_116),
.C(n_103),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_126),
.Y(n_164)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_82),
.B(n_97),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_124),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_167),
.B(n_142),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_132),
.C(n_127),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_143),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_156),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_150),
.B(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_192),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_128),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_128),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_203),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_194),
.B(n_195),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_129),
.C(n_142),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_163),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_200),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_164),
.B(n_186),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_163),
.A2(n_131),
.B1(n_147),
.B2(n_136),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_201),
.Y(n_215)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_134),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_205),
.B(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_170),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_221),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_188),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_202),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_173),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_191),
.C(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_182),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_177),
.B1(n_184),
.B2(n_180),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_200),
.B1(n_198),
.B2(n_204),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_229),
.Y(n_240)
);

OAI322xp33_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_197),
.A3(n_191),
.B1(n_196),
.B2(n_203),
.C1(n_207),
.C2(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_231),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_233),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_179),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_179),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_236),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_225),
.B(n_209),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_238),
.Y(n_253)
);

A2O1A1O1Ixp25_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_213),
.B(n_222),
.C(n_218),
.D(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_214),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_213),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_235),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_240),
.A2(n_235),
.B(n_231),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_224),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_255),
.C(n_246),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_254),
.B(n_241),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_253),
.B1(n_239),
.B2(n_215),
.Y(n_257)
);

OAI322xp33_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_210),
.A3(n_237),
.B1(n_220),
.B2(n_223),
.C1(n_215),
.C2(n_183),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_165),
.C(n_174),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_242),
.B1(n_244),
.B2(n_249),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_259),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_260),
.B(n_172),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_165),
.B(n_180),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_257),
.A2(n_250),
.B(n_162),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_162),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_261),
.C(n_259),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_187),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_263),
.B(n_172),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_270),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_174),
.Y(n_273)
);


endmodule