module real_aes_6900_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_727, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_727;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g469 ( .A1(n_0), .A2(n_207), .B(n_470), .C(n_473), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_1), .B(n_464), .Y(n_474) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g242 ( .A(n_3), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_4), .B(n_159), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_5), .A2(n_459), .B(n_547), .Y(n_546) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_6), .A2(n_182), .B(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_7), .A2(n_39), .B1(n_152), .B2(n_176), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_8), .A2(n_105), .B1(n_118), .B2(n_725), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_9), .B(n_182), .Y(n_254) );
AND2x6_ASAP7_75t_L g167 ( .A(n_10), .B(n_168), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_11), .A2(n_167), .B(n_450), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_12), .B(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_12), .B(n_40), .Y(n_128) );
INVx1_ASAP7_75t_L g148 ( .A(n_13), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_14), .B(n_157), .Y(n_190) );
INVx1_ASAP7_75t_L g234 ( .A(n_15), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_16), .A2(n_76), .B1(n_718), .B2(n_719), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_16), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_17), .B(n_159), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_18), .B(n_183), .Y(n_221) );
AO32x2_ASAP7_75t_L g204 ( .A1(n_19), .A2(n_181), .A3(n_182), .B1(n_205), .B2(n_209), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_20), .B(n_152), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_21), .B(n_183), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_22), .A2(n_56), .B1(n_152), .B2(n_176), .Y(n_208) );
AOI22xp33_ASAP7_75t_SL g179 ( .A1(n_23), .A2(n_83), .B1(n_152), .B2(n_157), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_24), .B(n_152), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_25), .A2(n_181), .B(n_450), .C(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_26), .A2(n_181), .B(n_450), .C(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_27), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_28), .B(n_144), .Y(n_263) );
OAI22xp5_ASAP7_75t_SL g704 ( .A1(n_29), .A2(n_94), .B1(n_705), .B2(n_706), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_29), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_30), .A2(n_703), .B1(n_704), .B2(n_707), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_30), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_31), .A2(n_459), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_32), .B(n_144), .Y(n_169) );
INVx2_ASAP7_75t_L g154 ( .A(n_33), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_34), .A2(n_456), .B(n_482), .C(n_483), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_35), .B(n_152), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_36), .B(n_144), .Y(n_197) );
OAI22xp5_ASAP7_75t_SL g722 ( .A1(n_37), .A2(n_44), .B1(n_440), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_37), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_38), .B(n_192), .Y(n_513) );
INVx1_ASAP7_75t_L g117 ( .A(n_40), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_41), .B(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_42), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_43), .B(n_159), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_44), .A2(n_135), .B1(n_440), .B2(n_441), .Y(n_134) );
INVx1_ASAP7_75t_L g440 ( .A(n_44), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_45), .B(n_459), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_46), .A2(n_456), .B(n_482), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_47), .B(n_152), .Y(n_249) );
INVx1_ASAP7_75t_L g471 ( .A(n_48), .Y(n_471) );
AOI22xp5_ASAP7_75t_SL g130 ( .A1(n_49), .A2(n_126), .B1(n_131), .B2(n_710), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_50), .A2(n_92), .B1(n_176), .B2(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g534 ( .A(n_51), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_52), .B(n_152), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_53), .B(n_152), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_54), .B(n_459), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_55), .B(n_240), .Y(n_253) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_57), .A2(n_61), .B1(n_152), .B2(n_157), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_58), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_59), .B(n_152), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_60), .B(n_152), .Y(n_262) );
INVx1_ASAP7_75t_L g168 ( .A(n_62), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_63), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_64), .B(n_464), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_65), .A2(n_237), .B(n_240), .C(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_66), .B(n_152), .Y(n_243) );
INVx1_ASAP7_75t_L g147 ( .A(n_67), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_68), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_69), .B(n_159), .Y(n_487) );
AO32x2_ASAP7_75t_L g173 ( .A1(n_70), .A2(n_174), .A3(n_180), .B1(n_181), .B2(n_182), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_71), .B(n_160), .Y(n_524) );
INVx1_ASAP7_75t_L g261 ( .A(n_72), .Y(n_261) );
INVx1_ASAP7_75t_L g155 ( .A(n_73), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_74), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_75), .B(n_486), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_76), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_77), .A2(n_450), .B(n_452), .C(n_456), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_78), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_79), .B(n_157), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_80), .Y(n_548) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_82), .B(n_485), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_84), .B(n_176), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_85), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_86), .B(n_157), .Y(n_164) );
INVx2_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_88), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_89), .B(n_178), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_90), .B(n_157), .Y(n_250) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_91), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g125 ( .A(n_91), .B(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_93), .A2(n_103), .B1(n_157), .B2(n_158), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_94), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_95), .B(n_459), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_96), .Y(n_484) );
INVxp67_ASAP7_75t_L g551 ( .A(n_97), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_98), .B(n_157), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g453 ( .A(n_100), .Y(n_453) );
INVx1_ASAP7_75t_L g520 ( .A(n_101), .Y(n_520) );
AND2x2_ASAP7_75t_L g536 ( .A(n_102), .B(n_144), .Y(n_536) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g725 ( .A(n_108), .Y(n_725) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_115), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g127 ( .A(n_111), .B(n_128), .Y(n_127) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_130), .B1(n_713), .B2(n_714), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g713 ( .A(n_121), .Y(n_713) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_123), .A2(n_715), .B(n_724), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_129), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g724 ( .A(n_125), .Y(n_724) );
NOR2x2_ASAP7_75t_L g712 ( .A(n_126), .B(n_133), .Y(n_712) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp33_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_702), .B1(n_708), .B2(n_709), .Y(n_131) );
INVx1_ASAP7_75t_L g708 ( .A(n_132), .Y(n_708) );
AO22x2_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_134), .B1(n_442), .B2(n_701), .Y(n_132) );
INVx1_ASAP7_75t_L g701 ( .A(n_133), .Y(n_701) );
INVx1_ASAP7_75t_L g441 ( .A(n_135), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_135), .A2(n_441), .B1(n_721), .B2(n_722), .Y(n_720) );
OR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_361), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_310), .C(n_352), .Y(n_136) );
AOI211xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_215), .B(n_264), .C(n_286), .Y(n_137) );
OAI211xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_170), .B(n_198), .C(n_210), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_140), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g373 ( .A(n_140), .B(n_290), .Y(n_373) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g275 ( .A(n_141), .B(n_201), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_141), .B(n_186), .Y(n_392) );
INVx1_ASAP7_75t_L g410 ( .A(n_141), .Y(n_410) );
AND2x2_ASAP7_75t_L g419 ( .A(n_141), .B(n_307), .Y(n_419) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g302 ( .A(n_142), .B(n_186), .Y(n_302) );
AND2x2_ASAP7_75t_L g360 ( .A(n_142), .B(n_307), .Y(n_360) );
INVx1_ASAP7_75t_L g404 ( .A(n_142), .Y(n_404) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g281 ( .A(n_143), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g289 ( .A(n_143), .Y(n_289) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_143), .Y(n_329) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_149), .B(n_169), .Y(n_143) );
INVx2_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_144), .A2(n_187), .B(n_197), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_144), .A2(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g503 ( .A(n_144), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_144), .A2(n_531), .B(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_L g183 ( .A(n_145), .B(n_146), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_162), .B(n_167), .Y(n_149) );
O2A1O1Ixp5_ASAP7_75t_SL g150 ( .A1(n_151), .A2(n_155), .B(n_156), .C(n_159), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_152), .Y(n_455) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
AND2x6_ASAP7_75t_L g450 ( .A(n_153), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g158 ( .A(n_154), .Y(n_158) );
INVx1_ASAP7_75t_L g241 ( .A(n_154), .Y(n_241) );
INVx2_ASAP7_75t_L g235 ( .A(n_157), .Y(n_235) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_159), .A2(n_249), .B(n_250), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_159), .A2(n_258), .B(n_259), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_159), .B(n_551), .Y(n_550) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g174 ( .A1(n_160), .A2(n_175), .B1(n_178), .B2(n_179), .Y(n_174) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_161), .Y(n_166) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
INVx1_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
INVx1_ASAP7_75t_L g451 ( .A(n_161), .Y(n_451) );
AND2x2_ASAP7_75t_L g460 ( .A(n_161), .B(n_241), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .Y(n_162) );
INVx1_ASAP7_75t_L g237 ( .A(n_165), .Y(n_237) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g486 ( .A(n_166), .Y(n_486) );
BUFx3_ASAP7_75t_L g181 ( .A(n_167), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_167), .A2(n_188), .B(n_193), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_167), .A2(n_233), .B(n_238), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_167), .A2(n_248), .B(n_251), .Y(n_247) );
INVx4_ASAP7_75t_SL g457 ( .A(n_167), .Y(n_457) );
AND2x4_ASAP7_75t_L g459 ( .A(n_167), .B(n_460), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_167), .B(n_460), .Y(n_521) );
INVxp67_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_184), .Y(n_171) );
AND2x2_ASAP7_75t_L g268 ( .A(n_172), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g301 ( .A(n_172), .Y(n_301) );
OR2x2_ASAP7_75t_L g427 ( .A(n_172), .B(n_428), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_172), .B(n_186), .Y(n_431) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
INVx1_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
AND2x2_ASAP7_75t_L g290 ( .A(n_173), .B(n_203), .Y(n_290) );
AND2x2_ASAP7_75t_L g330 ( .A(n_173), .B(n_204), .Y(n_330) );
INVx2_ASAP7_75t_L g473 ( .A(n_177), .Y(n_473) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_177), .Y(n_488) );
INVx2_ASAP7_75t_L g196 ( .A(n_178), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_178), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_178), .A2(n_207), .B1(n_224), .B2(n_225), .Y(n_223) );
INVx4_ASAP7_75t_L g472 ( .A(n_178), .Y(n_472) );
INVx1_ASAP7_75t_L g500 ( .A(n_180), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_181), .B(n_223), .C(n_226), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_181), .A2(n_257), .B(n_260), .Y(n_256) );
INVx4_ASAP7_75t_L g226 ( .A(n_182), .Y(n_226) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_182), .A2(n_247), .B(n_254), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_182), .A2(n_510), .B(n_511), .Y(n_509) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_182), .Y(n_545) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g209 ( .A(n_183), .Y(n_209) );
INVxp67_ASAP7_75t_L g372 ( .A(n_184), .Y(n_372) );
AND2x4_ASAP7_75t_L g397 ( .A(n_184), .B(n_290), .Y(n_397) );
BUFx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_SL g288 ( .A(n_185), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g202 ( .A(n_186), .B(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g276 ( .A(n_186), .B(n_204), .Y(n_276) );
INVx1_ASAP7_75t_L g282 ( .A(n_186), .Y(n_282) );
INVx2_ASAP7_75t_L g308 ( .A(n_186), .Y(n_308) );
AND2x2_ASAP7_75t_L g324 ( .A(n_186), .B(n_325), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .Y(n_193) );
O2A1O1Ixp5_ASAP7_75t_L g260 ( .A1(n_196), .A2(n_239), .B(n_261), .C(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_199), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_202), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g279 ( .A(n_201), .Y(n_279) );
AND2x2_ASAP7_75t_L g387 ( .A(n_201), .B(n_203), .Y(n_387) );
AND2x2_ASAP7_75t_L g304 ( .A(n_202), .B(n_289), .Y(n_304) );
AND2x2_ASAP7_75t_L g403 ( .A(n_202), .B(n_404), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g325 ( .A(n_203), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g428 ( .A(n_203), .B(n_289), .Y(n_428) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
BUFx2_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
AND2x2_ASAP7_75t_L g307 ( .A(n_204), .B(n_308), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_207), .A2(n_239), .B(n_242), .C(n_243), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_207), .A2(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g231 ( .A(n_209), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_209), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_214), .Y(n_211) );
AND2x2_ASAP7_75t_L g353 ( .A(n_212), .B(n_288), .Y(n_353) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_213), .B(n_289), .Y(n_338) );
INVx2_ASAP7_75t_L g337 ( .A(n_214), .Y(n_337) );
OAI222xp33_ASAP7_75t_L g341 ( .A1(n_214), .A2(n_281), .B1(n_342), .B2(n_344), .C1(n_345), .C2(n_348), .Y(n_341) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g266 ( .A(n_219), .Y(n_266) );
OR2x2_ASAP7_75t_L g377 ( .A(n_219), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx3_ASAP7_75t_L g299 ( .A(n_220), .Y(n_299) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_220), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g356 ( .A(n_220), .B(n_270), .Y(n_356) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g317 ( .A(n_221), .Y(n_317) );
AO21x1_ASAP7_75t_L g316 ( .A1(n_223), .A2(n_226), .B(n_317), .Y(n_316) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_226), .A2(n_448), .B(n_461), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_226), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g464 ( .A(n_226), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_226), .B(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_226), .A2(n_519), .B(n_526), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_227), .A2(n_320), .B1(n_359), .B2(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_245), .Y(n_227) );
INVx3_ASAP7_75t_L g292 ( .A(n_228), .Y(n_292) );
OR2x2_ASAP7_75t_L g425 ( .A(n_228), .B(n_301), .Y(n_425) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g298 ( .A(n_229), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g314 ( .A(n_229), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g322 ( .A(n_229), .B(n_270), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_229), .B(n_246), .Y(n_378) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g269 ( .A(n_230), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g273 ( .A(n_230), .B(n_246), .Y(n_273) );
AND2x2_ASAP7_75t_L g349 ( .A(n_230), .B(n_296), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_230), .B(n_255), .Y(n_389) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_244), .Y(n_230) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_231), .A2(n_256), .B(n_263), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .C(n_237), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_235), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_235), .A2(n_524), .B(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_237), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_239), .A2(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_245), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g305 ( .A(n_245), .B(n_266), .Y(n_305) );
AND2x2_ASAP7_75t_L g309 ( .A(n_245), .B(n_299), .Y(n_309) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
INVx3_ASAP7_75t_L g270 ( .A(n_246), .Y(n_270) );
AND2x2_ASAP7_75t_L g295 ( .A(n_246), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g430 ( .A(n_246), .B(n_413), .Y(n_430) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_255), .Y(n_284) );
INVx2_ASAP7_75t_L g296 ( .A(n_255), .Y(n_296) );
AND2x2_ASAP7_75t_L g340 ( .A(n_255), .B(n_316), .Y(n_340) );
INVx1_ASAP7_75t_L g383 ( .A(n_255), .Y(n_383) );
OR2x2_ASAP7_75t_L g414 ( .A(n_255), .B(n_316), .Y(n_414) );
AND2x2_ASAP7_75t_L g434 ( .A(n_255), .B(n_270), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B(n_271), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g272 ( .A(n_266), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_266), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g391 ( .A(n_268), .Y(n_391) );
INVx2_ASAP7_75t_SL g285 ( .A(n_269), .Y(n_285) );
AND2x2_ASAP7_75t_L g405 ( .A(n_269), .B(n_299), .Y(n_405) );
INVx2_ASAP7_75t_L g351 ( .A(n_270), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_270), .B(n_383), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B1(n_277), .B2(n_283), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_273), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g439 ( .A(n_273), .Y(n_439) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g364 ( .A(n_275), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_275), .B(n_307), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_276), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g380 ( .A(n_276), .B(n_329), .Y(n_380) );
INVx2_ASAP7_75t_L g436 ( .A(n_276), .Y(n_436) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g306 ( .A(n_279), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_279), .B(n_324), .Y(n_357) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_281), .B(n_301), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g418 ( .A(n_284), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_SL g368 ( .A1(n_285), .A2(n_369), .B(n_371), .C(n_374), .Y(n_368) );
OR2x2_ASAP7_75t_L g395 ( .A(n_285), .B(n_299), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_291), .B1(n_293), .B2(n_300), .C(n_303), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_288), .B(n_337), .Y(n_344) );
AND2x2_ASAP7_75t_L g386 ( .A(n_288), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g422 ( .A(n_288), .Y(n_422) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
INVx1_ASAP7_75t_L g326 ( .A(n_289), .Y(n_326) );
NOR2xp67_ASAP7_75t_L g346 ( .A(n_292), .B(n_347), .Y(n_346) );
INVxp67_ASAP7_75t_L g400 ( .A(n_292), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_292), .B(n_340), .Y(n_416) );
INVx2_ASAP7_75t_L g402 ( .A(n_293), .Y(n_402) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g343 ( .A(n_295), .B(n_314), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g352 ( .A1(n_295), .A2(n_311), .B(n_353), .C(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g321 ( .A(n_296), .B(n_316), .Y(n_321) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_300), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OR2x2_ASAP7_75t_L g369 ( .A(n_301), .B(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_306), .B2(n_309), .Y(n_303) );
INVx1_ASAP7_75t_L g423 ( .A(n_305), .Y(n_423) );
INVx1_ASAP7_75t_L g370 ( .A(n_307), .Y(n_370) );
INVx1_ASAP7_75t_L g421 ( .A(n_309), .Y(n_421) );
AOI211xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_314), .B(n_318), .C(n_341), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g333 ( .A(n_313), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g384 ( .A(n_314), .Y(n_384) );
AND2x2_ASAP7_75t_L g433 ( .A(n_314), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_323), .B(n_331), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx2_ASAP7_75t_L g347 ( .A(n_321), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_321), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g339 ( .A(n_322), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g415 ( .A(n_322), .Y(n_415) );
OAI32xp33_ASAP7_75t_L g426 ( .A1(n_322), .A2(n_374), .A3(n_381), .B1(n_422), .B2(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_SL g394 ( .A(n_324), .Y(n_394) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g334 ( .A(n_330), .Y(n_334) );
OAI21xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_333), .A2(n_381), .B1(n_407), .B2(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_337), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g367 ( .A(n_351), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_360), .A2(n_402), .B1(n_403), .B2(n_405), .C(n_406), .Y(n_401) );
NAND5xp2_ASAP7_75t_L g361 ( .A(n_362), .B(n_385), .C(n_401), .D(n_411), .E(n_429), .Y(n_361) );
AOI211xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_365), .B(n_368), .C(n_375), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g432 ( .A(n_369), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_379), .B2(n_381), .Y(n_375) );
INVx1_ASAP7_75t_SL g408 ( .A(n_378), .Y(n_408) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI322xp33_ASAP7_75t_L g390 ( .A1(n_381), .A2(n_391), .A3(n_392), .B1(n_393), .B2(n_394), .C1(n_395), .C2(n_396), .Y(n_390) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g393 ( .A(n_383), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_383), .B(n_408), .Y(n_407) );
AOI211xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_388), .B(n_390), .C(n_398), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_420) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_419), .B1(n_420), .B2(n_424), .C(n_426), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_415), .B(n_416), .C(n_417), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g438 ( .A(n_414), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B1(n_432), .B2(n_433), .C(n_435), .Y(n_429) );
AOI21xp33_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_437), .B(n_438), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_443), .B(n_644), .Y(n_442) );
AND4x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_584), .C(n_599), .D(n_624), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g444 ( .A(n_445), .B(n_557), .Y(n_444) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_475), .B(n_537), .Y(n_445) );
AND2x2_ASAP7_75t_L g587 ( .A(n_446), .B(n_492), .Y(n_587) );
AND2x2_ASAP7_75t_L g600 ( .A(n_446), .B(n_491), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_446), .B(n_476), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_446), .Y(n_654) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_463), .Y(n_446) );
INVx2_ASAP7_75t_L g571 ( .A(n_447), .Y(n_571) );
BUFx2_ASAP7_75t_L g598 ( .A(n_447), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_458), .Y(n_448) );
INVx5_ASAP7_75t_L g468 ( .A(n_450), .Y(n_468) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_SL g466 ( .A1(n_457), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_457), .A2(n_468), .B(n_548), .C(n_549), .Y(n_547) );
BUFx2_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
AND2x2_ASAP7_75t_L g538 ( .A(n_463), .B(n_492), .Y(n_538) );
INVx2_ASAP7_75t_L g554 ( .A(n_463), .Y(n_554) );
AND2x2_ASAP7_75t_L g563 ( .A(n_463), .B(n_491), .Y(n_563) );
AND2x2_ASAP7_75t_L g642 ( .A(n_463), .B(n_571), .Y(n_642) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_474), .Y(n_463) );
INVx2_ASAP7_75t_L g482 ( .A(n_468), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_504), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_476), .B(n_569), .Y(n_607) );
INVx1_ASAP7_75t_L g695 ( .A(n_476), .Y(n_695) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_491), .Y(n_476) );
AND2x2_ASAP7_75t_L g553 ( .A(n_477), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g567 ( .A(n_477), .B(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_477), .Y(n_596) );
OR2x2_ASAP7_75t_L g628 ( .A(n_477), .B(n_570), .Y(n_628) );
AND2x2_ASAP7_75t_L g636 ( .A(n_477), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g669 ( .A(n_477), .B(n_638), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_477), .B(n_538), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_477), .B(n_598), .Y(n_694) );
AND2x2_ASAP7_75t_L g700 ( .A(n_477), .B(n_587), .Y(n_700) );
INVx5_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g560 ( .A(n_478), .Y(n_560) );
AND2x2_ASAP7_75t_L g590 ( .A(n_478), .B(n_570), .Y(n_590) );
AND2x2_ASAP7_75t_L g623 ( .A(n_478), .B(n_583), .Y(n_623) );
AND2x2_ASAP7_75t_L g643 ( .A(n_478), .B(n_492), .Y(n_643) );
AND2x2_ASAP7_75t_L g677 ( .A(n_478), .B(n_543), .Y(n_677) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B(n_487), .C(n_488), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_485), .A2(n_488), .B(n_534), .C(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g583 ( .A(n_491), .B(n_554), .Y(n_583) );
AND2x2_ASAP7_75t_L g594 ( .A(n_491), .B(n_590), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_491), .B(n_570), .Y(n_633) );
INVx2_ASAP7_75t_L g648 ( .A(n_491), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_491), .B(n_582), .Y(n_671) );
AND2x2_ASAP7_75t_L g690 ( .A(n_491), .B(n_642), .Y(n_690) );
INVx5_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_492), .Y(n_589) );
AND2x2_ASAP7_75t_L g597 ( .A(n_492), .B(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g638 ( .A(n_492), .B(n_554), .Y(n_638) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
AOI21xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_496), .B(n_500), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
AND2x2_ASAP7_75t_L g561 ( .A(n_506), .B(n_544), .Y(n_561) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_507), .B(n_518), .Y(n_541) );
OR2x2_ASAP7_75t_L g574 ( .A(n_507), .B(n_544), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_507), .B(n_544), .Y(n_579) );
AND2x2_ASAP7_75t_L g606 ( .A(n_507), .B(n_543), .Y(n_606) );
AND2x2_ASAP7_75t_L g658 ( .A(n_507), .B(n_517), .Y(n_658) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_508), .B(n_528), .Y(n_566) );
AND2x2_ASAP7_75t_L g602 ( .A(n_508), .B(n_518), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_515), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g592 ( .A(n_516), .B(n_574), .Y(n_592) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_528), .Y(n_516) );
OAI322xp33_ASAP7_75t_L g557 ( .A1(n_517), .A2(n_558), .A3(n_562), .B1(n_564), .B2(n_567), .C1(n_572), .C2(n_580), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_517), .B(n_543), .Y(n_565) );
OR2x2_ASAP7_75t_L g575 ( .A(n_517), .B(n_529), .Y(n_575) );
AND2x2_ASAP7_75t_L g577 ( .A(n_517), .B(n_529), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_517), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_517), .B(n_544), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_517), .B(n_673), .Y(n_672) );
INVx5_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_518), .B(n_561), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_522), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_528), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g555 ( .A(n_528), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_528), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g617 ( .A(n_528), .B(n_544), .Y(n_617) );
AOI211xp5_ASAP7_75t_SL g645 ( .A1(n_528), .A2(n_646), .B(n_649), .C(n_661), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_528), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g683 ( .A(n_528), .B(n_658), .Y(n_683) );
INVx5_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g611 ( .A(n_529), .B(n_544), .Y(n_611) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_529), .Y(n_620) );
AND2x2_ASAP7_75t_L g660 ( .A(n_529), .B(n_658), .Y(n_660) );
AND2x2_ASAP7_75t_SL g691 ( .A(n_529), .B(n_561), .Y(n_691) );
AND2x2_ASAP7_75t_L g698 ( .A(n_529), .B(n_657), .Y(n_698) );
OR2x6_ASAP7_75t_L g529 ( .A(n_530), .B(n_536), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_553), .B2(n_555), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_538), .B(n_560), .Y(n_608) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g556 ( .A(n_541), .Y(n_556) );
OR2x2_ASAP7_75t_L g616 ( .A(n_541), .B(n_617), .Y(n_616) );
OAI221xp5_ASAP7_75t_SL g664 ( .A1(n_541), .A2(n_665), .B1(n_667), .B2(n_668), .C(n_670), .Y(n_664) );
INVx2_ASAP7_75t_L g603 ( .A(n_542), .Y(n_603) );
AND2x2_ASAP7_75t_L g576 ( .A(n_543), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g666 ( .A(n_543), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_543), .B(n_658), .Y(n_679) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVxp67_ASAP7_75t_L g621 ( .A(n_544), .Y(n_621) );
AND2x2_ASAP7_75t_L g657 ( .A(n_544), .B(n_658), .Y(n_657) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B(n_552), .Y(n_544) );
AND2x2_ASAP7_75t_L g659 ( .A(n_553), .B(n_598), .Y(n_659) );
AND2x2_ASAP7_75t_L g569 ( .A(n_554), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_554), .B(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_SL g640 ( .A(n_556), .B(n_603), .Y(n_640) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g646 ( .A(n_559), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
OR2x2_ASAP7_75t_L g632 ( .A(n_560), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g697 ( .A(n_560), .B(n_642), .Y(n_697) );
INVx2_ASAP7_75t_L g630 ( .A(n_561), .Y(n_630) );
NAND4xp25_ASAP7_75t_SL g693 ( .A(n_562), .B(n_694), .C(n_695), .D(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_563), .B(n_627), .Y(n_662) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_SL g699 ( .A(n_566), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_SL g661 ( .A1(n_567), .A2(n_630), .B(n_634), .C(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g656 ( .A(n_569), .B(n_648), .Y(n_656) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_570), .Y(n_582) );
INVx1_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_571), .Y(n_614) );
AOI211xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B(n_576), .C(n_578), .Y(n_572) );
AND2x2_ASAP7_75t_L g593 ( .A(n_573), .B(n_577), .Y(n_593) );
OAI322xp33_ASAP7_75t_SL g631 ( .A1(n_573), .A2(n_632), .A3(n_634), .B1(n_635), .B2(n_639), .C1(n_640), .C2(n_641), .Y(n_631) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g653 ( .A(n_575), .B(n_579), .Y(n_653) );
INVx1_ASAP7_75t_L g634 ( .A(n_577), .Y(n_634) );
INVx1_ASAP7_75t_SL g652 ( .A(n_579), .Y(n_652) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_591), .B1(n_593), .B2(n_594), .C1(n_595), .C2(n_727), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_586), .B(n_588), .Y(n_585) );
OAI322xp33_ASAP7_75t_L g674 ( .A1(n_586), .A2(n_648), .A3(n_653), .B1(n_675), .B2(n_676), .C1(n_678), .C2(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_587), .A2(n_601), .B1(n_625), .B2(n_629), .C(n_631), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
OAI222xp33_ASAP7_75t_L g604 ( .A1(n_592), .A2(n_605), .B1(n_607), .B2(n_608), .C1(n_609), .C2(n_612), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_594), .A2(n_601), .B1(n_671), .B2(n_672), .Y(n_670) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AOI211xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_604), .C(n_615), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_601), .A2(n_638), .B(n_681), .C(n_684), .Y(n_680) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g610 ( .A(n_602), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g673 ( .A(n_606), .Y(n_673) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_613), .B(n_638), .Y(n_667) );
BUFx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_618), .B(n_622), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g684 ( .A1(n_616), .A2(n_685), .B1(n_686), .B2(n_687), .C(n_688), .Y(n_684) );
INVxp33_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_620), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_627), .B(n_638), .Y(n_678) );
INVx2_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AND2x2_ASAP7_75t_L g689 ( .A(n_642), .B(n_648), .Y(n_689) );
AND4x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_663), .C(n_680), .D(n_692), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI221xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_651), .B1(n_653), .B2(n_654), .C(n_655), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_655) );
INVx1_ASAP7_75t_L g685 ( .A(n_656), .Y(n_685) );
INVx1_ASAP7_75t_SL g675 ( .A(n_660), .Y(n_675) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_674), .Y(n_663) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_676), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_683), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g709 ( .A(n_702), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx3_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
XNOR2xp5_ASAP7_75t_SL g716 ( .A(n_717), .B(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
endmodule