module fake_netlist_6_3122_n_1801 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1801);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1801;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_16),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_29),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_32),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_10),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_30),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_17),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_15),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_7),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_100),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_34),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_80),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_123),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_118),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_46),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_72),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_43),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_32),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_8),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_68),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_66),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_58),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_10),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_76),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

BUFx8_ASAP7_75t_SL g204 ( 
.A(n_143),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_55),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_83),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_46),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_22),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_33),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_115),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_152),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_36),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_149),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_78),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_151),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_131),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_104),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_119),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_94),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_125),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_20),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_65),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_12),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_81),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_79),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_7),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_30),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_33),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_145),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_24),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_18),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_89),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_97),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_63),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_52),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_31),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_19),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_116),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_117),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_28),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_40),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_11),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_128),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_45),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_110),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_37),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_18),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_154),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_67),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_127),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_157),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_12),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_25),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_41),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_108),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_20),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_122),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_38),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_29),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_156),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_35),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_84),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_126),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_48),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_9),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_95),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_134),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_4),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_139),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_59),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_93),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_136),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_25),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_41),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_133),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_158),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_70),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_51),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_45),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_27),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_69),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_13),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_35),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_31),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_82),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_147),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_64),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_56),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_90),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_2),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_51),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_38),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_144),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_96),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_148),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_146),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_43),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_135),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_57),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_120),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_153),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_140),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_28),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_141),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_193),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_167),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_193),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_193),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_193),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_204),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_187),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_193),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_231),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_185),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_246),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_246),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_298),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_191),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_246),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_194),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_246),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_288),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_246),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_163),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_163),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_200),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_179),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_202),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_165),
.Y(n_340)
);

INVxp33_ASAP7_75t_SL g341 ( 
.A(n_189),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_249),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_160),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_203),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_190),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_160),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_227),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_207),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_227),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_211),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_212),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_214),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_215),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_168),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_217),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_161),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_227),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_168),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_219),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_162),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_170),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_229),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_177),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_221),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_171),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_222),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_208),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_171),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_228),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_302),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_229),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_233),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_237),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_238),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_209),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_225),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_230),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_235),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_240),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_248),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_243),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_256),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_241),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_257),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_165),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_169),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_169),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_318),
.B(n_305),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_386),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_341),
.A2(n_265),
.B1(n_314),
.B2(n_259),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_333),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_386),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_325),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_319),
.B(n_175),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_319),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_322),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_351),
.B(n_175),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_374),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_376),
.B(n_362),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_323),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_328),
.A2(n_282),
.B1(n_181),
.B2(n_174),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_180),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_326),
.B(n_180),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_367),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_337),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_334),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_340),
.B(n_344),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_321),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_362),
.B(n_182),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_340),
.B(n_266),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_335),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_361),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_335),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_331),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_336),
.A2(n_263),
.B(n_255),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_345),
.A2(n_284),
.B1(n_174),
.B2(n_173),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_366),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_368),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_342),
.B(n_248),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_373),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_343),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_344),
.B(n_348),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_348),
.B(n_182),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_343),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_339),
.B(n_297),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_305),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_428),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_352),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_159),
.Y(n_469)
);

INVx6_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_412),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_353),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_394),
.B(n_355),
.Y(n_473)
);

NOR2x1p5_ASAP7_75t_L g474 ( 
.A(n_403),
.B(n_324),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_394),
.B(n_356),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

NOR2x1p5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_338),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_412),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_423),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_426),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_407),
.A2(n_347),
.B1(n_350),
.B2(n_346),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_397),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_423),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_439),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_434),
.B(n_359),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_423),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_407),
.B(n_360),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_439),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_408),
.Y(n_493)
);

BUFx6f_ASAP7_75t_SL g494 ( 
.A(n_433),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_458),
.B(n_317),
.C(n_369),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_435),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_425),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_461),
.B(n_372),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_425),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_445),
.A2(n_266),
.B1(n_358),
.B2(n_303),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_413),
.B(n_375),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_379),
.Y(n_504)
);

AO21x2_ASAP7_75t_L g505 ( 
.A1(n_395),
.A2(n_166),
.B(n_164),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_395),
.B(n_380),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_458),
.B(n_390),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_427),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

AND3x2_ASAP7_75t_L g511 ( 
.A(n_414),
.B(n_195),
.C(n_159),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_415),
.B(n_357),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_SL g513 ( 
.A1(n_417),
.A2(n_302),
.B1(n_181),
.B2(n_284),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_405),
.B(n_261),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_438),
.B(n_364),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_435),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_405),
.B(n_378),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_418),
.B(n_387),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_396),
.B(n_382),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_392),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_422),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_399),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_397),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_436),
.B(n_352),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_418),
.B(n_264),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_397),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_399),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_406),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_427),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_397),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_410),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_442),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_445),
.A2(n_268),
.B1(n_283),
.B2(n_293),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_422),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_401),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_411),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_419),
.B(n_388),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_442),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_411),
.Y(n_543)
);

NOR2x1p5_ASAP7_75t_L g544 ( 
.A(n_456),
.B(n_173),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_420),
.B(n_354),
.Y(n_545)
);

AOI21x1_ASAP7_75t_L g546 ( 
.A1(n_424),
.A2(n_205),
.B(n_195),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_424),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_442),
.Y(n_548)
);

AND3x2_ASAP7_75t_L g549 ( 
.A(n_420),
.B(n_205),
.C(n_196),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_393),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_401),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_435),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_442),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_431),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_419),
.B(n_183),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_442),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_393),
.B(n_183),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_431),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_397),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_398),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_417),
.A2(n_287),
.B1(n_236),
.B2(n_307),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_446),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_444),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_444),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_445),
.A2(n_308),
.B1(n_365),
.B2(n_248),
.Y(n_566)
);

NAND3xp33_ASAP7_75t_L g567 ( 
.A(n_400),
.B(n_354),
.C(n_186),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_436),
.B(n_383),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_400),
.A2(n_281),
.B1(n_282),
.B2(n_289),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_445),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_446),
.A2(n_242),
.B1(n_239),
.B2(n_251),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_445),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_456),
.B(n_184),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_433),
.B(n_184),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_433),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_433),
.B(n_236),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_435),
.B(n_267),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_441),
.B(n_389),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_396),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_441),
.B(n_285),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_448),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_435),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_448),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_435),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_437),
.B(n_273),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_437),
.B(n_274),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_449),
.B(n_285),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_437),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_444),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_437),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_437),
.B(n_248),
.Y(n_591)
);

AND2x2_ASAP7_75t_SL g592 ( 
.A(n_437),
.B(n_248),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_402),
.B(n_404),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_444),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_460),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_449),
.Y(n_597)
);

OAI21xp33_ASAP7_75t_SL g598 ( 
.A1(n_450),
.A2(n_389),
.B(n_385),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_398),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_450),
.B(n_286),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_452),
.B(n_383),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_444),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_459),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_452),
.B(n_286),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_402),
.B(n_404),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_402),
.B(n_277),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_459),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_460),
.A2(n_295),
.B1(n_385),
.B2(n_384),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_453),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_459),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_460),
.A2(n_295),
.B1(n_384),
.B2(n_199),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_453),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_459),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_507),
.B(n_447),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_570),
.A2(n_201),
.B1(n_295),
.B2(n_229),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_570),
.A2(n_572),
.B1(n_501),
.B2(n_537),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_447),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_473),
.B(n_287),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_504),
.B(n_457),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_581),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_475),
.B(n_296),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_562),
.A2(n_281),
.B1(n_289),
.B2(n_290),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_447),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_SL g625 ( 
.A(n_572),
.B(n_295),
.Y(n_625)
);

OAI22xp33_ASAP7_75t_L g626 ( 
.A1(n_561),
.A2(n_290),
.B1(n_301),
.B2(n_294),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_469),
.B(n_229),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_613),
.B(n_447),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_550),
.B(n_457),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_459),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_550),
.B(n_462),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_568),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_476),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_519),
.B(n_296),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_568),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_476),
.B(n_416),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_592),
.B(n_295),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_545),
.A2(n_292),
.B1(n_301),
.B2(n_294),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_583),
.B(n_304),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_583),
.B(n_462),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_601),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_578),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_480),
.B(n_416),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_583),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_578),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_506),
.B(n_304),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_472),
.B(n_307),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_592),
.B(n_229),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_502),
.A2(n_279),
.B1(n_315),
.B2(n_280),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_573),
.B(n_192),
.C(n_210),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_468),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_592),
.B(n_229),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_597),
.B(n_463),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_469),
.B(n_229),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_524),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_525),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_471),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_525),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_480),
.B(n_416),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_481),
.B(n_416),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_524),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_481),
.B(n_579),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_471),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_478),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_597),
.B(n_311),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_L g669 ( 
.A(n_515),
.B(n_541),
.C(n_518),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_488),
.B(n_311),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_579),
.B(n_416),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_467),
.B(n_463),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_495),
.B(n_213),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_517),
.B(n_292),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_555),
.A2(n_526),
.B(n_514),
.C(n_521),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_467),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_520),
.B(n_172),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_503),
.B(n_416),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_486),
.B(n_216),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_503),
.B(n_521),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_478),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_523),
.B(n_421),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_523),
.B(n_421),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_465),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_469),
.A2(n_178),
.B1(n_313),
.B2(n_312),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_566),
.B(n_229),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_601),
.B(n_463),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_528),
.B(n_421),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_528),
.B(n_421),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_575),
.B(n_232),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_482),
.B(n_176),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_529),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_529),
.B(n_421),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_497),
.B(n_234),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_474),
.B(n_188),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_601),
.Y(n_696)
);

AND2x6_ASAP7_75t_SL g697 ( 
.A(n_513),
.B(n_197),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_520),
.B(n_250),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_577),
.A2(n_398),
.B(n_404),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_479),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_490),
.B(n_245),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_465),
.B(n_440),
.Y(n_702)
);

OAI221xp5_ASAP7_75t_L g703 ( 
.A1(n_598),
.A2(n_198),
.B1(n_206),
.B2(n_220),
.C(n_223),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_499),
.B(n_247),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_469),
.B(n_250),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_567),
.B(n_252),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_600),
.B(n_258),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_530),
.B(n_421),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_520),
.B(n_224),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_580),
.B(n_226),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_604),
.B(n_260),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_469),
.B(n_250),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_532),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_587),
.A2(n_291),
.B(n_253),
.C(n_254),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_535),
.B(n_250),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_535),
.B(n_429),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_505),
.A2(n_250),
.B1(n_270),
.B2(n_244),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_540),
.B(n_429),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_479),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_543),
.B(n_250),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_543),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_485),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_SL g723 ( 
.A(n_494),
.B(n_276),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_547),
.B(n_429),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_470),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_574),
.B(n_576),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_465),
.B(n_306),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_547),
.B(n_429),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_554),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_554),
.B(n_262),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_549),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_558),
.B(n_271),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_558),
.B(n_275),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_470),
.B(n_429),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_469),
.B(n_250),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_469),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_470),
.B(n_429),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_596),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_534),
.B(n_250),
.Y(n_739)
);

AND2x6_ASAP7_75t_SL g740 ( 
.A(n_522),
.B(n_310),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_470),
.B(n_430),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_SL g742 ( 
.A(n_494),
.B(n_269),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_596),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_569),
.B(n_571),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_512),
.A2(n_309),
.B1(n_299),
.B2(n_278),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_485),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_505),
.B(n_430),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_505),
.B(n_496),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_582),
.B(n_430),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_606),
.B(n_455),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_582),
.B(n_430),
.Y(n_751)
);

BUFx6f_ASAP7_75t_SL g752 ( 
.A(n_494),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_544),
.A2(n_270),
.B1(n_451),
.B2(n_440),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_584),
.B(n_430),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_584),
.B(n_588),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_493),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_585),
.B(n_455),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_588),
.B(n_430),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_590),
.B(n_409),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_522),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_538),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_590),
.B(n_409),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_474),
.B(n_455),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_586),
.B(n_270),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_516),
.B(n_552),
.Y(n_765)
);

INVx8_ASAP7_75t_L g766 ( 
.A(n_538),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_487),
.A2(n_440),
.B(n_409),
.C(n_451),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_608),
.B(n_270),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_516),
.B(n_398),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_593),
.Y(n_770)
);

NOR2x1p5_ASAP7_75t_L g771 ( 
.A(n_551),
.B(n_0),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_516),
.B(n_398),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_489),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_544),
.B(n_150),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_552),
.B(n_451),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_605),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_552),
.B(n_451),
.Y(n_777)
);

INVx8_ASAP7_75t_L g778 ( 
.A(n_551),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_483),
.B(n_451),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_539),
.B(n_270),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_477),
.B(n_270),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_483),
.B(n_451),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_620),
.B(n_477),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_702),
.Y(n_784)
);

NOR2x1p5_ASAP7_75t_L g785 ( 
.A(n_645),
.B(n_466),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_629),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_725),
.B(n_614),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_687),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_687),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_641),
.B(n_524),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_648),
.B(n_487),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_692),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_725),
.B(n_534),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_648),
.B(n_491),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_642),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_713),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_655),
.B(n_492),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_657),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_639),
.Y(n_799)
);

BUFx8_ASAP7_75t_SL g800 ( 
.A(n_761),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_615),
.B(n_536),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_756),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_619),
.A2(n_614),
.B(n_536),
.C(n_611),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_721),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_729),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_631),
.B(n_511),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_672),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_654),
.B(n_492),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_657),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_647),
.B(n_483),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_621),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_756),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_760),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_738),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_743),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_632),
.B(n_542),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_642),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_726),
.A2(n_553),
.B1(n_611),
.B2(n_610),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_696),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_766),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_616),
.A2(n_270),
.B1(n_489),
.B2(n_498),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_619),
.B(n_484),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_622),
.B(n_484),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_616),
.B(n_270),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_622),
.B(n_484),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_696),
.B(n_542),
.Y(n_826)
);

CKINVDCx11_ASAP7_75t_R g827 ( 
.A(n_740),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_635),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_645),
.B(n_524),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_647),
.B(n_527),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_657),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_662),
.B(n_524),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_652),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_633),
.B(n_527),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_717),
.A2(n_500),
.B1(n_510),
.B2(n_509),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_736),
.B(n_548),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_665),
.B(n_527),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_662),
.B(n_533),
.Y(n_838)
);

AND2x6_ASAP7_75t_SL g839 ( 
.A(n_744),
.B(n_0),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_770),
.B(n_776),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_643),
.B(n_548),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_646),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_680),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_617),
.B(n_591),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_659),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_617),
.B(n_658),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_657),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_684),
.B(n_553),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_674),
.B(n_556),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_676),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_760),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_660),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_763),
.B(n_556),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_666),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_667),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_744),
.A2(n_531),
.B1(n_510),
.B2(n_509),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_681),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_766),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_726),
.A2(n_564),
.B1(n_610),
.B2(n_607),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_675),
.B(n_564),
.Y(n_860)
);

NOR2xp67_ASAP7_75t_L g861 ( 
.A(n_651),
.B(n_589),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_763),
.B(n_595),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_731),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_634),
.B(n_565),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_669),
.B(n_594),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_781),
.B(n_565),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_700),
.Y(n_867)
);

BUFx12f_ASAP7_75t_SL g868 ( 
.A(n_695),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_730),
.B(n_565),
.Y(n_869)
);

AO21x2_ASAP7_75t_L g870 ( 
.A1(n_748),
.A2(n_546),
.B(n_607),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_679),
.B(n_612),
.C(n_603),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_719),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_730),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_742),
.A2(n_498),
.B1(n_500),
.B2(n_508),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_732),
.B(n_560),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_766),
.B(n_546),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_722),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_746),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_717),
.A2(n_508),
.B1(n_531),
.B2(n_591),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_773),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_778),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_752),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_763),
.B(n_695),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_664),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_732),
.B(n_560),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_618),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_706),
.A2(n_603),
.B1(n_602),
.B2(n_563),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_664),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_679),
.B(n_602),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_755),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_R g891 ( 
.A(n_778),
.B(n_101),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_706),
.A2(n_563),
.B1(n_595),
.B2(n_594),
.Y(n_892)
);

CKINVDCx6p67_ASAP7_75t_R g893 ( 
.A(n_752),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_664),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_664),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_626),
.B(n_694),
.Y(n_896)
);

AND2x6_ASAP7_75t_L g897 ( 
.A(n_736),
.B(n_589),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_624),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_628),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_677),
.A2(n_560),
.B1(n_599),
.B2(n_591),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_759),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_626),
.B(n_599),
.Y(n_902)
);

NOR2x1_ASAP7_75t_L g903 ( 
.A(n_695),
.B(n_599),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_733),
.B(n_559),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_677),
.A2(n_591),
.B1(n_559),
.B2(n_533),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_774),
.B(n_559),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_750),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_734),
.A2(n_559),
.B(n_533),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_677),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_678),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_682),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_694),
.B(n_1),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_762),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_774),
.B(n_559),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_636),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_778),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_650),
.B(n_130),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_709),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_677),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_690),
.B(n_533),
.Y(n_920)
);

NOR2x2_ASAP7_75t_L g921 ( 
.A(n_697),
.B(n_1),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_644),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_750),
.B(n_533),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_670),
.B(n_3),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_637),
.A2(n_591),
.B1(n_124),
.B2(n_112),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_SL g926 ( 
.A(n_623),
.B(n_3),
.C(n_4),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_661),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_677),
.Y(n_928)
);

BUFx4f_ASAP7_75t_L g929 ( 
.A(n_771),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_757),
.B(n_591),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_683),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_698),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_701),
.B(n_704),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_704),
.B(n_5),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_SL g935 ( 
.A1(n_701),
.A2(n_591),
.B1(n_6),
.B2(n_8),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_688),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_SL g937 ( 
.A1(n_673),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_689),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_693),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_673),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_757),
.B(n_451),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_707),
.B(n_451),
.Y(n_942)
);

BUFx10_ASAP7_75t_L g943 ( 
.A(n_707),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_708),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_671),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_640),
.B(n_13),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_711),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_649),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_723),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_780),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_SL g951 ( 
.A1(n_711),
.A2(n_14),
.B1(n_19),
.B2(n_21),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_668),
.B(n_21),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_691),
.B(n_23),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_698),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_745),
.B(n_105),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_710),
.B(n_23),
.Y(n_956)
);

CKINVDCx11_ASAP7_75t_R g957 ( 
.A(n_623),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_630),
.B(n_24),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_716),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_718),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_779),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_637),
.B(n_27),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_782),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_625),
.B(n_36),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_745),
.B(n_103),
.Y(n_965)
);

OAI21xp33_ASAP7_75t_L g966 ( 
.A1(n_638),
.A2(n_37),
.B(n_39),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_727),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_663),
.B(n_39),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_765),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_753),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_798),
.Y(n_971)
);

AOI33xp33_ASAP7_75t_L g972 ( 
.A1(n_948),
.A2(n_638),
.A3(n_685),
.B1(n_767),
.B2(n_703),
.B3(n_714),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_786),
.B(n_747),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_907),
.A2(n_686),
.B1(n_649),
.B2(n_653),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_843),
.B(n_728),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_933),
.B(n_724),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_896),
.A2(n_686),
.B1(n_653),
.B2(n_720),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_SL g978 ( 
.A(n_947),
.B(n_715),
.C(n_720),
.Y(n_978)
);

OAI22x1_ASAP7_75t_L g979 ( 
.A1(n_896),
.A2(n_715),
.B1(n_739),
.B2(n_768),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_934),
.A2(n_627),
.B(n_705),
.C(n_712),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_802),
.B(n_739),
.Y(n_981)
);

BUFx12f_ASAP7_75t_L g982 ( 
.A(n_882),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_784),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_816),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_792),
.Y(n_985)
);

BUFx12f_ASAP7_75t_L g986 ( 
.A(n_785),
.Y(n_986)
);

CKINVDCx11_ASAP7_75t_R g987 ( 
.A(n_827),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_934),
.A2(n_656),
.B(n_735),
.C(n_764),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_812),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_841),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_844),
.A2(n_737),
.B(n_741),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_873),
.B(n_758),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_873),
.B(n_775),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_786),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_860),
.A2(n_754),
.B(n_751),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_799),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_SL g997 ( 
.A(n_949),
.B(n_777),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_783),
.A2(n_749),
.B(n_769),
.C(n_772),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_940),
.B(n_699),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_800),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_943),
.B(n_102),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_863),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_849),
.B(n_42),
.Y(n_1003)
);

INVx8_ASAP7_75t_L g1004 ( 
.A(n_897),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_813),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_840),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_884),
.A2(n_62),
.B(n_91),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_SL g1008 ( 
.A1(n_949),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_796),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_L g1010 ( 
.A(n_946),
.B(n_49),
.C(n_50),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_943),
.B(n_73),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_879),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_863),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_R g1014 ( 
.A(n_970),
.B(n_71),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_883),
.B(n_75),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_SL g1016 ( 
.A(n_884),
.B(n_53),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_833),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_890),
.B(n_85),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_845),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_804),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_946),
.A2(n_952),
.B(n_966),
.C(n_912),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_851),
.B(n_807),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_952),
.A2(n_902),
.B(n_846),
.C(n_918),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_953),
.A2(n_92),
.B1(n_932),
.B2(n_789),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_897),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_798),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_811),
.B(n_850),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_806),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_908),
.A2(n_860),
.B(n_961),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_884),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_805),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_956),
.A2(n_902),
.B(n_924),
.C(n_955),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_SL g1033 ( 
.A(n_951),
.B(n_917),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_798),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_850),
.B(n_819),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_884),
.A2(n_894),
.B(n_923),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_965),
.A2(n_811),
.B(n_962),
.C(n_865),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_808),
.B(n_886),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_798),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_808),
.B(n_898),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_820),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_803),
.A2(n_824),
.B(n_871),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_858),
.B(n_881),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_899),
.B(n_915),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_809),
.Y(n_1045)
);

CKINVDCx6p67_ASAP7_75t_R g1046 ( 
.A(n_893),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_814),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_819),
.B(n_903),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_879),
.A2(n_948),
.B1(n_821),
.B2(n_935),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_922),
.B(n_927),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_815),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_865),
.A2(n_914),
.B(n_906),
.C(n_918),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_828),
.Y(n_1053)
);

BUFx10_ASAP7_75t_L g1054 ( 
.A(n_853),
.Y(n_1054)
);

OA22x2_ASAP7_75t_L g1055 ( 
.A1(n_937),
.A2(n_852),
.B1(n_842),
.B2(n_967),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_821),
.A2(n_935),
.B1(n_954),
.B2(n_932),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_950),
.B(n_788),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_901),
.B(n_913),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_855),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_957),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_SL g1061 ( 
.A(n_891),
.B(n_926),
.C(n_876),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_797),
.B(n_910),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_911),
.B(n_931),
.Y(n_1063)
);

AO21x2_ASAP7_75t_L g1064 ( 
.A1(n_856),
.A2(n_904),
.B(n_801),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_967),
.B(n_954),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_889),
.B(n_791),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_894),
.A2(n_866),
.B(n_822),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_958),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_894),
.A2(n_823),
.B(n_825),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_894),
.B(n_809),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_795),
.B(n_969),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_809),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_929),
.B(n_916),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_810),
.A2(n_830),
.B(n_864),
.C(n_794),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_854),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_906),
.A2(n_914),
.B1(n_835),
.B2(n_926),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_809),
.Y(n_1077)
);

BUFx8_ASAP7_75t_L g1078 ( 
.A(n_853),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_936),
.B(n_938),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_826),
.A2(n_817),
.B1(n_862),
.B2(n_848),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_857),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_969),
.B(n_929),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_969),
.B(n_862),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_867),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_891),
.B(n_944),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_848),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_868),
.B(n_810),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_847),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_969),
.B(n_826),
.Y(n_1089)
);

AOI22x1_ASAP7_75t_L g1090 ( 
.A1(n_939),
.A2(n_960),
.B1(n_959),
.B2(n_945),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_968),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_830),
.B(n_945),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_864),
.A2(n_875),
.B(n_869),
.C(n_885),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_847),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_835),
.A2(n_836),
.B1(n_930),
.B2(n_928),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_921),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_861),
.A2(n_942),
.B(n_909),
.C(n_963),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_847),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_909),
.A2(n_963),
.B(n_961),
.C(n_818),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_872),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_847),
.B(n_888),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_834),
.A2(n_837),
.B(n_793),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_856),
.B(n_880),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_919),
.B(n_928),
.Y(n_1104)
);

NOR2xp67_ASAP7_75t_L g1105 ( 
.A(n_920),
.B(n_877),
.Y(n_1105)
);

INVxp67_ASAP7_75t_L g1106 ( 
.A(n_878),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_964),
.A2(n_790),
.B(n_874),
.C(n_838),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_888),
.Y(n_1108)
);

O2A1O1Ixp5_ASAP7_75t_L g1109 ( 
.A1(n_801),
.A2(n_941),
.B(n_832),
.C(n_829),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_859),
.A2(n_892),
.B(n_887),
.C(n_900),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_839),
.B(n_831),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_876),
.B(n_870),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_831),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_895),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_919),
.B(n_928),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_874),
.A2(n_787),
.B(n_793),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_888),
.B(n_928),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_787),
.A2(n_888),
.B(n_836),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_897),
.B(n_895),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_919),
.B(n_905),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_919),
.B(n_897),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_925),
.A2(n_870),
.B(n_897),
.Y(n_1122)
);

AO22x1_ASAP7_75t_L g1123 ( 
.A1(n_947),
.A2(n_896),
.B1(n_934),
.B2(n_946),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_980),
.A2(n_988),
.B(n_1093),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1074),
.A2(n_1042),
.B(n_1110),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1073),
.B(n_1048),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1042),
.A2(n_977),
.B(n_974),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_987),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1102),
.A2(n_1069),
.B(n_1092),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1085),
.B(n_1033),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1029),
.A2(n_995),
.B(n_991),
.Y(n_1131)
);

AO21x1_ASAP7_75t_L g1132 ( 
.A1(n_1049),
.A2(n_1021),
.B(n_1032),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1028),
.Y(n_1133)
);

OAI22x1_ASAP7_75t_L g1134 ( 
.A1(n_1111),
.A2(n_1065),
.B1(n_1087),
.B2(n_1123),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_985),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1040),
.B(n_1062),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1049),
.A2(n_1012),
.B1(n_1056),
.B2(n_1023),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_1025),
.B(n_1030),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_SL g1140 ( 
.A1(n_1006),
.A2(n_976),
.B(n_1012),
.C(n_1001),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1118),
.A2(n_1122),
.B(n_1067),
.Y(n_1141)
);

CKINVDCx11_ASAP7_75t_R g1142 ( 
.A(n_982),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_1097),
.A2(n_1099),
.A3(n_1095),
.B(n_979),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1063),
.B(n_1079),
.Y(n_1144)
);

OA22x2_ASAP7_75t_L g1145 ( 
.A1(n_1096),
.A2(n_1006),
.B1(n_1013),
.B2(n_1002),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_974),
.A2(n_1095),
.B(n_977),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1036),
.A2(n_1116),
.B(n_1090),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1048),
.B(n_1082),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1116),
.A2(n_1109),
.B(n_998),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1026),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_989),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1058),
.B(n_984),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1056),
.A2(n_1076),
.B(n_1037),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1078),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1046),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1027),
.B(n_1033),
.Y(n_1156)
);

NAND2x1_ASAP7_75t_L g1157 ( 
.A(n_1030),
.B(n_1104),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1004),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1061),
.A2(n_1055),
.B1(n_1015),
.B2(n_1091),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1103),
.A2(n_993),
.B(n_1105),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1004),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_990),
.B(n_1068),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1103),
.A2(n_1071),
.B(n_1120),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_975),
.A2(n_1025),
.B(n_999),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1055),
.A2(n_1010),
.B1(n_1024),
.B2(n_983),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1025),
.A2(n_1064),
.B(n_997),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_1005),
.Y(n_1167)
);

NOR4xp25_ASAP7_75t_L g1168 ( 
.A(n_1076),
.B(n_1091),
.C(n_1068),
.D(n_1052),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_SL g1169 ( 
.A(n_1025),
.B(n_1016),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1121),
.A2(n_1107),
.B(n_1119),
.Y(n_1170)
);

AO22x2_ASAP7_75t_L g1171 ( 
.A1(n_1112),
.A2(n_1003),
.B1(n_1035),
.B2(n_973),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1009),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1008),
.B(n_978),
.C(n_992),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1080),
.B(n_972),
.C(n_1011),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1044),
.B(n_1050),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1050),
.B(n_1020),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1018),
.A2(n_1059),
.B(n_1084),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1106),
.B(n_1022),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1064),
.A2(n_997),
.B(n_1089),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1026),
.Y(n_1180)
);

NOR4xp25_ASAP7_75t_L g1181 ( 
.A(n_1053),
.B(n_1083),
.C(n_1051),
.D(n_1031),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1004),
.A2(n_1121),
.B(n_1101),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_1007),
.A2(n_1117),
.B(n_1113),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1047),
.B(n_1017),
.Y(n_1184)
);

AOI21xp33_ASAP7_75t_L g1185 ( 
.A1(n_1014),
.A2(n_1100),
.B(n_981),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_996),
.A2(n_1019),
.B(n_1075),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1086),
.B(n_1081),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1114),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1057),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1104),
.A2(n_1115),
.B(n_971),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1104),
.A2(n_1115),
.B(n_1070),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_SL g1192 ( 
.A1(n_1115),
.A2(n_1117),
.B(n_1015),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_981),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1043),
.B(n_981),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1034),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1060),
.A2(n_1043),
.B(n_1034),
.C(n_1088),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1039),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1077),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1077),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1060),
.B(n_1054),
.Y(n_1200)
);

OAI21xp33_ASAP7_75t_L g1201 ( 
.A1(n_1094),
.A2(n_1108),
.B(n_1088),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1070),
.A2(n_1039),
.B(n_1045),
.Y(n_1202)
);

CKINVDCx14_ASAP7_75t_R g1203 ( 
.A(n_986),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1039),
.A2(n_1045),
.B(n_1072),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1072),
.A2(n_725),
.B(n_980),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1098),
.A2(n_1029),
.B(n_995),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1098),
.B(n_1066),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1073),
.B(n_1048),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_985),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_1025),
.B(n_1030),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1028),
.B(n_786),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_SL g1218 ( 
.A1(n_1052),
.A2(n_1037),
.B(n_1021),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1028),
.B(n_786),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1029),
.A2(n_995),
.B(n_991),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1021),
.A2(n_896),
.B1(n_1123),
.B2(n_947),
.C(n_934),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_987),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_994),
.B(n_493),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1074),
.A2(n_1093),
.B(n_896),
.Y(n_1226)
);

BUFx8_ASAP7_75t_SL g1227 ( 
.A(n_1000),
.Y(n_1227)
);

O2A1O1Ixp5_ASAP7_75t_L g1228 ( 
.A1(n_1123),
.A2(n_934),
.B(n_907),
.C(n_896),
.Y(n_1228)
);

BUFx4f_ASAP7_75t_SL g1229 ( 
.A(n_982),
.Y(n_1229)
);

OAI31xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1049),
.A2(n_934),
.A3(n_896),
.B(n_912),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1029),
.A2(n_995),
.B(n_991),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_994),
.Y(n_1232)
);

OAI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1111),
.A2(n_896),
.B1(n_947),
.B2(n_934),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1042),
.A2(n_1093),
.B(n_1029),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1093),
.A2(n_1074),
.A3(n_1110),
.B(n_1097),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1123),
.B(n_934),
.C(n_896),
.Y(n_1236)
);

AOI21xp33_ASAP7_75t_L g1237 ( 
.A1(n_1021),
.A2(n_907),
.B(n_934),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1026),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_L g1239 ( 
.A1(n_1033),
.A2(n_896),
.B(n_934),
.Y(n_1239)
);

AO21x1_ASAP7_75t_L g1240 ( 
.A1(n_1049),
.A2(n_934),
.B(n_907),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1029),
.A2(n_995),
.B(n_991),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1073),
.B(n_1048),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_983),
.B(n_949),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1041),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1248)
);

AOI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1021),
.A2(n_896),
.B1(n_1123),
.B2(n_947),
.C(n_934),
.Y(n_1249)
);

AOI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1069),
.A2(n_860),
.B(n_995),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1029),
.A2(n_995),
.B(n_991),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1074),
.A2(n_1093),
.B(n_896),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_983),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1123),
.B(n_947),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_982),
.Y(n_1255)
);

OAI21xp33_ASAP7_75t_L g1256 ( 
.A1(n_1033),
.A2(n_896),
.B(n_934),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1066),
.B(n_907),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1026),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1028),
.B(n_786),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1066),
.B(n_907),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_985),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1029),
.A2(n_995),
.B(n_991),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1123),
.B(n_947),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1066),
.B(n_1038),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_980),
.A2(n_725),
.B(n_988),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_983),
.B(n_949),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1021),
.A2(n_896),
.B(n_934),
.C(n_933),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1028),
.B(n_786),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1042),
.A2(n_1093),
.B(n_1029),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1004),
.B(n_858),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1066),
.B(n_907),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_983),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1172),
.Y(n_1275)
);

NAND2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1157),
.B(n_1158),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1236),
.A2(n_1256),
.B1(n_1239),
.B2(n_1156),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1158),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1153),
.A2(n_1149),
.B(n_1129),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1241),
.A2(n_1262),
.B(n_1251),
.Y(n_1280)
);

AOI21xp33_ASAP7_75t_L g1281 ( 
.A1(n_1236),
.A2(n_1249),
.B(n_1223),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1136),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1130),
.B(n_1135),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1141),
.A2(n_1250),
.B(n_1206),
.Y(n_1284)
);

AOI31xp67_ASAP7_75t_L g1285 ( 
.A1(n_1145),
.A2(n_1159),
.A3(n_1260),
.B(n_1273),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1186),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1209),
.A2(n_1215),
.B(n_1211),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1217),
.B(n_1219),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1259),
.B(n_1270),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1148),
.B(n_1161),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1218),
.A2(n_1127),
.B(n_1166),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1147),
.A2(n_1216),
.B(n_1222),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1127),
.A2(n_1237),
.B(n_1153),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1212),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1142),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1146),
.A2(n_1125),
.B(n_1252),
.Y(n_1296)
);

NOR2x1_ASAP7_75t_SL g1297 ( 
.A(n_1160),
.B(n_1272),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1155),
.B(n_1229),
.Y(n_1298)
);

OR3x4_ASAP7_75t_SL g1299 ( 
.A(n_1233),
.B(n_1254),
.C(n_1265),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1133),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1132),
.A2(n_1138),
.B1(n_1237),
.B2(n_1240),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1208),
.B(n_1214),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1221),
.B(n_1243),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1227),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1138),
.A2(n_1269),
.A3(n_1124),
.B(n_1179),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1263),
.A2(n_1264),
.B(n_1267),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1261),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1125),
.A2(n_1252),
.B(n_1226),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1184),
.Y(n_1309)
);

AO21x1_ASAP7_75t_L g1310 ( 
.A1(n_1226),
.A2(n_1164),
.B(n_1273),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1183),
.A2(n_1205),
.A3(n_1230),
.B(n_1134),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1163),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1181),
.A2(n_1168),
.B(n_1170),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1244),
.B(n_1246),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1248),
.B(n_1266),
.Y(n_1315)
);

BUFx5_ASAP7_75t_L g1316 ( 
.A(n_1198),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1230),
.A2(n_1260),
.A3(n_1257),
.B(n_1181),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1148),
.B(n_1161),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_SL g1319 ( 
.A1(n_1192),
.A2(n_1196),
.B(n_1191),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1257),
.A2(n_1182),
.A3(n_1168),
.B(n_1190),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1228),
.A2(n_1173),
.B(n_1144),
.C(n_1137),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1174),
.A2(n_1185),
.B(n_1173),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1126),
.B(n_1242),
.Y(n_1323)
);

CKINVDCx9p33_ASAP7_75t_R g1324 ( 
.A(n_1154),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1174),
.A2(n_1165),
.B(n_1137),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1144),
.B(n_1185),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1234),
.A2(n_1271),
.A3(n_1143),
.B(n_1207),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1271),
.A2(n_1140),
.B(n_1177),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1193),
.A2(n_1207),
.B(n_1167),
.C(n_1232),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1184),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1171),
.A2(n_1177),
.B(n_1145),
.Y(n_1331)
);

OAI221xp5_ASAP7_75t_L g1332 ( 
.A1(n_1225),
.A2(n_1162),
.B1(n_1178),
.B2(n_1193),
.C(n_1189),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1210),
.B(n_1242),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1169),
.A2(n_1171),
.B1(n_1194),
.B2(n_1175),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1169),
.A2(n_1176),
.B(n_1139),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1176),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1139),
.A2(n_1213),
.B(n_1202),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1152),
.B(n_1210),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_SL g1339 ( 
.A(n_1200),
.B(n_1201),
.C(n_1187),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1188),
.A2(n_1143),
.B(n_1235),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1204),
.A2(n_1199),
.B(n_1195),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1245),
.B(n_1268),
.C(n_1151),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1253),
.A2(n_1274),
.B(n_1143),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1235),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1203),
.A2(n_1255),
.B(n_1224),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1150),
.B(n_1180),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1150),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1258),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1197),
.A2(n_1238),
.B(n_1128),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1350)
);

NAND2x1p5_ASAP7_75t_L g1351 ( 
.A(n_1157),
.B(n_1025),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1162),
.B(n_1144),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1153),
.A2(n_1149),
.B(n_1129),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1172),
.Y(n_1354)
);

AO21x1_ASAP7_75t_L g1355 ( 
.A1(n_1237),
.A2(n_934),
.B(n_1138),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1247),
.Y(n_1356)
);

OAI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1239),
.A2(n_1256),
.B1(n_933),
.B2(n_896),
.C(n_947),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1228),
.A2(n_933),
.B(n_1269),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1172),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1150),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1135),
.B(n_1208),
.Y(n_1362)
);

AOI221x1_ASAP7_75t_L g1363 ( 
.A1(n_1239),
.A2(n_1256),
.B1(n_1236),
.B2(n_1237),
.C(n_1269),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1172),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1228),
.A2(n_933),
.B(n_1269),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1239),
.A2(n_947),
.B1(n_1256),
.B2(n_1033),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1247),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1148),
.B(n_1158),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1172),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1239),
.A2(n_1256),
.B1(n_896),
.B2(n_1249),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1172),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1236),
.A2(n_947),
.B1(n_1256),
.B2(n_1239),
.Y(n_1373)
);

AND2x6_ASAP7_75t_L g1374 ( 
.A(n_1158),
.B(n_1161),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1247),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1228),
.A2(n_933),
.B(n_1269),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1143),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1247),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1223),
.B(n_1249),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1247),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1157),
.B(n_1025),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1228),
.A2(n_933),
.B(n_1269),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1386)
);

BUFx10_ASAP7_75t_L g1387 ( 
.A(n_1155),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1218),
.A2(n_1127),
.B(n_1166),
.Y(n_1388)
);

INVx4_ASAP7_75t_SL g1389 ( 
.A(n_1272),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1236),
.A2(n_947),
.B1(n_1256),
.B2(n_1239),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1232),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1172),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1228),
.A2(n_933),
.B(n_1269),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1131),
.A2(n_1231),
.B(n_1220),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1239),
.A2(n_1256),
.B1(n_896),
.B2(n_1249),
.Y(n_1395)
);

INVx4_ASAP7_75t_SL g1396 ( 
.A(n_1272),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1172),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1239),
.A2(n_1256),
.B1(n_896),
.B2(n_1249),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1230),
.A2(n_1256),
.B(n_1239),
.C(n_1127),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1239),
.B(n_1256),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1162),
.B(n_1144),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1355),
.A2(n_1380),
.B(n_1281),
.C(n_1377),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1366),
.A2(n_1398),
.B1(n_1395),
.B2(n_1371),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1302),
.B(n_1303),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1371),
.A2(n_1398),
.B1(n_1395),
.B2(n_1315),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1302),
.B(n_1303),
.Y(n_1406)
);

O2A1O1Ixp5_ASAP7_75t_L g1407 ( 
.A1(n_1380),
.A2(n_1383),
.B(n_1365),
.C(n_1393),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1399),
.A2(n_1321),
.B(n_1357),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1315),
.A2(n_1283),
.B1(n_1314),
.B2(n_1362),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1328),
.A2(n_1306),
.B(n_1292),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1283),
.A2(n_1399),
.B1(n_1332),
.B2(n_1342),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1308),
.B(n_1317),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1317),
.B(n_1296),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1294),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1296),
.B(n_1291),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1300),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1296),
.B(n_1291),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1286),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1391),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1389),
.B(n_1396),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1373),
.A2(n_1390),
.B(n_1321),
.C(n_1277),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1388),
.B(n_1378),
.Y(n_1422)
);

O2A1O1Ixp5_ASAP7_75t_L g1423 ( 
.A1(n_1358),
.A2(n_1310),
.B(n_1400),
.C(n_1331),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1352),
.B(n_1401),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1326),
.B(n_1336),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1388),
.B(n_1293),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1293),
.B(n_1327),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1340),
.B(n_1326),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1400),
.A2(n_1301),
.B1(n_1334),
.B2(n_1338),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1391),
.Y(n_1430)
);

OA22x2_ASAP7_75t_L g1431 ( 
.A1(n_1319),
.A2(n_1363),
.B1(n_1309),
.B2(n_1330),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1301),
.A2(n_1334),
.B1(n_1329),
.B2(n_1325),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1292),
.A2(n_1287),
.B(n_1284),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1294),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1335),
.A2(n_1339),
.B(n_1344),
.C(n_1307),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1340),
.B(n_1344),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1307),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1279),
.A2(n_1353),
.B(n_1297),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1340),
.B(n_1320),
.Y(n_1439)
);

CKINVDCx16_ASAP7_75t_R g1440 ( 
.A(n_1304),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1389),
.B(n_1396),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1356),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1374),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1279),
.A2(n_1353),
.B(n_1325),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1295),
.A2(n_1304),
.B1(n_1299),
.B2(n_1345),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1320),
.B(n_1327),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1322),
.B(n_1313),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1322),
.B(n_1313),
.Y(n_1448)
);

AOI221xp5_ASAP7_75t_L g1449 ( 
.A1(n_1339),
.A2(n_1289),
.B1(n_1288),
.B2(n_1392),
.C(n_1275),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1305),
.B(n_1311),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1305),
.B(n_1311),
.Y(n_1451)
);

NAND4xp25_ASAP7_75t_L g1452 ( 
.A(n_1282),
.B(n_1354),
.C(n_1397),
.D(n_1359),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1312),
.B(n_1343),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1381),
.A2(n_1356),
.B1(n_1369),
.B2(n_1290),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1364),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1370),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_L g1457 ( 
.A(n_1381),
.B(n_1379),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1372),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1351),
.A2(n_1382),
.B(n_1276),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1279),
.B(n_1353),
.Y(n_1460)
);

AOI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1368),
.A2(n_1375),
.B1(n_1299),
.B2(n_1333),
.C(n_1323),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1333),
.B(n_1318),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1318),
.B(n_1348),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1367),
.A2(n_1350),
.B(n_1394),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1316),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1337),
.A2(n_1351),
.B(n_1382),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1295),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1349),
.B(n_1278),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1316),
.B(n_1341),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1276),
.A2(n_1360),
.B(n_1396),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1285),
.A2(n_1347),
.B(n_1361),
.C(n_1384),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1324),
.A2(n_1360),
.B1(n_1387),
.B2(n_1298),
.Y(n_1473)
);

AOI221x1_ASAP7_75t_SL g1474 ( 
.A1(n_1316),
.A2(n_1374),
.B1(n_1280),
.B2(n_1376),
.C(n_1385),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1316),
.A2(n_896),
.B(n_1256),
.C(n_1239),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1386),
.B(n_1374),
.Y(n_1476)
);

AOI221x1_ASAP7_75t_SL g1477 ( 
.A1(n_1281),
.A2(n_626),
.B1(n_1239),
.B2(n_1256),
.C(n_896),
.Y(n_1477)
);

O2A1O1Ixp5_ASAP7_75t_L g1478 ( 
.A1(n_1355),
.A2(n_1123),
.B(n_1380),
.C(n_1127),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1389),
.B(n_1396),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1308),
.B(n_1317),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1308),
.B(n_1317),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1304),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1328),
.A2(n_1306),
.B(n_1292),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1391),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1366),
.A2(n_947),
.B1(n_896),
.B2(n_1156),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1366),
.A2(n_947),
.B1(n_896),
.B2(n_1156),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1308),
.B(n_1317),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1300),
.Y(n_1488)
);

AOI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1281),
.A2(n_896),
.B1(n_1256),
.B2(n_1239),
.C(n_1123),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1294),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1476),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1476),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1470),
.B(n_1466),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1437),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1425),
.B(n_1409),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1418),
.Y(n_1496)
);

BUFx4f_ASAP7_75t_SL g1497 ( 
.A(n_1442),
.Y(n_1497)
);

AOI322xp5_ASAP7_75t_L g1498 ( 
.A1(n_1489),
.A2(n_1404),
.A3(n_1406),
.B1(n_1461),
.B2(n_1449),
.C1(n_1477),
.C2(n_1428),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1428),
.B(n_1424),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1453),
.Y(n_1500)
);

AO21x2_ASAP7_75t_L g1501 ( 
.A1(n_1444),
.A2(n_1438),
.B(n_1472),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1423),
.A2(n_1407),
.B(n_1460),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1405),
.A2(n_1403),
.B1(n_1485),
.B2(n_1486),
.Y(n_1503)
);

OR2x6_ASAP7_75t_L g1504 ( 
.A(n_1408),
.B(n_1467),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1459),
.B(n_1420),
.Y(n_1505)
);

OAI21xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1431),
.A2(n_1443),
.B(n_1432),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1435),
.A2(n_1426),
.B(n_1448),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1410),
.A2(n_1483),
.B(n_1433),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1490),
.B(n_1414),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1413),
.A2(n_1487),
.B(n_1481),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1412),
.B(n_1480),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1453),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1434),
.B(n_1411),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1436),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1412),
.B(n_1480),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1455),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1465),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1429),
.B(n_1421),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1456),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1481),
.B(n_1487),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1458),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1410),
.A2(n_1483),
.B(n_1433),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1439),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1445),
.A2(n_1452),
.B1(n_1431),
.B2(n_1473),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1439),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1454),
.A2(n_1488),
.B1(n_1416),
.B2(n_1468),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1465),
.Y(n_1527)
);

BUFx8_ASAP7_75t_L g1528 ( 
.A(n_1420),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1419),
.A2(n_1430),
.B1(n_1484),
.B2(n_1468),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1518),
.B(n_1495),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1500),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1500),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1528),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1510),
.B(n_1427),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1512),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1504),
.B(n_1469),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1510),
.B(n_1417),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1499),
.B(n_1448),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1504),
.B(n_1505),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1510),
.B(n_1415),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1518),
.B(n_1464),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1505),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1510),
.B(n_1426),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1510),
.B(n_1450),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1517),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1496),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1493),
.B(n_1446),
.Y(n_1548)
);

NOR2x1_ASAP7_75t_L g1549 ( 
.A(n_1504),
.B(n_1447),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1493),
.B(n_1446),
.Y(n_1550)
);

NAND2x1_ASAP7_75t_L g1551 ( 
.A(n_1504),
.B(n_1441),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1511),
.B(n_1422),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1495),
.B(n_1447),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1511),
.B(n_1422),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1540),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1531),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1531),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1552),
.B(n_1511),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1532),
.Y(n_1559)
);

OAI221xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1530),
.A2(n_1498),
.B1(n_1506),
.B2(n_1524),
.C(n_1504),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1548),
.B(n_1550),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1552),
.B(n_1515),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1530),
.A2(n_1503),
.B1(n_1504),
.B2(n_1506),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1540),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1542),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1546),
.A2(n_1522),
.B(n_1508),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1536),
.B(n_1503),
.C(n_1402),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

NAND2xp33_ASAP7_75t_R g1569 ( 
.A(n_1542),
.B(n_1482),
.Y(n_1569)
);

AO21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1553),
.A2(n_1524),
.B(n_1513),
.Y(n_1570)
);

OAI33xp33_ASAP7_75t_L g1571 ( 
.A1(n_1553),
.A2(n_1513),
.A3(n_1525),
.B1(n_1523),
.B2(n_1521),
.B3(n_1519),
.Y(n_1571)
);

OAI211xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1553),
.A2(n_1498),
.B(n_1529),
.C(n_1478),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1539),
.A2(n_1526),
.B1(n_1505),
.B2(n_1497),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1539),
.A2(n_1505),
.B1(n_1526),
.B2(n_1529),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1545),
.A2(n_1499),
.B1(n_1475),
.B2(n_1494),
.C(n_1519),
.Y(n_1575)
);

AO21x1_ASAP7_75t_SL g1576 ( 
.A1(n_1534),
.A2(n_1451),
.B(n_1525),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1552),
.B(n_1515),
.Y(n_1577)
);

OAI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1549),
.A2(n_1505),
.B1(n_1462),
.B2(n_1474),
.C(n_1457),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1536),
.B(n_1502),
.C(n_1494),
.Y(n_1579)
);

OAI221xp5_ASAP7_75t_L g1580 ( 
.A1(n_1549),
.A2(n_1505),
.B1(n_1442),
.B2(n_1491),
.C(n_1492),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1552),
.B(n_1515),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1520),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1535),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1535),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1547),
.Y(n_1585)
);

AO21x2_ASAP7_75t_L g1586 ( 
.A1(n_1546),
.A2(n_1527),
.B(n_1501),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1539),
.A2(n_1497),
.B1(n_1443),
.B2(n_1479),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1547),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1547),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1549),
.A2(n_1491),
.B1(n_1492),
.B2(n_1463),
.C(n_1482),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1538),
.B(n_1507),
.Y(n_1591)
);

OAI211xp5_ASAP7_75t_L g1592 ( 
.A1(n_1536),
.A2(n_1502),
.B(n_1451),
.C(n_1516),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1533),
.Y(n_1593)
);

OAI33xp33_ASAP7_75t_L g1594 ( 
.A1(n_1534),
.A2(n_1523),
.A3(n_1521),
.B1(n_1516),
.B2(n_1514),
.B3(n_1509),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1554),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1561),
.B(n_1543),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1575),
.B(n_1544),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1586),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1561),
.Y(n_1599)
);

AND2x6_ASAP7_75t_SL g1600 ( 
.A(n_1569),
.B(n_1440),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1586),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1579),
.B(n_1592),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1555),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1586),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1566),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1555),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1576),
.B(n_1545),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1591),
.B(n_1534),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1545),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1585),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1588),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1589),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1561),
.B(n_1545),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1570),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1591),
.B(n_1534),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1564),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_SL g1620 ( 
.A(n_1567),
.B(n_1544),
.C(n_1551),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1556),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1595),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1557),
.B(n_1544),
.Y(n_1623)
);

INVx4_ASAP7_75t_SL g1624 ( 
.A(n_1558),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1624),
.B(n_1562),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1610),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1560),
.C(n_1572),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1624),
.B(n_1562),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1624),
.B(n_1577),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1565),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1597),
.B(n_1565),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1617),
.B(n_1602),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1617),
.B(n_1582),
.Y(n_1633)
);

NAND2xp33_ASAP7_75t_SL g1634 ( 
.A(n_1600),
.B(n_1563),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1624),
.B(n_1577),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1622),
.B(n_1559),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1622),
.B(n_1581),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1622),
.B(n_1583),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1624),
.B(n_1581),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1603),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1624),
.B(n_1570),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1622),
.B(n_1584),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1624),
.B(n_1544),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1600),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1610),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1603),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1609),
.B(n_1612),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1609),
.B(n_1537),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1537),
.Y(n_1649)
);

NAND4xp25_ASAP7_75t_L g1650 ( 
.A(n_1620),
.B(n_1574),
.C(n_1590),
.D(n_1580),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1619),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1620),
.B(n_1593),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1623),
.B(n_1537),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1599),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1599),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1603),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1619),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1599),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1612),
.B(n_1616),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1607),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1621),
.B(n_1541),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1621),
.A2(n_1571),
.B1(n_1594),
.B2(n_1573),
.C(n_1541),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1621),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1607),
.Y(n_1664)
);

OAI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1611),
.A2(n_1578),
.B(n_1502),
.C(n_1551),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1663),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1626),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1625),
.B(n_1616),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1640),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1640),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1625),
.B(n_1596),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1613),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1646),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1625),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1632),
.B(n_1613),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1625),
.B(n_1596),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1627),
.A2(n_1539),
.B1(n_1543),
.B2(n_1587),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1627),
.B(n_1644),
.Y(n_1679)
);

XNOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1630),
.B(n_1593),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1662),
.B(n_1614),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1654),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1637),
.B(n_1611),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1641),
.B(n_1596),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1634),
.A2(n_1551),
.B(n_1539),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1646),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1650),
.B(n_1596),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1652),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1636),
.B(n_1614),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1656),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1656),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1641),
.B(n_1596),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1655),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1618),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1636),
.B(n_1618),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1639),
.Y(n_1698)
);

NOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1665),
.B(n_1638),
.Y(n_1699)
);

AOI211xp5_ASAP7_75t_L g1700 ( 
.A1(n_1658),
.A2(n_1471),
.B(n_1598),
.C(n_1601),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1638),
.B(n_1615),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1695),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1698),
.B(n_1639),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1647),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1669),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1695),
.Y(n_1706)
);

INVx3_ASAP7_75t_SL g1707 ( 
.A(n_1680),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1674),
.B(n_1647),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1679),
.A2(n_1639),
.B1(n_1539),
.B2(n_1635),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1685),
.B(n_1639),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1694),
.B(n_1628),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1671),
.B(n_1628),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1670),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1673),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1679),
.B(n_1654),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1688),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1681),
.A2(n_1635),
.B1(n_1629),
.B2(n_1643),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1683),
.Y(n_1718)
);

OR2x6_ASAP7_75t_L g1719 ( 
.A(n_1667),
.B(n_1629),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1699),
.B(n_1660),
.Y(n_1720)
);

INVx4_ASAP7_75t_L g1721 ( 
.A(n_1671),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1668),
.B(n_1659),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1692),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1666),
.Y(n_1724)
);

NAND2x1_ASAP7_75t_L g1725 ( 
.A(n_1676),
.B(n_1643),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1668),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1693),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1720),
.B(n_1690),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1724),
.Y(n_1729)
);

OAI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1707),
.A2(n_1681),
.B1(n_1696),
.B2(n_1677),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1712),
.B(n_1682),
.Y(n_1731)
);

NAND2xp33_ASAP7_75t_L g1732 ( 
.A(n_1707),
.B(n_1675),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1707),
.A2(n_1689),
.B1(n_1700),
.B2(n_1687),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1724),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1722),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1702),
.A2(n_1675),
.B1(n_1672),
.B2(n_1676),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1712),
.B(n_1659),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1715),
.B(n_1672),
.C(n_1691),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1706),
.A2(n_1701),
.B(n_1691),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1721),
.B(n_1678),
.Y(n_1740)
);

NAND2x1_ASAP7_75t_L g1741 ( 
.A(n_1719),
.B(n_1701),
.Y(n_1741)
);

NAND2x1_ASAP7_75t_L g1742 ( 
.A(n_1719),
.B(n_1697),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1722),
.B(n_1686),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1718),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1726),
.B(n_1684),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1719),
.B(n_1653),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1717),
.A2(n_1664),
.B1(n_1660),
.B2(n_1649),
.C(n_1648),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1732),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1728),
.A2(n_1719),
.B1(n_1709),
.B2(n_1721),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1730),
.A2(n_1722),
.B1(n_1711),
.B2(n_1721),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1742),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1729),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1734),
.B(n_1726),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1735),
.B(n_1704),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1736),
.B(n_1704),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1744),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1736),
.B(n_1708),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1731),
.B(n_1711),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1758),
.B(n_1740),
.Y(n_1759)
);

AOI221xp5_ASAP7_75t_L g1760 ( 
.A1(n_1748),
.A2(n_1739),
.B1(n_1733),
.B2(n_1738),
.C(n_1741),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1750),
.A2(n_1748),
.B1(n_1728),
.B2(n_1751),
.C(n_1749),
.Y(n_1761)
);

NOR2x1_ASAP7_75t_L g1762 ( 
.A(n_1752),
.B(n_1728),
.Y(n_1762)
);

AOI211xp5_ASAP7_75t_L g1763 ( 
.A1(n_1755),
.A2(n_1743),
.B(n_1745),
.C(n_1747),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1754),
.Y(n_1764)
);

AOI222xp33_ASAP7_75t_L g1765 ( 
.A1(n_1757),
.A2(n_1716),
.B1(n_1713),
.B2(n_1714),
.C1(n_1705),
.C2(n_1727),
.Y(n_1765)
);

NAND3xp33_ASAP7_75t_SL g1766 ( 
.A(n_1753),
.B(n_1746),
.C(n_1725),
.Y(n_1766)
);

AOI21xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1756),
.A2(n_1713),
.B(n_1705),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1764),
.B(n_1737),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1759),
.B(n_1708),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1762),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1760),
.A2(n_1703),
.B(n_1722),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1767),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1768),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1770),
.B(n_1763),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1772),
.B(n_1765),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1769),
.Y(n_1776)
);

INVx3_ASAP7_75t_L g1777 ( 
.A(n_1771),
.Y(n_1777)
);

NOR3xp33_ASAP7_75t_L g1778 ( 
.A(n_1770),
.B(n_1761),
.C(n_1766),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1773),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1778),
.B(n_1714),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1777),
.Y(n_1781)
);

AOI222xp33_ASAP7_75t_L g1782 ( 
.A1(n_1774),
.A2(n_1727),
.B1(n_1716),
.B2(n_1723),
.C1(n_1703),
.C2(n_1710),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1775),
.B(n_1723),
.Y(n_1783)
);

NOR2xp67_ASAP7_75t_L g1784 ( 
.A(n_1779),
.B(n_1776),
.Y(n_1784)
);

AND4x1_ASAP7_75t_L g1785 ( 
.A(n_1783),
.B(n_1710),
.C(n_1725),
.D(n_1648),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1780),
.B(n_1703),
.C(n_1664),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1785),
.Y(n_1787)
);

INVx4_ASAP7_75t_L g1788 ( 
.A(n_1787),
.Y(n_1788)
);

AOI22x1_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1781),
.B1(n_1782),
.B2(n_1784),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1788),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1790),
.B(n_1786),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1789),
.A2(n_1703),
.B1(n_1657),
.B2(n_1651),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1791),
.A2(n_1651),
.B1(n_1657),
.B2(n_1661),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1792),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1604),
.B1(n_1598),
.B2(n_1601),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1793),
.Y(n_1796)
);

AO22x1_ASAP7_75t_L g1797 ( 
.A1(n_1796),
.A2(n_1605),
.B1(n_1606),
.B2(n_1608),
.Y(n_1797)
);

OR2x6_ASAP7_75t_L g1798 ( 
.A(n_1797),
.B(n_1795),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1604),
.B1(n_1598),
.B2(n_1601),
.Y(n_1799)
);

AO22x1_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1606),
.B1(n_1608),
.B2(n_1605),
.Y(n_1800)
);

AOI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1604),
.B(n_1598),
.C(n_1601),
.Y(n_1801)
);


endmodule