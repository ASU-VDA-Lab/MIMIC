module fake_netlist_1_7407_n_23 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_23;
wire n_20;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
NAND2xp33_ASAP7_75t_R g10 ( .A(n_2), .B(n_5), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_7), .B(n_5), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
O2A1O1Ixp33_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_1), .B(n_2), .C(n_3), .Y(n_16) );
AO21x1_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_13), .B(n_10), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_18), .B(n_14), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g20 ( .A(n_19), .B(n_12), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_13), .B(n_15), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_4), .B1(n_8), .B2(n_9), .Y(n_23) );
endmodule