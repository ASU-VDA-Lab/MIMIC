module fake_netlist_5_339_n_1911 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1911);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1911;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_315;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1817;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g173 ( 
.A(n_65),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_46),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_51),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_84),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_16),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_19),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_32),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_23),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_88),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_90),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_45),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_140),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_124),
.Y(n_193)
);

INVxp33_ASAP7_75t_SL g194 ( 
.A(n_95),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_17),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

CKINVDCx11_ASAP7_75t_R g198 ( 
.A(n_17),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_117),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_56),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_66),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_37),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_39),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_85),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_60),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_42),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_51),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_21),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_47),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_104),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_49),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_91),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_110),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_48),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_46),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_7),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_74),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_31),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_41),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_49),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_36),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_75),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_144),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_13),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_148),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_25),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_64),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_129),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_93),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_44),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_162),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_61),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_5),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_133),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_161),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_18),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_116),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_19),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_52),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_79),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_10),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_23),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_128),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_149),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_153),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_145),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_62),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_97),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_31),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_154),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_34),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_96),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_5),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_35),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_99),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_143),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_102),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_165),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_120),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_100),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_82),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_24),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_136),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_26),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_138),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_10),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_43),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_9),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_172),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_53),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_32),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_103),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_156),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_141),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_4),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_35),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_52),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_168),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_29),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_107),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_98),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_2),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_105),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_1),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_3),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_86),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_25),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_26),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_41),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_24),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_6),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_56),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_57),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_63),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_130),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_123),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_7),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_59),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_164),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_6),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_118),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_4),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_142),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_14),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_115),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_147),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_89),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_12),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_69),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_27),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_59),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_114),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_87),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_36),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_22),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_159),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_131),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_43),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_167),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_47),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_18),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_111),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_53),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_77),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_108),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_28),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_8),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_29),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_15),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_70),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_173),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_173),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_177),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_198),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_174),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_190),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_226),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_295),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_177),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_329),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_179),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_313),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_181),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_179),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_192),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_183),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_192),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_323),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_205),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_183),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_174),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_184),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_251),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_331),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_336),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_186),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_295),
.B(n_0),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_205),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_251),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_196),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_189),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_271),
.B(n_0),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_175),
.B(n_3),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_202),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_207),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_207),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_215),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_215),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_203),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_199),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_333),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_R g387 ( 
.A(n_176),
.B(n_121),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_208),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_209),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_231),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_231),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_233),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_210),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_211),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_233),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_234),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_212),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_217),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_221),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_194),
.B(n_9),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_234),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_213),
.B(n_11),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_222),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_238),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_235),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_223),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_235),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_248),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_248),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_237),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_227),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_252),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_213),
.B(n_13),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_304),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_228),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_252),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_232),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_178),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_180),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_182),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_246),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_191),
.B(n_14),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_296),
.B(n_15),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_311),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_250),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_261),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_185),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_311),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_314),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_R g432 ( 
.A(n_357),
.B(n_187),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_419),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_428),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_351),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_345),
.B(n_322),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_428),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_356),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_413),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_420),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_428),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_428),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_421),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_428),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_R g450 ( 
.A(n_357),
.B(n_188),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_366),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_403),
.B(n_344),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_366),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_346),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_425),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_371),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_371),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_349),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_347),
.B(n_322),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_349),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g462 ( 
.A(n_414),
.B(n_296),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_430),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_365),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_365),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_376),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_429),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_350),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_353),
.B(n_249),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_367),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_355),
.B(n_193),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_377),
.B(n_242),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_362),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_358),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_359),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_376),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_378),
.B(n_307),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_379),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_361),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_363),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_379),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_373),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_380),
.Y(n_486)
);

NOR2x1_ASAP7_75t_L g487 ( 
.A(n_423),
.B(n_191),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_372),
.B(n_300),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_381),
.B(n_249),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_352),
.A2(n_260),
.B1(n_280),
.B2(n_283),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_382),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_401),
.B(n_300),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_368),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_378),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_390),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_395),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_384),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_384),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_406),
.B(n_204),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_408),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_409),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_470),
.B(n_410),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_475),
.B(n_254),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_434),
.Y(n_511)
);

AND3x2_ASAP7_75t_L g512 ( 
.A(n_475),
.B(n_254),
.C(n_360),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_477),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_452),
.B(n_411),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_452),
.B(n_404),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_259),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_388),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_488),
.B(n_185),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_388),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_478),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_L g524 ( 
.A(n_487),
.B(n_201),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_470),
.B(n_490),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_442),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_488),
.B(n_389),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_472),
.B(n_185),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_489),
.B(n_389),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

INVx11_ASAP7_75t_L g533 ( 
.A(n_446),
.Y(n_533)
);

INVx5_ASAP7_75t_L g534 ( 
.A(n_463),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_451),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_453),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_455),
.B(n_230),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_489),
.A2(n_386),
.B1(n_385),
.B2(n_375),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_478),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_486),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_496),
.B(n_393),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_496),
.B(n_405),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_472),
.B(n_393),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_470),
.B(n_364),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_498),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_432),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_496),
.B(n_394),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_440),
.B(n_415),
.C(n_469),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_503),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_185),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_490),
.B(n_259),
.Y(n_552)
);

BUFx4f_ASAP7_75t_L g553 ( 
.A(n_478),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_505),
.B(n_394),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_478),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_440),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_455),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_485),
.B(n_185),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_453),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_506),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_478),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_480),
.B(n_370),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_483),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_483),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_490),
.B(n_272),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_485),
.B(n_397),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_469),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_478),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_437),
.B(n_272),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_485),
.B(n_197),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_453),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_453),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_437),
.B(n_273),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_436),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_480),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_485),
.B(n_197),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_480),
.A2(n_398),
.B1(n_307),
.B2(n_424),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_397),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_450),
.B(n_197),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_445),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_460),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_445),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_483),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_450),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_462),
.A2(n_460),
.B1(n_502),
.B2(n_500),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_445),
.B(n_399),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_507),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_460),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_507),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_507),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_445),
.B(n_399),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_507),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_507),
.Y(n_597)
);

AO22x2_ASAP7_75t_L g598 ( 
.A1(n_491),
.A2(n_241),
.B1(n_244),
.B2(n_263),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_507),
.B(n_400),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_507),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_454),
.B(n_400),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_491),
.A2(n_247),
.B1(n_305),
.B2(n_328),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_463),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_435),
.B(n_273),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_482),
.B(n_197),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_482),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

NOR2x1p5_ASAP7_75t_L g608 ( 
.A(n_457),
.B(n_348),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_435),
.B(n_407),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_435),
.B(n_276),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_438),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_458),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_467),
.B(n_407),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_492),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_456),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_439),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_462),
.A2(n_314),
.B1(n_340),
.B2(n_342),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_476),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_492),
.Y(n_619)
);

INVx6_ASAP7_75t_L g620 ( 
.A(n_463),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_456),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_438),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_438),
.B(n_412),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_459),
.B(n_461),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_492),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_463),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_494),
.Y(n_627)
);

AO21x2_ASAP7_75t_L g628 ( 
.A1(n_444),
.A2(n_387),
.B(n_310),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_459),
.B(n_412),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_494),
.B(n_416),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_444),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_479),
.B(n_416),
.Y(n_632)
);

AND2x2_ASAP7_75t_SL g633 ( 
.A(n_494),
.B(n_276),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_481),
.B(n_418),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_484),
.B(n_418),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_463),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_501),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_461),
.B(n_422),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_444),
.B(n_422),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_504),
.B(n_427),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_497),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_447),
.B(n_497),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_495),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_463),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_502),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_497),
.Y(n_646)
);

AND2x2_ASAP7_75t_SL g647 ( 
.A(n_499),
.B(n_282),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_499),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_499),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_463),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_500),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_471),
.B(n_282),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_500),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_471),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_502),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_473),
.B(n_348),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_473),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_474),
.B(n_285),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_576),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_584),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_529),
.B(n_427),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_514),
.B(n_466),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_543),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_515),
.B(n_354),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_517),
.B(n_354),
.Y(n_665)
);

O2A1O1Ixp5_ASAP7_75t_L g666 ( 
.A1(n_510),
.A2(n_447),
.B(n_315),
.C(n_297),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_526),
.B(n_466),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_526),
.B(n_466),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_520),
.A2(n_369),
.B1(n_318),
.B2(n_300),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_526),
.B(n_466),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_645),
.B(n_464),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_645),
.B(n_464),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_585),
.B(n_253),
.Y(n_673)
);

OAI22x1_ASAP7_75t_L g674 ( 
.A1(n_539),
.A2(n_214),
.B1(n_342),
.B2(n_218),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_510),
.A2(n_297),
.B1(n_285),
.B2(n_315),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_651),
.B(n_464),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_655),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_584),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_592),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_585),
.B(n_293),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_547),
.B(n_588),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_576),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_651),
.B(n_464),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_523),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_625),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_625),
.B(n_464),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_649),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_531),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_544),
.A2(n_308),
.B1(n_339),
.B2(n_268),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_563),
.B(n_175),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_615),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_649),
.B(n_599),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_654),
.B(n_464),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_523),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_554),
.B(n_509),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_509),
.B(n_464),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_509),
.B(n_468),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_579),
.A2(n_317),
.B1(n_320),
.B2(n_338),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_657),
.B(n_468),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_572),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_624),
.B(n_468),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_615),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_552),
.A2(n_317),
.B1(n_320),
.B2(n_338),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_547),
.B(n_206),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_552),
.B(n_197),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_538),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_568),
.A2(n_255),
.B1(n_327),
.B2(n_326),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_624),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_588),
.B(n_216),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_621),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_624),
.B(n_468),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_582),
.A2(n_245),
.B1(n_321),
.B2(n_319),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_542),
.A2(n_243),
.B1(n_309),
.B2(n_291),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_552),
.A2(n_330),
.B1(n_468),
.B2(n_340),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_548),
.B(n_220),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_538),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_592),
.B(n_468),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_621),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_606),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_513),
.B(n_468),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_607),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_579),
.B(n_225),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_552),
.A2(n_229),
.B1(n_236),
.B2(n_239),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_552),
.A2(n_330),
.B1(n_288),
.B2(n_337),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_584),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_630),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_518),
.B(n_447),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_519),
.A2(n_583),
.B(n_530),
.C(n_551),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_557),
.B(n_474),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_602),
.B(n_302),
.C(n_266),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_532),
.B(n_240),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_614),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_557),
.Y(n_733)
);

BUFx12f_ASAP7_75t_SL g734 ( 
.A(n_601),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_619),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_627),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_629),
.B(n_256),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_521),
.B(n_465),
.Y(n_738)
);

AND2x2_ASAP7_75t_SL g739 ( 
.A(n_551),
.B(n_330),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_629),
.B(n_638),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_571),
.B(n_431),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_638),
.B(n_257),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_541),
.B(n_465),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_631),
.A2(n_465),
.B(n_449),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_523),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_546),
.B(n_433),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_633),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_641),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_550),
.B(n_433),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_646),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_552),
.A2(n_330),
.B1(n_337),
.B2(n_335),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_567),
.A2(n_258),
.B1(n_262),
.B2(n_265),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_567),
.A2(n_330),
.B1(n_335),
.B2(n_200),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_613),
.B(n_267),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_SL g756 ( 
.A(n_519),
.B(n_195),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_545),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_571),
.A2(n_195),
.B(n_325),
.C(n_324),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_511),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_633),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_632),
.B(n_275),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_559),
.B(n_441),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_537),
.B(n_269),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_648),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_634),
.B(n_277),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_653),
.Y(n_766)
);

OAI221xp5_ASAP7_75t_L g767 ( 
.A1(n_617),
.A2(n_200),
.B1(n_214),
.B2(n_218),
.C(n_219),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_567),
.B(n_270),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_537),
.B(n_274),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_564),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_567),
.A2(n_294),
.B1(n_224),
.B2(n_241),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_561),
.B(n_443),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_567),
.A2(n_294),
.B1(n_224),
.B2(n_244),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_565),
.B(n_443),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_569),
.B(n_219),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_556),
.B(n_263),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_571),
.B(n_448),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_637),
.B(n_448),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_567),
.A2(n_299),
.B1(n_281),
.B2(n_288),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_566),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_587),
.B(n_449),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_635),
.B(n_279),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_642),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_523),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_SL g785 ( 
.A(n_535),
.B(n_304),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_524),
.B(n_278),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_516),
.A2(n_301),
.B1(n_281),
.B2(n_299),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_647),
.B(n_287),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_577),
.B(n_264),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_516),
.A2(n_264),
.B1(n_301),
.B2(n_325),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_647),
.B(n_286),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_524),
.B(n_341),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_586),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_577),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_577),
.B(n_658),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_609),
.B(n_334),
.Y(n_796)
);

O2A1O1Ixp5_ASAP7_75t_L g797 ( 
.A1(n_530),
.A2(n_558),
.B(n_573),
.C(n_580),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_652),
.B(n_324),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_656),
.B(n_332),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_516),
.A2(n_304),
.B1(n_312),
.B2(n_306),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_623),
.B(n_316),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_652),
.B(n_80),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_586),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_612),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_516),
.A2(n_303),
.B1(n_298),
.B2(n_292),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_586),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_640),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_639),
.B(n_290),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_578),
.B(n_289),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_516),
.B(n_284),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_652),
.B(n_68),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_589),
.B(n_20),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_516),
.A2(n_67),
.B1(n_170),
.B2(n_169),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_590),
.B(n_171),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_595),
.B(n_163),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_658),
.B(n_157),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_611),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_611),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_658),
.B(n_155),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_581),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_583),
.B(n_27),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_611),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_558),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_643),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_622),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_616),
.Y(n_826)
);

AND2x4_ASAP7_75t_SL g827 ( 
.A(n_535),
.B(n_150),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_512),
.B(n_137),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_775),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_706),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_802),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_659),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_670),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_660),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_SL g835 ( 
.A(n_748),
.B(n_760),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_659),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_670),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_660),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_748),
.B(n_535),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_700),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_759),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_804),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_795),
.B(n_608),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_733),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_760),
.B(n_628),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_795),
.B(n_549),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_695),
.B(n_628),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_706),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_775),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_682),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_733),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_733),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_682),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_679),
.B(n_622),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_708),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_SL g856 ( 
.A(n_820),
.B(n_616),
.C(n_511),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_746),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_691),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_679),
.B(n_622),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_795),
.B(n_591),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_662),
.B(n_596),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_688),
.B(n_593),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_687),
.Y(n_863)
);

BUFx10_ASAP7_75t_L g864 ( 
.A(n_759),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_783),
.B(n_755),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_783),
.B(n_597),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_687),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_757),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_SL g869 ( 
.A(n_669),
.B(n_527),
.C(n_618),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_804),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_691),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_793),
.Y(n_872)
);

AO22x1_ASAP7_75t_L g873 ( 
.A1(n_761),
.A2(n_782),
.B1(n_765),
.B2(n_730),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_776),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_726),
.B(n_527),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_793),
.Y(n_876)
);

AND3x1_ASAP7_75t_SL g877 ( 
.A(n_767),
.B(n_598),
.C(n_33),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_716),
.B(n_525),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_660),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_803),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_716),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_802),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_812),
.A2(n_598),
.B1(n_604),
.B2(n_610),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_777),
.B(n_594),
.Y(n_884)
);

CKINVDCx20_ASAP7_75t_R g885 ( 
.A(n_734),
.Y(n_885)
);

AND2x6_ASAP7_75t_L g886 ( 
.A(n_811),
.B(n_525),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_R g887 ( 
.A(n_734),
.B(n_643),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_733),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_777),
.B(n_794),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_794),
.B(n_522),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_729),
.B(n_522),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_685),
.B(n_508),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_702),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_R g894 ( 
.A(n_785),
.B(n_533),
.Y(n_894)
);

INVxp67_ASAP7_75t_SL g895 ( 
.A(n_733),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_671),
.B(n_508),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_802),
.A2(n_598),
.B1(n_604),
.B2(n_610),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_672),
.B(n_575),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_803),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_729),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_676),
.B(n_575),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_780),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_683),
.B(n_536),
.Y(n_903)
);

CKINVDCx14_ASAP7_75t_R g904 ( 
.A(n_826),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_702),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_780),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_710),
.Y(n_907)
);

INVx6_ASAP7_75t_L g908 ( 
.A(n_729),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_824),
.Y(n_909)
);

BUFx4_ASAP7_75t_SL g910 ( 
.A(n_809),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_693),
.B(n_536),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_678),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_741),
.B(n_574),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_811),
.B(n_667),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_663),
.B(n_573),
.Y(n_915)
);

BUFx4f_ASAP7_75t_L g916 ( 
.A(n_828),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_692),
.B(n_560),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_668),
.B(n_591),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_741),
.B(n_560),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_741),
.B(n_574),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_828),
.B(n_650),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_710),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_809),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_718),
.Y(n_924)
);

INVx5_ASAP7_75t_L g925 ( 
.A(n_802),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_802),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_740),
.A2(n_580),
.B1(n_604),
.B2(n_610),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_690),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_802),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_684),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_718),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_719),
.Y(n_932)
);

AOI22x1_ASAP7_75t_L g933 ( 
.A1(n_678),
.A2(n_725),
.B1(n_806),
.B2(n_770),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_726),
.B(n_553),
.Y(n_934)
);

OAI221xp5_ASAP7_75t_L g935 ( 
.A1(n_800),
.A2(n_605),
.B1(n_644),
.B2(n_636),
.C(n_626),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_684),
.Y(n_936)
);

BUFx8_ASAP7_75t_L g937 ( 
.A(n_828),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_796),
.B(n_801),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_807),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_789),
.B(n_798),
.Y(n_940)
);

NOR3xp33_ASAP7_75t_SL g941 ( 
.A(n_820),
.B(n_605),
.C(n_34),
.Y(n_941)
);

NOR3xp33_ASAP7_75t_SL g942 ( 
.A(n_758),
.B(n_30),
.C(n_37),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_678),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_770),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_684),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_732),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_787),
.A2(n_610),
.B1(n_604),
.B2(n_636),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_732),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_664),
.B(n_650),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_735),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_735),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_661),
.B(n_644),
.C(n_626),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_677),
.Y(n_953)
);

BUFx12f_ASAP7_75t_L g954 ( 
.A(n_690),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_751),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_789),
.B(n_528),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_776),
.B(n_38),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_681),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_798),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_816),
.B(n_570),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_751),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_674),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_694),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_756),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_725),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_665),
.B(n_778),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_827),
.Y(n_967)
);

AOI211xp5_ASAP7_75t_L g968 ( 
.A1(n_799),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_788),
.B(n_528),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_764),
.Y(n_970)
);

INVx5_ASAP7_75t_L g971 ( 
.A(n_694),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_674),
.B(n_562),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_758),
.B(n_603),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_694),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_745),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_827),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_764),
.Y(n_977)
);

AND2x6_ASAP7_75t_L g978 ( 
.A(n_813),
.B(n_600),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_745),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_791),
.B(n_528),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_725),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_721),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_786),
.B(n_603),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_766),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_756),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_766),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_696),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_747),
.B(n_750),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_697),
.B(n_603),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_810),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_721),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_745),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_717),
.B(n_540),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_SL g994 ( 
.A(n_698),
.B(n_40),
.C(n_42),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_736),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_822),
.Y(n_996)
);

INVx5_ASAP7_75t_L g997 ( 
.A(n_825),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_736),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_749),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_749),
.Y(n_1000)
);

AO22x1_ASAP7_75t_L g1001 ( 
.A1(n_819),
.A2(n_610),
.B1(n_604),
.B2(n_600),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_806),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_737),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_728),
.A2(n_591),
.B(n_570),
.C(n_553),
.Y(n_1004)
);

AO22x1_ASAP7_75t_L g1005 ( 
.A1(n_814),
.A2(n_610),
.B1(n_604),
.B2(n_600),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_817),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_727),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_704),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_817),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_818),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_763),
.B(n_540),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_769),
.B(n_540),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_762),
.B(n_562),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_772),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_742),
.B(n_555),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_792),
.B(n_555),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_818),
.Y(n_1017)
);

NOR2xp67_ASAP7_75t_L g1018 ( 
.A(n_841),
.B(n_709),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_936),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_832),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_865),
.B(n_673),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_936),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_916),
.A2(n_703),
.B1(n_711),
.B2(n_701),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_941),
.A2(n_938),
.B(n_968),
.C(n_994),
.Y(n_1024)
);

NOR2x1_ASAP7_75t_SL g1025 ( 
.A(n_831),
.B(n_815),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_933),
.A2(n_797),
.B(n_686),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_832),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_916),
.A2(n_675),
.B1(n_784),
.B2(n_714),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_960),
.A2(n_699),
.B(n_720),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_829),
.B(n_715),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_831),
.B(n_743),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_930),
.A2(n_570),
.B(n_553),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_831),
.A2(n_754),
.B1(n_724),
.B2(n_752),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_988),
.B(n_680),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_930),
.A2(n_705),
.B(n_768),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_840),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_1004),
.A2(n_774),
.A3(n_781),
.B(n_738),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_928),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_923),
.B(n_808),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_887),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_849),
.B(n_857),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_930),
.A2(n_705),
.B(n_768),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_941),
.A2(n_821),
.B(n_823),
.C(n_790),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_855),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1014),
.B(n_689),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_928),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1014),
.B(n_771),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_SL g1048 ( 
.A(n_831),
.B(n_722),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_960),
.A2(n_825),
.B(n_822),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_882),
.B(n_825),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_896),
.A2(n_822),
.B(n_666),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_898),
.A2(n_744),
.B(n_779),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_882),
.A2(n_739),
.B1(n_713),
.B2(n_773),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_847),
.A2(n_753),
.B(n_723),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_930),
.A2(n_600),
.B(n_739),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_940),
.B(n_707),
.Y(n_1056)
);

BUFx2_ASAP7_75t_SL g1057 ( 
.A(n_885),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_936),
.Y(n_1058)
);

INVxp67_ASAP7_75t_SL g1059 ( 
.A(n_936),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_945),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_994),
.A2(n_805),
.B(n_712),
.C(n_731),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_901),
.A2(n_620),
.B(n_534),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_963),
.A2(n_534),
.B(n_620),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_SL g1064 ( 
.A1(n_929),
.A2(n_620),
.B(n_534),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_873),
.B(n_534),
.C(n_45),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_945),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_940),
.B(n_44),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_944),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_940),
.B(n_50),
.Y(n_1069)
);

AO21x1_ASAP7_75t_L g1070 ( 
.A1(n_914),
.A2(n_50),
.B(n_54),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_945),
.Y(n_1071)
);

OA21x2_ASAP7_75t_L g1072 ( 
.A1(n_1004),
.A2(n_534),
.B(n_92),
.Y(n_1072)
);

AO21x2_ASAP7_75t_L g1073 ( 
.A1(n_934),
.A2(n_83),
.B(n_132),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_903),
.A2(n_81),
.B(n_125),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_842),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_918),
.A2(n_76),
.B(n_122),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_932),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_874),
.B(n_54),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_SL g1079 ( 
.A1(n_897),
.A2(n_94),
.B(n_113),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_836),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_L g1081 ( 
.A1(n_962),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_917),
.A2(n_71),
.B(n_112),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_836),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_889),
.B(n_55),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_987),
.B(n_58),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_963),
.A2(n_134),
.B(n_971),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_850),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_870),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_918),
.A2(n_914),
.B(n_911),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_987),
.B(n_833),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_875),
.B(n_857),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_845),
.A2(n_980),
.A3(n_969),
.B(n_861),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_887),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_837),
.B(n_959),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_862),
.B(n_1007),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_956),
.A2(n_884),
.B(n_919),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_894),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_920),
.A2(n_866),
.B(n_949),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_868),
.B(n_939),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_934),
.A2(n_860),
.B(n_1006),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_840),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_860),
.A2(n_1017),
.B(n_1006),
.Y(n_1102)
);

AO32x2_ASAP7_75t_L g1103 ( 
.A1(n_851),
.A2(n_852),
.A3(n_877),
.B1(n_856),
.B2(n_979),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_892),
.A2(n_989),
.B(n_935),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_856),
.A2(n_948),
.B(n_984),
.C(n_950),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_868),
.B(n_953),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_953),
.B(n_954),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_946),
.B(n_951),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_989),
.A2(n_993),
.B(n_927),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_955),
.B(n_961),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_945),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1005),
.A2(n_1001),
.B(n_890),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_882),
.A2(n_925),
.B1(n_926),
.B2(n_929),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1009),
.A2(n_1017),
.B(n_1010),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_915),
.B(n_954),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_909),
.Y(n_1116)
);

NOR2xp67_ASAP7_75t_SL g1117 ( 
.A(n_971),
.B(n_925),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_910),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_L g1119 ( 
.A(n_1008),
.B(n_958),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_970),
.B(n_977),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_885),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_986),
.B(n_966),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_863),
.B(n_867),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1009),
.A2(n_1010),
.B(n_872),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_850),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_925),
.B(n_926),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_990),
.B(n_982),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_869),
.B(n_1003),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_982),
.B(n_991),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_830),
.Y(n_1130)
);

BUFx4f_ASAP7_75t_SL g1131 ( 
.A(n_864),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_991),
.B(n_998),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_904),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_876),
.A2(n_880),
.B(n_899),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1013),
.A2(n_993),
.B(n_975),
.Y(n_1135)
);

AO21x1_ASAP7_75t_L g1136 ( 
.A1(n_835),
.A2(n_973),
.B(n_839),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_926),
.B(n_974),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_998),
.A2(n_999),
.A3(n_995),
.B(n_1000),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_843),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_853),
.A2(n_931),
.B(n_924),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_957),
.A2(n_942),
.B(n_835),
.C(n_883),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_974),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_839),
.B(n_843),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_974),
.A2(n_992),
.B(n_975),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_976),
.B(n_900),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_853),
.Y(n_1146)
);

BUFx4_ASAP7_75t_SL g1147 ( 
.A(n_830),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_858),
.A2(n_931),
.B(n_924),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_926),
.B(n_992),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_900),
.B(n_895),
.Y(n_1150)
);

AOI221x1_ASAP7_75t_L g1151 ( 
.A1(n_952),
.A2(n_973),
.B1(n_902),
.B2(n_906),
.C(n_983),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_858),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_992),
.A2(n_844),
.B(n_997),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_997),
.A2(n_979),
.B(n_1015),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_921),
.B(n_878),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_997),
.A2(n_983),
.B(n_1012),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_848),
.Y(n_1157)
);

AOI221x1_ASAP7_75t_L g1158 ( 
.A1(n_973),
.A2(n_983),
.B1(n_1012),
.B2(n_1011),
.C(n_1016),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1002),
.A2(n_905),
.A3(n_893),
.B(n_907),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_921),
.B(n_878),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_908),
.B(n_985),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_997),
.A2(n_1012),
.B(n_1011),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_891),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_871),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_871),
.A2(n_907),
.B(n_905),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1011),
.A2(n_859),
.B(n_854),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_883),
.A2(n_913),
.B(n_893),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_922),
.Y(n_1168)
);

OAI21xp33_ASAP7_75t_SL g1169 ( 
.A1(n_897),
.A2(n_972),
.B(n_838),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_1119),
.B(n_843),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1104),
.A2(n_1016),
.B(n_922),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1036),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1024),
.A2(n_964),
.B(n_904),
.C(n_846),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1128),
.A2(n_846),
.B1(n_908),
.B2(n_921),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1128),
.A2(n_894),
.B1(n_937),
.B2(n_846),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1034),
.B(n_1095),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1091),
.B(n_864),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1138),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1138),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1159),
.Y(n_1180)
);

AO21x2_ASAP7_75t_L g1181 ( 
.A1(n_1054),
.A2(n_1016),
.B(n_891),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1021),
.B(n_881),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1062),
.A2(n_1098),
.B(n_1026),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1045),
.A2(n_908),
.B1(n_848),
.B2(n_881),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1138),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1036),
.Y(n_1186)
);

INVx8_ASAP7_75t_L g1187 ( 
.A(n_1022),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1049),
.A2(n_834),
.B(n_838),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1099),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1122),
.B(n_972),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1126),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1106),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1022),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1090),
.B(n_891),
.Y(n_1194)
);

OR2x6_ASAP7_75t_L g1195 ( 
.A(n_1109),
.B(n_972),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1163),
.B(n_913),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1100),
.Y(n_1197)
);

AO21x2_ASAP7_75t_L g1198 ( 
.A1(n_1026),
.A2(n_942),
.B(n_878),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1116),
.B(n_967),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1040),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1151),
.A2(n_947),
.B(n_913),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1088),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1143),
.B(n_888),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1100),
.A2(n_1114),
.B(n_1124),
.Y(n_1204)
);

AOI22x1_ASAP7_75t_L g1205 ( 
.A1(n_1166),
.A2(n_834),
.B1(n_981),
.B2(n_965),
.Y(n_1205)
);

INVx4_ASAP7_75t_SL g1206 ( 
.A(n_1066),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1138),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1024),
.B(n_886),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1159),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1159),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_1075),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_1066),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1159),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1126),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1020),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1114),
.A2(n_943),
.B(n_981),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1105),
.A2(n_978),
.B(n_886),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1061),
.A2(n_965),
.B(n_943),
.C(n_912),
.Y(n_1218)
);

NOR2x1_ASAP7_75t_SL g1219 ( 
.A(n_1073),
.B(n_1031),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1061),
.A2(n_886),
.B(n_978),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1112),
.A2(n_1136),
.B(n_1031),
.Y(n_1221)
);

BUFx4f_ASAP7_75t_L g1222 ( 
.A(n_1066),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1129),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1027),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1089),
.A2(n_1029),
.B(n_1035),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1030),
.A2(n_1039),
.B1(n_1163),
.B2(n_1065),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1161),
.A2(n_888),
.B1(n_851),
.B2(n_852),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1167),
.B(n_879),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1050),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1127),
.B(n_886),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1043),
.A2(n_978),
.B(n_947),
.Y(n_1231)
);

OAI221xp5_ASAP7_75t_L g1232 ( 
.A1(n_1039),
.A2(n_877),
.B1(n_879),
.B2(n_912),
.C(n_937),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1027),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_1131),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1022),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1158),
.A2(n_978),
.A3(n_996),
.B(n_967),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1141),
.B(n_996),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1161),
.B(n_996),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1124),
.A2(n_978),
.B(n_996),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1080),
.Y(n_1240)
);

BUFx8_ASAP7_75t_L g1241 ( 
.A(n_1038),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1147),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1097),
.Y(n_1243)
);

OA21x2_ASAP7_75t_L g1244 ( 
.A1(n_1089),
.A2(n_1029),
.B(n_1074),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_SL g1245 ( 
.A1(n_1070),
.A2(n_1025),
.B(n_1048),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1108),
.B(n_1110),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1044),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1141),
.B(n_1077),
.Y(n_1248)
);

AO21x2_ASAP7_75t_L g1249 ( 
.A1(n_1105),
.A2(n_1096),
.B(n_1042),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1156),
.A2(n_1162),
.B(n_1135),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1148),
.A2(n_1165),
.B(n_1102),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1148),
.A2(n_1165),
.B(n_1102),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1120),
.B(n_1085),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1132),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1080),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1032),
.A2(n_1144),
.B(n_1055),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1088),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1130),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1130),
.B(n_1157),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1140),
.A2(n_1051),
.B(n_1076),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1051),
.A2(n_1076),
.B(n_1134),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1074),
.A2(n_1052),
.B(n_1134),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1043),
.A2(n_1053),
.B(n_1047),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1083),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1154),
.A2(n_1052),
.B(n_1063),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_L g1266 ( 
.A(n_1067),
.B(n_1069),
.C(n_1115),
.Y(n_1266)
);

INVx3_ASAP7_75t_SL g1267 ( 
.A(n_1097),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1056),
.A2(n_1131),
.B1(n_1093),
.B2(n_1018),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1086),
.A2(n_1072),
.B(n_1113),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1072),
.A2(n_1153),
.B(n_1137),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_L g1271 ( 
.A(n_1093),
.B(n_1101),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1157),
.B(n_1145),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1155),
.B(n_1160),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1041),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1041),
.B(n_1094),
.Y(n_1275)
);

AOI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1072),
.A2(n_1023),
.B(n_1082),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1083),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1084),
.A2(n_1164),
.B(n_1152),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1117),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1168),
.A2(n_1087),
.B(n_1125),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1087),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1125),
.B(n_1146),
.Y(n_1282)
);

AO21x2_ASAP7_75t_L g1283 ( 
.A1(n_1079),
.A2(n_1028),
.B(n_1149),
.Y(n_1283)
);

AO21x1_ASAP7_75t_L g1284 ( 
.A1(n_1033),
.A2(n_1149),
.B(n_1137),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1115),
.A2(n_1107),
.B1(n_1078),
.B2(n_1081),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1050),
.A2(n_1064),
.B(n_1146),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1123),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1082),
.A2(n_1150),
.B(n_1071),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1073),
.A2(n_1037),
.B(n_1092),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1037),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1037),
.A2(n_1092),
.B(n_1082),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1046),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1133),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1066),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1058),
.A2(n_1142),
.B(n_1060),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1169),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1121),
.B(n_1092),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1059),
.A2(n_1111),
.B(n_1071),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1019),
.A2(n_1060),
.B1(n_1057),
.B2(n_1103),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1092),
.B(n_1019),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1037),
.A2(n_1103),
.B(n_1139),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1103),
.B(n_1139),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_SL g1303 ( 
.A1(n_1103),
.A2(n_1118),
.B(n_1139),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1117),
.B(n_831),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1136),
.A2(n_1070),
.B(n_1109),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1038),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_R g1307 ( 
.A(n_1097),
.B(n_643),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1034),
.B(n_940),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1068),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1126),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1021),
.B(n_688),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1034),
.B(n_940),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1100),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1021),
.A2(n_785),
.B1(n_759),
.B2(n_928),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1100),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1128),
.A2(n_869),
.B1(n_517),
.B2(n_520),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1100),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1100),
.Y(n_1318)
);

AOI221x1_ASAP7_75t_L g1319 ( 
.A1(n_1105),
.A2(n_1024),
.B1(n_1104),
.B2(n_1065),
.C(n_1141),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1117),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1068),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1100),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1147),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1128),
.A2(n_869),
.B1(n_517),
.B2(n_520),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1100),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1151),
.A2(n_1026),
.B(n_1062),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1151),
.A2(n_1026),
.B(n_1062),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1311),
.B(n_1176),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1173),
.B(n_1195),
.Y(n_1329)
);

OAI221xp5_ASAP7_75t_L g1330 ( 
.A1(n_1316),
.A2(n_1324),
.B1(n_1285),
.B2(n_1266),
.C(n_1226),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1187),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1308),
.B(n_1312),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1263),
.A2(n_1231),
.B1(n_1195),
.B2(n_1308),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1280),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1314),
.A2(n_1312),
.B1(n_1268),
.B2(n_1200),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1195),
.A2(n_1176),
.B1(n_1253),
.B2(n_1220),
.Y(n_1336)
);

NAND3xp33_ASAP7_75t_L g1337 ( 
.A(n_1319),
.B(n_1174),
.C(n_1232),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_SL g1338 ( 
.A(n_1175),
.B(n_1246),
.C(n_1190),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1272),
.B(n_1192),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1200),
.A2(n_1170),
.B1(n_1177),
.B2(n_1184),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1247),
.Y(n_1341)
);

AOI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1190),
.A2(n_1297),
.B(n_1208),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1319),
.A2(n_1275),
.B1(n_1287),
.B2(n_1195),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1287),
.A2(n_1274),
.B1(n_1189),
.B2(n_1182),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1309),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1248),
.A2(n_1296),
.B1(n_1297),
.B2(n_1305),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1187),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1272),
.B(n_1196),
.Y(n_1348)
);

NAND2xp33_ASAP7_75t_R g1349 ( 
.A(n_1201),
.B(n_1307),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1296),
.B(n_1238),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1235),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1276),
.A2(n_1305),
.B(n_1245),
.Y(n_1352)
);

INVx4_ASAP7_75t_L g1353 ( 
.A(n_1187),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1242),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1321),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1259),
.B(n_1272),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1259),
.B(n_1258),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1276),
.A2(n_1245),
.B(n_1256),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1211),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1194),
.B(n_1273),
.Y(n_1360)
);

NAND2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1235),
.B(n_1193),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1259),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1199),
.A2(n_1172),
.B1(n_1271),
.B2(n_1293),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1258),
.Y(n_1364)
);

INVx6_ASAP7_75t_L g1365 ( 
.A(n_1187),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1248),
.A2(n_1217),
.B1(n_1284),
.B2(n_1273),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1273),
.B(n_1223),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1235),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1201),
.A2(n_1171),
.B1(n_1181),
.B2(n_1217),
.Y(n_1369)
);

AOI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1186),
.A2(n_1218),
.B1(n_1228),
.B2(n_1299),
.C(n_1284),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1202),
.A2(n_1230),
.B(n_1186),
.C(n_1300),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1257),
.B(n_1202),
.Y(n_1372)
);

NAND2xp33_ASAP7_75t_SL g1373 ( 
.A(n_1235),
.B(n_1193),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1204),
.A2(n_1251),
.B(n_1252),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1193),
.Y(n_1375)
);

OR2x6_ASAP7_75t_L g1376 ( 
.A(n_1237),
.B(n_1298),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1196),
.B(n_1257),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1237),
.B(n_1267),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1223),
.B(n_1254),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_R g1380 ( 
.A(n_1201),
.B(n_1203),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1292),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1267),
.A2(n_1243),
.B1(n_1320),
.B2(n_1279),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1280),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1215),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1243),
.A2(n_1292),
.B1(n_1254),
.B2(n_1234),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_L g1386 ( 
.A(n_1235),
.B(n_1304),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1212),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1215),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1201),
.A2(n_1217),
.B1(n_1198),
.B2(n_1302),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1222),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1212),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1306),
.Y(n_1392)
);

INVx4_ASAP7_75t_L g1393 ( 
.A(n_1212),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1282),
.B(n_1203),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1222),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1198),
.A2(n_1283),
.B1(n_1303),
.B2(n_1249),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1241),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1280),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1224),
.B(n_1233),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1233),
.B(n_1240),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1240),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1255),
.B(n_1264),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1206),
.B(n_1294),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1255),
.B(n_1264),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1277),
.B(n_1281),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1222),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1277),
.B(n_1281),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1278),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1278),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1212),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1283),
.A2(n_1249),
.B1(n_1198),
.B2(n_1278),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1178),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1241),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_SL g1414 ( 
.A(n_1234),
.B(n_1227),
.C(n_1242),
.Y(n_1414)
);

BUFx12f_ASAP7_75t_L g1415 ( 
.A(n_1323),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1241),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1323),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1212),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1206),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1294),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1304),
.A2(n_1221),
.B1(n_1278),
.B2(n_1214),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1191),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1178),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1304),
.A2(n_1221),
.B1(n_1214),
.B2(n_1310),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1283),
.A2(n_1250),
.B1(n_1249),
.B2(n_1191),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1191),
.A2(n_1214),
.B1(n_1310),
.B2(n_1229),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1250),
.A2(n_1205),
.B(n_1239),
.Y(n_1427)
);

BUFx4f_ASAP7_75t_L g1428 ( 
.A(n_1310),
.Y(n_1428)
);

NAND2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1229),
.B(n_1290),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1206),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1229),
.B(n_1295),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1179),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1180),
.Y(n_1433)
);

OAI211xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1290),
.A2(n_1179),
.B(n_1207),
.C(n_1185),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1303),
.A2(n_1185),
.B1(n_1207),
.B2(n_1289),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1225),
.A2(n_1265),
.B(n_1269),
.Y(n_1436)
);

CKINVDCx6p67_ASAP7_75t_R g1437 ( 
.A(n_1209),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1289),
.A2(n_1210),
.B1(n_1205),
.B2(n_1180),
.Y(n_1438)
);

OAI221xp5_ASAP7_75t_L g1439 ( 
.A1(n_1262),
.A2(n_1225),
.B1(n_1244),
.B2(n_1210),
.C(n_1291),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1213),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1236),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1213),
.A2(n_1291),
.B1(n_1327),
.B2(n_1326),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1239),
.A2(n_1301),
.B(n_1288),
.C(n_1269),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1262),
.B(n_1244),
.C(n_1291),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1236),
.B(n_1250),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1288),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1236),
.B(n_1301),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1204),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1219),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1236),
.B(n_1289),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1291),
.A2(n_1183),
.B1(n_1262),
.B2(n_1327),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1219),
.A2(n_1236),
.B1(n_1326),
.B2(n_1327),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1262),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1244),
.B(n_1188),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1188),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1265),
.A2(n_1183),
.B(n_1270),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1216),
.Y(n_1457)
);

NAND2x1_ASAP7_75t_L g1458 ( 
.A(n_1244),
.B(n_1327),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1286),
.B(n_1326),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1286),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1260),
.A2(n_1261),
.B(n_1197),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1261),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1356),
.B(n_1313),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1330),
.A2(n_1326),
.B1(n_1315),
.B2(n_1317),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1412),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1364),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1338),
.A2(n_1318),
.B1(n_1322),
.B2(n_1325),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1423),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1343),
.A2(n_1318),
.B1(n_1322),
.B2(n_1325),
.C(n_1337),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1367),
.B(n_1360),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1335),
.A2(n_1340),
.B1(n_1378),
.B2(n_1336),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1432),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1379),
.B(n_1344),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1338),
.A2(n_1329),
.B1(n_1336),
.B2(n_1333),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1357),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_L g1476 ( 
.A(n_1364),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1329),
.A2(n_1333),
.B1(n_1414),
.B2(n_1332),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1339),
.B(n_1348),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1378),
.A2(n_1363),
.B1(n_1419),
.B2(n_1385),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1343),
.A2(n_1342),
.B1(n_1370),
.B2(n_1371),
.C(n_1350),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1390),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1414),
.A2(n_1332),
.B1(n_1376),
.B2(n_1350),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1419),
.A2(n_1346),
.B1(n_1376),
.B2(n_1382),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1356),
.A2(n_1362),
.B1(n_1359),
.B2(n_1377),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1357),
.B(n_1394),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1346),
.A2(n_1413),
.B1(n_1416),
.B2(n_1397),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1366),
.A2(n_1392),
.B1(n_1381),
.B2(n_1437),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1428),
.A2(n_1381),
.B1(n_1420),
.B2(n_1406),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1428),
.A2(n_1406),
.B1(n_1395),
.B2(n_1449),
.Y(n_1489)
);

OAI33xp33_ASAP7_75t_L g1490 ( 
.A1(n_1341),
.A2(n_1355),
.A3(n_1345),
.B1(n_1434),
.B2(n_1421),
.B3(n_1442),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1395),
.A2(n_1372),
.B1(n_1430),
.B2(n_1365),
.Y(n_1491)
);

OAI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1417),
.A2(n_1425),
.B1(n_1349),
.B2(n_1396),
.C(n_1361),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1372),
.A2(n_1430),
.B1(n_1365),
.B2(n_1390),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1411),
.A2(n_1396),
.B1(n_1369),
.B2(n_1445),
.C(n_1435),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1415),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1422),
.A2(n_1352),
.B1(n_1431),
.B2(n_1441),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1422),
.A2(n_1352),
.B1(n_1431),
.B2(n_1441),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1369),
.A2(n_1429),
.B1(n_1386),
.B2(n_1361),
.Y(n_1498)
);

AOI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1411),
.A2(n_1435),
.B1(n_1434),
.B2(n_1438),
.C(n_1389),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1430),
.A2(n_1365),
.B1(n_1455),
.B2(n_1353),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1447),
.A2(n_1380),
.B1(n_1450),
.B2(n_1410),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1399),
.B(n_1404),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1424),
.A2(n_1426),
.B(n_1373),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1443),
.A2(n_1444),
.B(n_1451),
.Y(n_1504)
);

NOR3xp33_ASAP7_75t_L g1505 ( 
.A(n_1373),
.B(n_1331),
.C(n_1347),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1354),
.B(n_1368),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1440),
.Y(n_1507)
);

AO221x2_ASAP7_75t_L g1508 ( 
.A1(n_1446),
.A2(n_1409),
.B1(n_1408),
.B2(n_1401),
.C(n_1388),
.Y(n_1508)
);

CKINVDCx11_ASAP7_75t_R g1509 ( 
.A(n_1351),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1402),
.B(n_1407),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1353),
.A2(n_1331),
.B1(n_1347),
.B2(n_1368),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1410),
.A2(n_1418),
.B1(n_1391),
.B2(n_1387),
.Y(n_1512)
);

OAI211xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1438),
.A2(n_1389),
.B(n_1452),
.C(n_1384),
.Y(n_1513)
);

AOI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1429),
.A2(n_1439),
.B1(n_1452),
.B2(n_1405),
.C(n_1400),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1403),
.A2(n_1358),
.B1(n_1351),
.B2(n_1375),
.Y(n_1515)
);

BUFx5_ASAP7_75t_L g1516 ( 
.A(n_1462),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1403),
.A2(n_1358),
.B1(n_1351),
.B2(n_1375),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1387),
.A2(n_1391),
.B1(n_1393),
.B2(n_1418),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1410),
.A2(n_1418),
.B1(n_1393),
.B2(n_1460),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1410),
.A2(n_1418),
.B1(n_1433),
.B2(n_1459),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1460),
.Y(n_1521)
);

AOI221xp5_ASAP7_75t_L g1522 ( 
.A1(n_1451),
.A2(n_1433),
.B1(n_1457),
.B2(n_1453),
.C(n_1454),
.Y(n_1522)
);

NAND2xp33_ASAP7_75t_R g1523 ( 
.A(n_1374),
.B(n_1448),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1458),
.A2(n_1374),
.B1(n_1383),
.B2(n_1398),
.C(n_1436),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1374),
.A2(n_1316),
.B1(n_1324),
.B2(n_669),
.Y(n_1525)
);

BUFx4f_ASAP7_75t_SL g1526 ( 
.A(n_1461),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1461),
.A2(n_1158),
.B(n_1231),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1390),
.Y(n_1528)
);

AOI222xp33_ASAP7_75t_L g1529 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_488),
.B2(n_493),
.C1(n_520),
.C2(n_517),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1334),
.Y(n_1531)
);

AO221x2_ASAP7_75t_L g1532 ( 
.A1(n_1337),
.A2(n_1081),
.B1(n_873),
.B2(n_1314),
.C(n_1343),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1330),
.A2(n_785),
.B1(n_1231),
.B2(n_1263),
.Y(n_1533)
);

NAND4xp25_ASAP7_75t_L g1534 ( 
.A(n_1328),
.B(n_669),
.C(n_1311),
.D(n_1316),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1328),
.B(n_1176),
.Y(n_1537)
);

NAND4xp25_ASAP7_75t_L g1538 ( 
.A(n_1328),
.B(n_669),
.C(n_1311),
.D(n_1316),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1412),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1354),
.Y(n_1540)
);

BUFx4f_ASAP7_75t_SL g1541 ( 
.A(n_1415),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1542)
);

CKINVDCx11_ASAP7_75t_R g1543 ( 
.A(n_1392),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1330),
.A2(n_1324),
.B1(n_1316),
.B2(n_669),
.C(n_520),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1334),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1330),
.A2(n_1328),
.B1(n_1231),
.B2(n_785),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1427),
.A2(n_1443),
.B(n_1456),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1330),
.A2(n_1328),
.B1(n_1231),
.B2(n_785),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1330),
.A2(n_1316),
.B1(n_1324),
.B2(n_869),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1348),
.B(n_1377),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1364),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1412),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1381),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_1324),
.B2(n_1316),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1412),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1328),
.B(n_578),
.Y(n_1559)
);

AOI222xp33_ASAP7_75t_L g1560 ( 
.A1(n_1330),
.A2(n_869),
.B1(n_488),
.B2(n_493),
.C1(n_520),
.C2(n_517),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1356),
.B(n_1339),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1334),
.Y(n_1562)
);

OAI211xp5_ASAP7_75t_L g1563 ( 
.A1(n_1330),
.A2(n_669),
.B(n_1324),
.C(n_1316),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1354),
.Y(n_1564)
);

OAI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1330),
.A2(n_1324),
.B1(n_1316),
.B2(n_669),
.C(n_520),
.Y(n_1565)
);

NOR2x1_ASAP7_75t_L g1566 ( 
.A(n_1328),
.B(n_1266),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1501),
.B(n_1504),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1463),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1545),
.B(n_1562),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1473),
.B(n_1470),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1544),
.A2(n_1565),
.B1(n_1533),
.B2(n_1560),
.Y(n_1573)
);

AO31x2_ASAP7_75t_L g1574 ( 
.A1(n_1525),
.A2(n_1520),
.A3(n_1558),
.B(n_1539),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1547),
.B(n_1494),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1547),
.B(n_1508),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1508),
.B(n_1516),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1533),
.A2(n_1529),
.B1(n_1549),
.B2(n_1542),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1465),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1468),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1472),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1521),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1507),
.B(n_1554),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1530),
.A2(n_1557),
.B1(n_1535),
.B2(n_1536),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1524),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1526),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1469),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1527),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1551),
.B(n_1550),
.C(n_1555),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1499),
.B(n_1464),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1563),
.B(n_1546),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1522),
.B(n_1496),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1523),
.Y(n_1593)
);

BUFx2_ASAP7_75t_SL g1594 ( 
.A(n_1500),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1513),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1467),
.B(n_1503),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1497),
.B(n_1480),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1474),
.B(n_1514),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1502),
.B(n_1510),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1492),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1515),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1498),
.B(n_1482),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1566),
.B(n_1548),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1563),
.A2(n_1546),
.B1(n_1548),
.B2(n_1534),
.C(n_1538),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1485),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1532),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1517),
.B(n_1532),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1477),
.B(n_1471),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_L g1609 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1559),
.B(n_1487),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1519),
.Y(n_1611)
);

OAI211xp5_ASAP7_75t_L g1612 ( 
.A1(n_1486),
.A2(n_1479),
.B(n_1484),
.C(n_1519),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1589),
.A2(n_1490),
.B1(n_1478),
.B2(n_1552),
.C(n_1488),
.Y(n_1614)
);

AO21x2_ASAP7_75t_L g1615 ( 
.A1(n_1587),
.A2(n_1505),
.B(n_1512),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1582),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1568),
.B(n_1561),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1589),
.A2(n_1505),
.B(n_1489),
.Y(n_1619)
);

NAND2x1_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1466),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1572),
.B(n_1556),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1578),
.A2(n_1573),
.B1(n_1584),
.B2(n_1608),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1583),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1580),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_R g1625 ( 
.A(n_1568),
.B(n_1564),
.Y(n_1625)
);

OAI33xp33_ASAP7_75t_L g1626 ( 
.A1(n_1584),
.A2(n_1491),
.A3(n_1493),
.B1(n_1511),
.B2(n_1518),
.B3(n_1490),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1570),
.B(n_1466),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1573),
.A2(n_1561),
.B1(n_1475),
.B2(n_1495),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1593),
.B(n_1466),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1604),
.A2(n_1506),
.B1(n_1553),
.B2(n_1476),
.C(n_1528),
.Y(n_1630)
);

NAND2xp33_ASAP7_75t_SL g1631 ( 
.A(n_1598),
.B(n_1476),
.Y(n_1631)
);

INVxp67_ASAP7_75t_SL g1632 ( 
.A(n_1567),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1604),
.B(n_1476),
.C(n_1553),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1578),
.A2(n_1543),
.B1(n_1541),
.B2(n_1553),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1568),
.B(n_1528),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1581),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1572),
.B(n_1540),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1579),
.B(n_1481),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1581),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1591),
.A2(n_1481),
.B1(n_1509),
.B2(n_1598),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1568),
.B(n_1481),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1583),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1581),
.Y(n_1643)
);

OAI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1608),
.A2(n_1600),
.B1(n_1595),
.B2(n_1591),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1599),
.Y(n_1645)
);

OR2x6_ASAP7_75t_L g1646 ( 
.A(n_1594),
.B(n_1588),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1569),
.B(n_1605),
.Y(n_1647)
);

OAI33xp33_ASAP7_75t_L g1648 ( 
.A1(n_1587),
.A2(n_1595),
.A3(n_1600),
.B1(n_1603),
.B2(n_1579),
.B3(n_1610),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1598),
.A2(n_1600),
.B1(n_1595),
.B2(n_1609),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1587),
.B(n_1603),
.C(n_1597),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1598),
.A2(n_1597),
.B1(n_1612),
.B2(n_1610),
.C(n_1590),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1569),
.B(n_1605),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1569),
.B(n_1605),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1612),
.B(n_1597),
.C(n_1590),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1609),
.A2(n_1606),
.B1(n_1590),
.B2(n_1597),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1569),
.B(n_1605),
.Y(n_1656)
);

INVx4_ASAP7_75t_L g1657 ( 
.A(n_1586),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_R g1658 ( 
.A(n_1582),
.B(n_1601),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1582),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1618),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1613),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1623),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1613),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1636),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1636),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1647),
.B(n_1576),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1643),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1643),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1647),
.B(n_1576),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1652),
.B(n_1593),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1657),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1652),
.B(n_1585),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1653),
.B(n_1576),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1653),
.B(n_1576),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1656),
.B(n_1575),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1656),
.B(n_1575),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1632),
.B(n_1585),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1645),
.B(n_1585),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1629),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1624),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1635),
.B(n_1575),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1620),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1642),
.B(n_1585),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1629),
.B(n_1571),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1617),
.B(n_1641),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1617),
.B(n_1641),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1624),
.B(n_1583),
.Y(n_1687)
);

OR2x6_ASAP7_75t_L g1688 ( 
.A(n_1646),
.B(n_1594),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_1583),
.Y(n_1689)
);

AND2x4_ASAP7_75t_SL g1690 ( 
.A(n_1646),
.B(n_1657),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1620),
.B(n_1575),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1657),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1627),
.B(n_1577),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1679),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1682),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1661),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1660),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1660),
.Y(n_1698)
);

INVxp67_ASAP7_75t_SL g1699 ( 
.A(n_1677),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1684),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1682),
.B(n_1627),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1672),
.B(n_1574),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1677),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1679),
.B(n_1621),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1672),
.B(n_1638),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1681),
.B(n_1684),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1691),
.A2(n_1654),
.B1(n_1622),
.B2(n_1596),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1661),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1627),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1660),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1663),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1670),
.B(n_1574),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1680),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1663),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.B(n_1574),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1678),
.B(n_1582),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1664),
.Y(n_1717)
);

NOR2x1p5_ASAP7_75t_SL g1718 ( 
.A(n_1680),
.B(n_1588),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1664),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1682),
.B(n_1570),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1675),
.B(n_1588),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1681),
.B(n_1616),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1665),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1678),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1682),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1667),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1688),
.A2(n_1651),
.B(n_1648),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1675),
.B(n_1588),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1667),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1668),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1687),
.B(n_1574),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1681),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1707),
.B(n_1650),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1716),
.B(n_1637),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1697),
.Y(n_1736)
);

AOI32xp33_ASAP7_75t_L g1737 ( 
.A1(n_1694),
.A2(n_1655),
.A3(n_1644),
.B1(n_1649),
.B2(n_1590),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1703),
.B(n_1699),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1705),
.B(n_1676),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1701),
.B(n_1685),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1704),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1725),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1722),
.B(n_1659),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1695),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1697),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1700),
.B(n_1676),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1696),
.Y(n_1747)
);

AOI31xp67_ASAP7_75t_SL g1748 ( 
.A1(n_1706),
.A2(n_1619),
.A3(n_1625),
.B(n_1633),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1701),
.B(n_1685),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1701),
.B(n_1709),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1698),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1695),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1702),
.B(n_1634),
.C(n_1630),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1709),
.B(n_1685),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1702),
.B(n_1658),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1726),
.Y(n_1756)
);

AOI21xp33_ASAP7_75t_L g1757 ( 
.A1(n_1726),
.A2(n_1688),
.B(n_1601),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1698),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1676),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1720),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1721),
.B(n_1686),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1711),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1710),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1696),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1708),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1720),
.Y(n_1766)
);

INVxp67_ASAP7_75t_SL g1767 ( 
.A(n_1708),
.Y(n_1767)
);

NAND4xp25_ASAP7_75t_L g1768 ( 
.A(n_1732),
.B(n_1614),
.C(n_1609),
.D(n_1628),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_L g1769 ( 
.A(n_1712),
.B(n_1606),
.C(n_1602),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1729),
.B(n_1686),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1712),
.B(n_1687),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1715),
.B(n_1689),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1729),
.B(n_1686),
.Y(n_1773)
);

NOR2xp67_ASAP7_75t_L g1774 ( 
.A(n_1715),
.B(n_1732),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1719),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1750),
.B(n_1720),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1775),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1756),
.Y(n_1778)
);

NOR2x1_ASAP7_75t_L g1779 ( 
.A(n_1753),
.B(n_1659),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1750),
.B(n_1693),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1740),
.B(n_1693),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1741),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1737),
.B(n_1666),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1767),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1747),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1747),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1737),
.B(n_1666),
.Y(n_1787)
);

BUFx2_ASAP7_75t_L g1788 ( 
.A(n_1756),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1740),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1764),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1749),
.B(n_1693),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1764),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1765),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1734),
.B(n_1666),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1753),
.B(n_1631),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1744),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1765),
.Y(n_1797)
);

AO22x1_ASAP7_75t_L g1798 ( 
.A1(n_1748),
.A2(n_1606),
.B1(n_1691),
.B2(n_1671),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1775),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1748),
.A2(n_1733),
.B1(n_1606),
.B2(n_1769),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1762),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1768),
.A2(n_1631),
.B1(n_1596),
.B2(n_1607),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1749),
.B(n_1669),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1736),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1736),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1742),
.B(n_1669),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1768),
.A2(n_1626),
.B(n_1688),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1745),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1735),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1766),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1738),
.B(n_1691),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1779),
.B(n_1769),
.C(n_1748),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1795),
.A2(n_1757),
.B(n_1755),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1778),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1785),
.Y(n_1815)
);

NAND2x1_ASAP7_75t_SL g1816 ( 
.A(n_1802),
.B(n_1774),
.Y(n_1816)
);

CKINVDCx16_ASAP7_75t_R g1817 ( 
.A(n_1782),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1796),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1778),
.Y(n_1819)
);

NOR3xp33_ASAP7_75t_SL g1820 ( 
.A(n_1800),
.B(n_1743),
.C(n_1746),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1798),
.A2(n_1688),
.B1(n_1596),
.B2(n_1607),
.Y(n_1821)
);

AOI32xp33_ASAP7_75t_L g1822 ( 
.A1(n_1783),
.A2(n_1766),
.A3(n_1752),
.B1(n_1754),
.B2(n_1760),
.Y(n_1822)
);

OAI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1787),
.A2(n_1688),
.B1(n_1646),
.B2(n_1774),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1807),
.A2(n_1688),
.B1(n_1646),
.B2(n_1640),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1788),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1776),
.B(n_1754),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1798),
.A2(n_1596),
.B1(n_1607),
.B2(n_1602),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1785),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1789),
.A2(n_1596),
.B1(n_1602),
.B2(n_1592),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1809),
.A2(n_1596),
.B1(n_1611),
.B2(n_1760),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1784),
.B(n_1739),
.Y(n_1831)
);

OAI22xp33_ASAP7_75t_SL g1832 ( 
.A1(n_1796),
.A2(n_1752),
.B1(n_1772),
.B2(n_1771),
.Y(n_1832)
);

NAND2x1p5_ASAP7_75t_L g1833 ( 
.A(n_1788),
.B(n_1671),
.Y(n_1833)
);

NAND2x1_ASAP7_75t_L g1834 ( 
.A(n_1776),
.B(n_1745),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1780),
.Y(n_1835)
);

INVx2_ASAP7_75t_SL g1836 ( 
.A(n_1789),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1801),
.A2(n_1758),
.B1(n_1751),
.B2(n_1763),
.C(n_1772),
.Y(n_1837)
);

NOR3xp33_ASAP7_75t_SL g1838 ( 
.A(n_1817),
.B(n_1801),
.C(n_1784),
.Y(n_1838)
);

AOI221x1_ASAP7_75t_SL g1839 ( 
.A1(n_1812),
.A2(n_1797),
.B1(n_1777),
.B2(n_1792),
.C(n_1790),
.Y(n_1839)
);

NOR4xp25_ASAP7_75t_SL g1840 ( 
.A(n_1837),
.B(n_1811),
.C(n_1793),
.D(n_1786),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1818),
.B(n_1810),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1826),
.B(n_1780),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1812),
.A2(n_1794),
.B(n_1806),
.Y(n_1843)
);

XNOR2xp5_ASAP7_75t_L g1844 ( 
.A(n_1820),
.B(n_1824),
.Y(n_1844)
);

OAI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1827),
.A2(n_1813),
.B1(n_1821),
.B2(n_1814),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1814),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1819),
.B(n_1803),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1832),
.B(n_1781),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1834),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1825),
.Y(n_1850)
);

OAI21xp33_ASAP7_75t_L g1851 ( 
.A1(n_1816),
.A2(n_1799),
.B(n_1792),
.Y(n_1851)
);

CKINVDCx14_ASAP7_75t_R g1852 ( 
.A(n_1830),
.Y(n_1852)
);

AND2x2_ASAP7_75t_SL g1853 ( 
.A(n_1829),
.B(n_1786),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1815),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1831),
.B(n_1761),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1833),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1828),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1850),
.Y(n_1858)
);

NOR3xp33_ASAP7_75t_L g1859 ( 
.A(n_1841),
.B(n_1813),
.C(n_1831),
.Y(n_1859)
);

OAI221xp5_ASAP7_75t_L g1860 ( 
.A1(n_1838),
.A2(n_1822),
.B1(n_1836),
.B2(n_1833),
.C(n_1835),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1838),
.B(n_1803),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1842),
.B(n_1781),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1856),
.Y(n_1863)
);

O2A1O1Ixp5_ASAP7_75t_L g1864 ( 
.A1(n_1848),
.A2(n_1823),
.B(n_1808),
.C(n_1805),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1847),
.B(n_1770),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1846),
.B(n_1791),
.Y(n_1866)
);

OAI211xp5_ASAP7_75t_L g1867 ( 
.A1(n_1840),
.A2(n_1799),
.B(n_1793),
.C(n_1790),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1850),
.B(n_1791),
.Y(n_1868)
);

AOI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1845),
.A2(n_1805),
.B(n_1804),
.C(n_1808),
.Y(n_1869)
);

OAI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1867),
.A2(n_1851),
.B(n_1852),
.C(n_1843),
.Y(n_1870)
);

OAI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1860),
.A2(n_1839),
.B1(n_1844),
.B2(n_1849),
.C(n_1855),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1863),
.B(n_1854),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1863),
.B(n_1857),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1858),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1859),
.A2(n_1845),
.B1(n_1853),
.B2(n_1804),
.Y(n_1875)
);

AOI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1869),
.A2(n_1853),
.B(n_1771),
.C(n_1758),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1861),
.A2(n_1759),
.B1(n_1773),
.B2(n_1690),
.Y(n_1877)
);

OAI321xp33_ASAP7_75t_L g1878 ( 
.A1(n_1866),
.A2(n_1586),
.A3(n_1611),
.B1(n_1601),
.B2(n_1763),
.C(n_1751),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1864),
.A2(n_1710),
.B(n_1713),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1868),
.A2(n_1713),
.B(n_1719),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1870),
.A2(n_1862),
.B1(n_1865),
.B2(n_1671),
.Y(n_1881)
);

NAND2x1p5_ASAP7_75t_L g1882 ( 
.A(n_1872),
.B(n_1671),
.Y(n_1882)
);

AOI21xp33_ASAP7_75t_L g1883 ( 
.A1(n_1875),
.A2(n_1692),
.B(n_1615),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1874),
.B(n_1669),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1871),
.A2(n_1690),
.B(n_1586),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1873),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1882),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1886),
.B(n_1876),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1884),
.Y(n_1889)
);

INVx5_ASAP7_75t_L g1890 ( 
.A(n_1885),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1881),
.Y(n_1891)
);

XNOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1883),
.B(n_1877),
.Y(n_1892)
);

NOR2x1_ASAP7_75t_L g1893 ( 
.A(n_1888),
.B(n_1879),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1891),
.A2(n_1880),
.B1(n_1878),
.B2(n_1615),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1887),
.Y(n_1895)
);

OAI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1890),
.A2(n_1692),
.B(n_1611),
.C(n_1683),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1892),
.A2(n_1890),
.B1(n_1889),
.B2(n_1690),
.Y(n_1897)
);

CKINVDCx20_ASAP7_75t_R g1898 ( 
.A(n_1897),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1893),
.Y(n_1899)
);

CKINVDCx16_ASAP7_75t_R g1900 ( 
.A(n_1895),
.Y(n_1900)
);

BUFx4f_ASAP7_75t_SL g1901 ( 
.A(n_1898),
.Y(n_1901)
);

OAI22x1_ASAP7_75t_L g1902 ( 
.A1(n_1901),
.A2(n_1890),
.B1(n_1899),
.B2(n_1900),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1902),
.Y(n_1903)
);

NOR2xp67_ASAP7_75t_L g1904 ( 
.A(n_1902),
.B(n_1896),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1903),
.A2(n_1894),
.B1(n_1731),
.B2(n_1730),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1904),
.B(n_1731),
.Y(n_1906)
);

AOI222xp33_ASAP7_75t_SL g1907 ( 
.A1(n_1906),
.A2(n_1730),
.B1(n_1727),
.B2(n_1724),
.C1(n_1723),
.C2(n_1714),
.Y(n_1907)
);

AOI222xp33_ASAP7_75t_L g1908 ( 
.A1(n_1905),
.A2(n_1727),
.B1(n_1724),
.B2(n_1717),
.C1(n_1718),
.C2(n_1674),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1662),
.B1(n_1615),
.B2(n_1594),
.Y(n_1909)
);

AOI221xp5_ASAP7_75t_L g1910 ( 
.A1(n_1909),
.A2(n_1907),
.B1(n_1662),
.B2(n_1674),
.C(n_1673),
.Y(n_1910)
);

AOI211xp5_ASAP7_75t_L g1911 ( 
.A1(n_1910),
.A2(n_1683),
.B(n_1673),
.C(n_1674),
.Y(n_1911)
);


endmodule