module fake_aes_12436_n_712 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_712);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_712;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g93 ( .A(n_26), .Y(n_93) );
BUFx10_ASAP7_75t_L g94 ( .A(n_62), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_86), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_74), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_19), .Y(n_97) );
BUFx10_ASAP7_75t_L g98 ( .A(n_50), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_15), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_29), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_11), .Y(n_101) );
BUFx2_ASAP7_75t_SL g102 ( .A(n_11), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_81), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_45), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_34), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_88), .B(n_47), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_57), .Y(n_107) );
BUFx5_ASAP7_75t_L g108 ( .A(n_58), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_54), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_64), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_12), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_39), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_19), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_77), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_85), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_40), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_82), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_80), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_53), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_48), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_73), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_75), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_25), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_91), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_65), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_69), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_37), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_23), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_4), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_0), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_104), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_119), .B(n_1), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_119), .B(n_2), .Y(n_137) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_101), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_108), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_111), .B(n_3), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_103), .B(n_49), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_130), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_127), .B(n_5), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_130), .B(n_6), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_97), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_103), .A2(n_51), .B(n_90), .Y(n_151) );
INVxp33_ASAP7_75t_SL g152 ( .A(n_144), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_141), .B(n_100), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_137), .B(n_93), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_141), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_134), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_134), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_144), .Y(n_158) );
OAI22x1_ASAP7_75t_L g159 ( .A1(n_133), .A2(n_112), .B1(n_129), .B2(n_96), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_139), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_137), .B(n_105), .Y(n_161) );
OR2x6_ASAP7_75t_L g162 ( .A(n_138), .B(n_102), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_139), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
OAI22xp33_ASAP7_75t_L g165 ( .A1(n_135), .A2(n_101), .B1(n_114), .B2(n_131), .Y(n_165) );
NAND3xp33_ASAP7_75t_L g166 ( .A(n_148), .B(n_117), .C(n_120), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_148), .A2(n_107), .B1(n_109), .B2(n_121), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_150), .B(n_125), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_132), .B(n_94), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_147), .B(n_94), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_140), .A2(n_98), .B1(n_95), .B2(n_116), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_154), .B(n_147), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_162), .B(n_143), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_154), .B(n_141), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_161), .B(n_115), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_161), .B(n_110), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_159), .A2(n_95), .B1(n_118), .B2(n_116), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_176), .B(n_151), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_176), .B(n_151), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_152), .B(n_98), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_178), .B(n_126), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_166), .B(n_128), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_166), .B(n_124), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_171), .B(n_123), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_160), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_177), .B(n_118), .Y(n_201) );
INVx4_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_158), .B(n_106), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_183), .B(n_122), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_153), .A2(n_122), .B(n_46), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_164), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
INVx1_ASAP7_75t_SL g209 ( .A(n_164), .Y(n_209) );
NOR3xp33_ASAP7_75t_L g210 ( .A(n_165), .B(n_6), .C(n_7), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_7), .B(n_8), .C(n_9), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_155), .B(n_122), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_180), .B(n_122), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_182), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_155), .B(n_52), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_180), .B(n_8), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_167), .B(n_170), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_167), .B(n_9), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_159), .B(n_10), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_170), .Y(n_223) );
NOR2x1_ASAP7_75t_L g224 ( .A(n_209), .B(n_162), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_218), .Y(n_225) );
BUFx2_ASAP7_75t_L g226 ( .A(n_209), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_184), .B(n_159), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_219), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_191), .A2(n_162), .B(n_173), .C(n_174), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_191), .B(n_181), .Y(n_231) );
BUFx8_ASAP7_75t_L g232 ( .A(n_207), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_207), .B(n_179), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_193), .A2(n_182), .B(n_183), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_189), .B(n_179), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_200), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_185), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_193), .A2(n_182), .B(n_183), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_202), .B(n_183), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_199), .B(n_155), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_185), .B(n_169), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_211), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_194), .A2(n_182), .B(n_169), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_211), .B(n_174), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_210), .A2(n_162), .B1(n_173), .B2(n_172), .Y(n_245) );
AND2x6_ASAP7_75t_L g246 ( .A(n_216), .B(n_168), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_202), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_223), .B(n_203), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_223), .B(n_175), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_202), .B(n_168), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_185), .A2(n_162), .B1(n_182), .B2(n_168), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_194), .A2(n_182), .B(n_169), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_186), .A2(n_216), .B(n_204), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_220), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_187), .Y(n_255) );
AOI21xp5_ASAP7_75t_SL g256 ( .A1(n_216), .A2(n_217), .B(n_186), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_228), .A2(n_213), .B(n_222), .C(n_215), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_226), .B(n_185), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_243), .A2(n_205), .B(n_214), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_SL g260 ( .A1(n_252), .A2(n_198), .B(n_197), .C(n_188), .Y(n_260) );
AO21x1_ASAP7_75t_L g261 ( .A1(n_251), .A2(n_222), .B(n_221), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_231), .B(n_185), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_234), .A2(n_221), .B(n_190), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_238), .A2(n_187), .B(n_212), .C(n_208), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_253), .A2(n_212), .B(n_208), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_232), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_232), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_254), .A2(n_225), .B(n_236), .C(n_242), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_233), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_240), .A2(n_190), .B(n_206), .Y(n_270) );
AO31x2_ASAP7_75t_L g271 ( .A1(n_229), .A2(n_163), .A3(n_175), .B(n_188), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_230), .A2(n_206), .B(n_157), .C(n_172), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_216), .B(n_172), .Y(n_273) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_244), .A2(n_163), .B(n_175), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_232), .Y(n_275) );
AO31x2_ASAP7_75t_L g276 ( .A1(n_227), .A2(n_163), .A3(n_196), .B(n_201), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_248), .A2(n_172), .B(n_192), .C(n_195), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_235), .A2(n_192), .B1(n_216), .B2(n_162), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_278), .A2(n_245), .B1(n_237), .B2(n_240), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_275), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_273), .A2(n_250), .B(n_239), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_274), .Y(n_283) );
NAND3xp33_ASAP7_75t_L g284 ( .A(n_277), .B(n_245), .C(n_249), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_261), .A2(n_255), .B(n_250), .Y(n_285) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_272), .A2(n_239), .B(n_255), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
AOI21x1_ASAP7_75t_L g288 ( .A1(n_274), .A2(n_241), .B(n_246), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_267), .Y(n_289) );
OR2x6_ASAP7_75t_L g290 ( .A(n_258), .B(n_241), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_260), .A2(n_241), .B(n_247), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_269), .B(n_258), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_274), .Y(n_293) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_272), .A2(n_246), .B(n_247), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_257), .A2(n_246), .B(n_12), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_271), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_266), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_271), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_271), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_260), .A2(n_246), .B(n_59), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_283), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_283), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_283), .B(n_276), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_293), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_293), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_293), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_297), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_295), .A2(n_264), .B(n_268), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_290), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_299), .B(n_276), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_299), .B(n_276), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_297), .B(n_276), .Y(n_315) );
OR2x6_ASAP7_75t_L g316 ( .A(n_295), .B(n_279), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_297), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_284), .B(n_262), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_284), .A2(n_257), .B(n_277), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_300), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_300), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_300), .B(n_302), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_302), .B(n_270), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_292), .B(n_268), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_288), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_292), .B(n_265), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
AO21x2_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_264), .B(n_263), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_292), .B(n_259), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_290), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_285), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_285), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_313), .B(n_280), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_304), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_313), .B(n_280), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_313), .B(n_292), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_307), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_308), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_317), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_322), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_317), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_296), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_320), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_298), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_320), .Y(n_360) );
AND2x6_ASAP7_75t_L g361 ( .A(n_331), .B(n_287), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_321), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_321), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_311), .B(n_289), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_323), .B(n_298), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_319), .A2(n_301), .B(n_291), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_323), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_312), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_314), .B(n_305), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_314), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_314), .B(n_296), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_315), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_305), .B(n_294), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_328), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_315), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_305), .B(n_294), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_319), .B(n_286), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_315), .B(n_281), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_318), .B(n_287), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_330), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_312), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_330), .B(n_294), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_311), .B(n_287), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_318), .B(n_286), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_331), .A2(n_287), .B1(n_290), .B2(n_286), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_330), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_331), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_312), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_327), .B(n_286), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_312), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_369), .B(n_311), .Y(n_392) );
INVx4_ASAP7_75t_L g393 ( .A(n_361), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_380), .A2(n_331), .B1(n_386), .B2(n_336), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_342), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_369), .B(n_325), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_374), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_355), .B(n_316), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_374), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_374), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_355), .B(n_327), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_380), .B(n_327), .Y(n_403) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_337), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_386), .B(n_370), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_342), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_350), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_370), .B(n_335), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_359), .B(n_325), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_372), .B(n_375), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_343), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_343), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_351), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_378), .B(n_316), .Y(n_414) );
BUFx2_ASAP7_75t_L g415 ( .A(n_340), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_372), .B(n_335), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_378), .B(n_316), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_350), .Y(n_418) );
AND2x2_ASAP7_75t_SL g419 ( .A(n_339), .B(n_312), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_375), .B(n_334), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_368), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_390), .B(n_333), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_388), .B(n_326), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_351), .Y(n_424) );
NAND2x1_ASAP7_75t_L g425 ( .A(n_361), .B(n_326), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_390), .B(n_333), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_359), .B(n_316), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_365), .Y(n_428) );
INVx2_ASAP7_75t_SL g429 ( .A(n_340), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_364), .B(n_371), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_388), .B(n_326), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_352), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_373), .B(n_333), .Y(n_433) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_354), .B(n_316), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_350), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_337), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_339), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_340), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_353), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_356), .B(n_316), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_353), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_371), .B(n_316), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_373), .B(n_332), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_345), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_349), .B(n_332), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_376), .B(n_332), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_376), .B(n_328), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_353), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_357), .B(n_324), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_358), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_358), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_360), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_349), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_362), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_345), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_382), .B(n_360), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_348), .B(n_328), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_357), .B(n_324), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_336), .B(n_310), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_382), .B(n_326), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_360), .B(n_326), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_362), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_345), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_367), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_363), .B(n_310), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_338), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_363), .B(n_310), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_367), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_387), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_338), .B(n_291), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_348), .B(n_310), .Y(n_471) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_393), .B(n_425), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_410), .B(n_387), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_402), .B(n_388), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_428), .B(n_379), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_395), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_393), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_470), .A2(n_381), .B(n_310), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_392), .B(n_379), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_410), .B(n_384), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_403), .B(n_338), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_395), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_393), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_406), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_403), .B(n_363), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_405), .B(n_456), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_429), .B(n_389), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_405), .B(n_384), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_411), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_420), .B(n_377), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_429), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_456), .B(n_347), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_398), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_420), .B(n_377), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_436), .B(n_385), .C(n_383), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_412), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_397), .B(n_347), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_413), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_469), .B(n_344), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_457), .B(n_341), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_430), .B(n_346), .Y(n_501) );
INVxp33_ASAP7_75t_L g502 ( .A(n_425), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_469), .B(n_344), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_413), .Y(n_504) );
NAND2x1_ASAP7_75t_L g505 ( .A(n_434), .B(n_361), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_457), .B(n_341), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_424), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_424), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_440), .A2(n_381), .B(n_361), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_398), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_422), .B(n_346), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_400), .Y(n_512) );
OAI21xp33_ASAP7_75t_L g513 ( .A1(n_419), .A2(n_391), .B(n_389), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_449), .B(n_346), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_432), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_458), .B(n_344), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_400), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_422), .B(n_426), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_432), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_415), .B(n_391), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_401), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_464), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_426), .B(n_433), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_464), .Y(n_524) );
AND2x4_ASAP7_75t_SL g525 ( .A(n_437), .B(n_341), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_414), .B(n_391), .Y(n_526) );
OA211x2_ASAP7_75t_L g527 ( .A1(n_455), .A2(n_361), .B(n_389), .C(n_391), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_414), .B(n_389), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_433), .B(n_368), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_468), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_401), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_468), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_407), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_443), .B(n_446), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_407), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_415), .B(n_368), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_423), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_443), .B(n_368), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_417), .B(n_366), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_459), .B(n_366), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_446), .B(n_368), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_450), .B(n_366), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_451), .B(n_366), .Y(n_543) );
NOR2x1_ASAP7_75t_R g544 ( .A(n_438), .B(n_361), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_447), .B(n_361), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_417), .B(n_396), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_454), .B(n_361), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_462), .B(n_329), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_418), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_444), .B(n_329), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_418), .Y(n_551) );
AND3x1_ASAP7_75t_L g552 ( .A(n_394), .B(n_10), .C(n_13), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_435), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_435), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_408), .B(n_329), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_463), .B(n_329), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_473), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_492), .B(n_408), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_473), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_546), .B(n_409), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_490), .B(n_416), .Y(n_561) );
AOI21xp33_ASAP7_75t_SL g562 ( .A1(n_483), .A2(n_419), .B(n_399), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_518), .B(n_460), .Y(n_563) );
NOR4xp25_ASAP7_75t_L g564 ( .A(n_495), .B(n_399), .C(n_404), .D(n_427), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_500), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_501), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_525), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_486), .B(n_416), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_534), .B(n_453), .Y(n_569) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_540), .A2(n_442), .B(n_460), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_523), .B(n_463), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_497), .B(n_427), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_480), .B(n_445), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_474), .B(n_423), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_476), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_525), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_490), .B(n_465), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_482), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_484), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g580 ( .A1(n_540), .A2(n_471), .B(n_466), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_491), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_505), .A2(n_544), .B(n_509), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_494), .B(n_467), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_506), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_489), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_502), .A2(n_471), .B(n_431), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_481), .B(n_431), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_511), .Y(n_588) );
NOR2x1p5_ASAP7_75t_L g589 ( .A(n_477), .B(n_431), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_480), .B(n_445), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_552), .A2(n_461), .B1(n_467), .B2(n_465), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_494), .B(n_452), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_452), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_488), .B(n_448), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_485), .B(n_461), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_475), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_497), .B(n_479), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_514), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_545), .B(n_448), .Y(n_599) );
NOR2x2_ASAP7_75t_L g600 ( .A(n_527), .B(n_290), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_477), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_529), .B(n_441), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_516), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_538), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_537), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_496), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_472), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_498), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_509), .A2(n_441), .B1(n_439), .B2(n_290), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_504), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_542), .B(n_439), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_507), .Y(n_612) );
OR2x6_ASAP7_75t_L g613 ( .A(n_513), .B(n_421), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_539), .A2(n_421), .B1(n_329), .B2(n_282), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_510), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g616 ( .A(n_537), .B(n_421), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_541), .B(n_282), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_502), .A2(n_13), .B(n_14), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_508), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_515), .B(n_14), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_542), .B(n_16), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_557), .B(n_519), .Y(n_622) );
AOI322xp5_ASAP7_75t_L g623 ( .A1(n_597), .A2(n_555), .A3(n_556), .B1(n_530), .B2(n_532), .C1(n_524), .C2(n_522), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_564), .A2(n_547), .B(n_543), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_574), .B(n_520), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_581), .B(n_526), .Y(n_626) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_565), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_591), .A2(n_520), .B1(n_547), .B2(n_528), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_564), .A2(n_478), .B1(n_543), .B2(n_555), .C(n_499), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_592), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_570), .A2(n_478), .B(n_550), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_580), .A2(n_503), .B(n_499), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_592), .Y(n_633) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_586), .A2(n_503), .B(n_548), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_562), .A2(n_487), .B1(n_536), .B2(n_549), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_593), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_581), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_594), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_618), .A2(n_553), .B1(n_548), .B2(n_533), .C1(n_551), .C2(n_554), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_573), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_590), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_596), .B(n_487), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_607), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_559), .B(n_551), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_582), .B(n_536), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_575), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g647 ( .A1(n_621), .A2(n_533), .B1(n_535), .B2(n_521), .C1(n_517), .C2(n_531), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_578), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_586), .A2(n_521), .B(n_517), .C(n_512), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_609), .A2(n_600), .B(n_601), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_609), .A2(n_493), .B(n_17), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_579), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_584), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_587), .B(n_16), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_572), .A2(n_246), .B1(n_18), .B2(n_17), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_585), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_560), .A2(n_18), .A3(n_20), .B1(n_21), .B2(n_22), .C1(n_24), .C2(n_27), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_588), .Y(n_658) );
NOR4xp25_ASAP7_75t_L g659 ( .A(n_643), .B(n_621), .C(n_620), .D(n_598), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_637), .Y(n_660) );
OAI222xp33_ASAP7_75t_L g661 ( .A1(n_645), .A2(n_613), .B1(n_605), .B2(n_576), .C1(n_567), .C2(n_569), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_653), .B(n_571), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_627), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_623), .B(n_603), .Y(n_664) );
AOI21xp33_ASAP7_75t_SL g665 ( .A1(n_650), .A2(n_613), .B(n_604), .Y(n_665) );
OAI322xp33_ASAP7_75t_L g666 ( .A1(n_653), .A2(n_561), .A3(n_577), .B1(n_583), .B2(n_566), .C1(n_558), .C2(n_568), .Y(n_666) );
OAI221xp5_ASAP7_75t_SL g667 ( .A1(n_650), .A2(n_613), .B1(n_561), .B2(n_583), .C(n_577), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_628), .A2(n_631), .B1(n_624), .B2(n_635), .C(n_632), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_654), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_634), .A2(n_616), .B1(n_614), .B2(n_608), .C(n_606), .Y(n_670) );
AOI221x1_ASAP7_75t_SL g671 ( .A1(n_640), .A2(n_619), .B1(n_612), .B2(n_610), .C(n_611), .Y(n_671) );
OAI22xp33_ASAP7_75t_SL g672 ( .A1(n_629), .A2(n_611), .B1(n_589), .B2(n_615), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_630), .A2(n_563), .B1(n_602), .B2(n_599), .C(n_595), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_633), .A2(n_617), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_622), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_658), .A2(n_642), .B1(n_649), .B2(n_626), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_651), .A2(n_28), .B(n_33), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_641), .A2(n_35), .B1(n_36), .B2(n_38), .C(n_41), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_639), .B(n_42), .C(n_43), .D(n_44), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_647), .A2(n_55), .B1(n_56), .B2(n_60), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_639), .B(n_61), .C(n_63), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_646), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g683 ( .A1(n_647), .A2(n_66), .B(n_67), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_636), .A2(n_68), .B1(n_70), .B2(n_71), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_638), .B(n_72), .Y(n_685) );
A2O1A1Ixp33_ASAP7_75t_L g686 ( .A1(n_657), .A2(n_76), .B(n_78), .C(n_79), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g687 ( .A1(n_644), .A2(n_83), .B(n_84), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_648), .B(n_87), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g689 ( .A1(n_652), .A2(n_89), .B(n_92), .C(n_656), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g690 ( .A1(n_655), .A2(n_650), .B1(n_628), .B2(n_631), .C(n_623), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_690), .B(n_668), .C(n_665), .Y(n_691) );
AOI221x1_ASAP7_75t_L g692 ( .A1(n_672), .A2(n_664), .B1(n_683), .B2(n_676), .C(n_681), .Y(n_692) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_667), .B(n_680), .C(n_663), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_671), .B(n_659), .Y(n_694) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_679), .B(n_661), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_675), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_691), .B(n_686), .C(n_677), .D(n_689), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_696), .Y(n_698) );
NOR3xp33_ASAP7_75t_SL g699 ( .A(n_693), .B(n_670), .C(n_677), .Y(n_699) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_694), .B(n_674), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_698), .B(n_697), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_700), .B(n_692), .Y(n_702) );
OR2x2_ASAP7_75t_L g703 ( .A(n_699), .B(n_660), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_702), .B(n_695), .Y(n_704) );
XNOR2x1_ASAP7_75t_L g705 ( .A(n_703), .B(n_684), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_704), .Y(n_706) );
AOI22x1_ASAP7_75t_L g707 ( .A1(n_705), .A2(n_701), .B1(n_669), .B2(n_662), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_682), .B1(n_685), .B2(n_666), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_708), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_709), .A2(n_707), .B1(n_706), .B2(n_673), .Y(n_710) );
OR2x6_ASAP7_75t_L g711 ( .A(n_710), .B(n_688), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_711), .A2(n_687), .B1(n_625), .B2(n_678), .Y(n_712) );
endmodule