module fake_jpeg_17641_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_49),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_50),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_17),
.A2(n_3),
.B(n_4),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_53),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_46),
.B1(n_39),
.B2(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_70),
.B1(n_74),
.B2(n_43),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_25),
.B1(n_33),
.B2(n_18),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_76),
.B1(n_47),
.B2(n_4),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_35),
.A2(n_23),
.B1(n_24),
.B2(n_18),
.Y(n_70)
);

OA22x2_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_33),
.B1(n_25),
.B2(n_32),
.Y(n_71)
);

AO22x1_ASAP7_75t_SL g93 ( 
.A1(n_71),
.A2(n_26),
.B1(n_16),
.B2(n_44),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_35),
.A2(n_24),
.B1(n_32),
.B2(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_32),
.B1(n_26),
.B2(n_16),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_30),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_34),
.B1(n_30),
.B2(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_82),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_40),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_50),
.C(n_45),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_97),
.Y(n_108)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_44),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_93),
.Y(n_110)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_100),
.B1(n_59),
.B2(n_68),
.Y(n_119)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_34),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_43),
.B1(n_41),
.B2(n_48),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_116)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_51),
.B1(n_50),
.B2(n_6),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_121),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_95),
.B(n_81),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_63),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_71),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_71),
.B(n_64),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_94),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_140),
.B(n_89),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_107),
.B(n_108),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_142),
.B(n_145),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_111),
.B1(n_119),
.B2(n_101),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_149),
.B1(n_125),
.B2(n_109),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_93),
.B(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_137),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_63),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_91),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_81),
.B1(n_64),
.B2(n_59),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_144),
.B1(n_148),
.B2(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_96),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_72),
.B1(n_68),
.B2(n_76),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_87),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_108),
.B(n_78),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_79),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_105),
.B1(n_104),
.B2(n_98),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_154),
.A2(n_160),
.B1(n_60),
.B2(n_114),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_109),
.B1(n_125),
.B2(n_103),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_115),
.B1(n_118),
.B2(n_124),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_164),
.B1(n_166),
.B2(n_72),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_166),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_165),
.B(n_138),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_132),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_131),
.B(n_128),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_149),
.B(n_114),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_125),
.Y(n_171)
);

XOR2x1_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_137),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_148),
.B1(n_141),
.B2(n_133),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_191),
.B1(n_160),
.B2(n_163),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_133),
.C(n_140),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_181),
.C(n_186),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_189),
.B(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_169),
.C(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_159),
.B1(n_151),
.B2(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_158),
.C(n_139),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_135),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_160),
.C(n_163),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_117),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_170),
.B(n_155),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_174),
.B(n_191),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_167),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_202),
.C(n_206),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_153),
.B1(n_159),
.B2(n_160),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_178),
.B1(n_180),
.B2(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_174),
.B(n_181),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_211),
.B(n_213),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_177),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_109),
.Y(n_217)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_186),
.B(n_187),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_198),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_212),
.A2(n_208),
.B1(n_207),
.B2(n_188),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_226),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_211),
.A2(n_193),
.B(n_205),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_230),
.C(n_210),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_201),
.C(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_221),
.C(n_220),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_14),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_231),
.B(n_217),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_193),
.A3(n_84),
.B1(n_99),
.B2(n_126),
.C1(n_106),
.C2(n_117),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_216),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_213),
.B(n_218),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_236),
.B(n_223),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_240),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_212),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_219),
.C(n_126),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_233),
.B(n_5),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_102),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_3),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_5),
.C(n_6),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.C(n_248),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_7),
.C(n_9),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_255),
.C(n_257),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_10),
.C(n_12),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_10),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_259),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_258),
.Y(n_262)
);


endmodule