module fake_jpeg_18484_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx11_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

OR2x4_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_27),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_23),
.B1(n_21),
.B2(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_13),
.B1(n_26),
.B2(n_18),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_20),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_36),
.B1(n_28),
.B2(n_18),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_58),
.B1(n_26),
.B2(n_13),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_29),
.B(n_19),
.C(n_25),
.Y(n_55)
);

AOI22x1_ASAP7_75t_R g71 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_15),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_31),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_61),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_63),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_15),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_34),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_70),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_19),
.B1(n_40),
.B2(n_37),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_55),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_15),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_80),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_45),
.B1(n_40),
.B2(n_37),
.Y(n_73)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_64),
.B1(n_50),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_50),
.B1(n_13),
.B2(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_65),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_15),
.C(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_53),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_20),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_69),
.B1(n_78),
.B2(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_49),
.B1(n_20),
.B2(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_59),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_72),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_104),
.C(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_98),
.B(n_105),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_73),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_82),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_73),
.C(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_82),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_73),
.C(n_9),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_12),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_104),
.C(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_112),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_92),
.B1(n_88),
.B2(n_94),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_99),
.Y(n_118)
);

AO221x1_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_83),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_116),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_98),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_119),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_100),
.C(n_94),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_111),
.B(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_122),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_4),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_83),
.B1(n_11),
.B2(n_10),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_117),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_0),
.B(n_3),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_127),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_0),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_0),
.Y(n_130)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_130),
.B(n_6),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_7),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_7),
.Y(n_135)
);


endmodule