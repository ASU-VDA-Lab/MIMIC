module fake_jpeg_1064_n_717 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_717);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_717;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_716;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_715;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_714;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_7),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_62),
.Y(n_193)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_64),
.Y(n_151)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_66),
.B(n_68),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_26),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_69),
.B(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_19),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_72),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_26),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_73),
.B(n_74),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_32),
.B(n_17),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_77),
.Y(n_155)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_79),
.B(n_83),
.Y(n_179)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_81),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_40),
.B(n_17),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_84),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_16),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_85),
.B(n_89),
.Y(n_224)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_20),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_86),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_106),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_96),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_98),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_99),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_102),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_103),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_23),
.B(n_16),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_123),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_16),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_116),
.Y(n_217)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_20),
.Y(n_121)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_47),
.B(n_15),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_20),
.B(n_1),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_124),
.B(n_6),
.Y(n_225)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_24),
.Y(n_125)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_20),
.Y(n_126)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_126),
.Y(n_216)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_35),
.Y(n_128)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_22),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_29),
.Y(n_159)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_35),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_131),
.A2(n_22),
.B1(n_14),
.B2(n_13),
.Y(n_178)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_30),
.Y(n_133)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_133),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_63),
.B1(n_67),
.B2(n_70),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_140),
.A2(n_147),
.B1(n_178),
.B2(n_186),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_64),
.A2(n_54),
.B1(n_48),
.B2(n_47),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_144),
.B(n_188),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_54),
.B1(n_48),
.B2(n_59),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_159),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_86),
.A2(n_29),
.B1(n_41),
.B2(n_59),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_181),
.Y(n_259)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_41),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_166),
.B(n_189),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_96),
.A2(n_55),
.B1(n_38),
.B2(n_22),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_65),
.A2(n_22),
.B1(n_55),
.B2(n_38),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_82),
.A2(n_44),
.B1(n_14),
.B2(n_4),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_87),
.A2(n_44),
.B1(n_3),
.B2(n_4),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_77),
.A2(n_44),
.B1(n_14),
.B2(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_81),
.B(n_2),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_103),
.B(n_2),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_192),
.B(n_196),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_103),
.B(n_2),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_110),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_197),
.A2(n_210),
.B1(n_218),
.B2(n_182),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_199),
.A2(n_200),
.B1(n_204),
.B2(n_214),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_124),
.A2(n_128),
.B1(n_113),
.B2(n_115),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_80),
.Y(n_202)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_120),
.B(n_3),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_205),
.B(n_209),
.Y(n_251)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_207),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_117),
.B(n_5),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_92),
.Y(n_213)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_99),
.Y(n_222)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_109),
.B(n_6),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_223),
.B(n_8),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g279 ( 
.A(n_225),
.B(n_10),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_104),
.A2(n_107),
.B1(n_112),
.B2(n_119),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_132),
.Y(n_253)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

BUFx4f_ASAP7_75t_SL g358 ( 
.A(n_231),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_161),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_232),
.B(n_236),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_122),
.B1(n_94),
.B2(n_75),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_233),
.A2(n_283),
.B1(n_293),
.B2(n_259),
.Y(n_343)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_235),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_161),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_142),
.B(n_62),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_237),
.B(n_244),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_199),
.A2(n_130),
.B1(n_72),
.B2(n_121),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_238),
.A2(n_291),
.B1(n_305),
.B2(n_171),
.Y(n_325)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_239),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_139),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_241),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_139),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_242),
.Y(n_357)
);

INVx11_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_243),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_150),
.B(n_7),
.Y(n_244)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_246),
.Y(n_328)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_247),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_186),
.A2(n_126),
.B1(n_100),
.B2(n_101),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_249),
.B(n_295),
.Y(n_365)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_198),
.Y(n_250)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_250),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_252),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_253),
.A2(n_254),
.B1(n_262),
.B2(n_292),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_201),
.A2(n_108),
.B1(n_114),
.B2(n_95),
.Y(n_254)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_149),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_134),
.B(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_258),
.B(n_271),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_151),
.Y(n_261)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_148),
.A2(n_95),
.B1(n_84),
.B2(n_10),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_263),
.Y(n_316)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_170),
.Y(n_265)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_265),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_164),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_267),
.B(n_268),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_180),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_269),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_153),
.B(n_8),
.C(n_9),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_270),
.B(n_279),
.C(n_252),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_8),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_273),
.Y(n_361)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_141),
.A2(n_8),
.B(n_9),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_275),
.B(n_278),
.Y(n_330)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_143),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_277),
.B(n_307),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_298),
.Y(n_326)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_172),
.Y(n_280)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g283 ( 
.A1(n_226),
.A2(n_167),
.B1(n_163),
.B2(n_197),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_155),
.Y(n_284)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_284),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_177),
.B(n_10),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_244),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_177),
.B(n_138),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_286),
.B(n_312),
.Y(n_346)
);

CKINVDCx6p67_ASAP7_75t_R g287 ( 
.A(n_185),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_287),
.Y(n_370)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_155),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_294),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_147),
.A2(n_226),
.B1(n_176),
.B2(n_174),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_152),
.A2(n_143),
.B1(n_136),
.B2(n_146),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_210),
.A2(n_184),
.B1(n_154),
.B2(n_135),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_136),
.Y(n_294)
);

AOI32xp33_ASAP7_75t_L g295 ( 
.A1(n_191),
.A2(n_169),
.A3(n_145),
.B1(n_146),
.B2(n_214),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_296),
.A2(n_299),
.B1(n_208),
.B2(n_195),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_156),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_301),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_193),
.Y(n_298)
);

BUFx8_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_135),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_173),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_304),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_162),
.A2(n_229),
.B(n_206),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_221),
.B(n_204),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_309),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_137),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_173),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_310),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_228),
.B(n_183),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_137),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_228),
.B(n_208),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_281),
.A2(n_171),
.B1(n_227),
.B2(n_162),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_314),
.A2(n_349),
.B1(n_350),
.B2(n_368),
.Y(n_423)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_303),
.A2(n_194),
.B1(n_206),
.B2(n_227),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_317),
.A2(n_325),
.B1(n_263),
.B2(n_242),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_329),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_281),
.A2(n_305),
.B1(n_253),
.B2(n_237),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_342),
.B1(n_272),
.B2(n_256),
.Y(n_382)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_249),
.A2(n_175),
.B1(n_190),
.B2(n_194),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_SL g395 ( 
.A1(n_337),
.A2(n_299),
.B(n_246),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_303),
.A2(n_175),
.B1(n_190),
.B2(n_158),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_339),
.A2(n_352),
.B1(n_287),
.B2(n_243),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_253),
.A2(n_158),
.B1(n_195),
.B2(n_160),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_343),
.B(n_337),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_344),
.B(n_348),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_285),
.B(n_258),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g349 ( 
.A1(n_283),
.A2(n_293),
.B1(n_301),
.B2(n_273),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_L g350 ( 
.A1(n_241),
.A2(n_247),
.B1(n_310),
.B2(n_257),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_233),
.A2(n_306),
.B1(n_309),
.B2(n_274),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_300),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_251),
.A2(n_306),
.B1(n_309),
.B2(n_271),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_266),
.B(n_264),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_376),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_364),
.B(n_366),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_279),
.B(n_270),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_372),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_230),
.A2(n_255),
.B1(n_260),
.B2(n_248),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_265),
.B(n_234),
.C(n_261),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_248),
.C(n_302),
.Y(n_390)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_261),
.A2(n_234),
.A3(n_288),
.B1(n_282),
.B2(n_260),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_245),
.B(n_255),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_308),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_297),
.B(n_250),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_324),
.A2(n_287),
.B(n_240),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_377),
.A2(n_424),
.B(n_425),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_378),
.A2(n_381),
.B(n_387),
.Y(n_445)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_358),
.Y(n_379)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_379),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_342),
.A2(n_287),
.B1(n_298),
.B2(n_231),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_382),
.A2(n_395),
.B1(n_415),
.B2(n_420),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_334),
.B(n_245),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_385),
.B(n_393),
.Y(n_439)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_313),
.A2(n_239),
.B1(n_289),
.B2(n_276),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_390),
.B(n_323),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_323),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_402),
.Y(n_432)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_347),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_394),
.B(n_399),
.Y(n_451)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_396),
.Y(n_431)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_318),
.B(n_235),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_375),
.Y(n_400)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_400),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_333),
.A2(n_299),
.B(n_294),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_401),
.A2(n_406),
.B(n_363),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_346),
.B(n_235),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_364),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_347),
.B(n_320),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_405),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_328),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_323),
.A2(n_365),
.B(n_370),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

AND2x2_ASAP7_75t_SL g408 ( 
.A(n_326),
.B(n_318),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_408),
.Y(n_442)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_409),
.Y(n_462)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_316),
.Y(n_410)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_410),
.Y(n_464)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_372),
.Y(n_411)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_341),
.B(n_369),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_416),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_363),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_414),
.A2(n_358),
.B1(n_357),
.B2(n_363),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_343),
.A2(n_365),
.B1(n_349),
.B2(n_360),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_417),
.B(n_421),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_338),
.B(n_348),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_418),
.B(n_422),
.Y(n_434)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_338),
.B(n_344),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_326),
.A2(n_353),
.B(n_370),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_326),
.A2(n_374),
.B(n_335),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_321),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_427),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_335),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_429),
.B(n_440),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_411),
.A2(n_314),
.B1(n_337),
.B2(n_330),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_438),
.A2(n_447),
.B1(n_456),
.B2(n_465),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_419),
.B(n_330),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_441),
.B(n_444),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_419),
.B(n_340),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_420),
.A2(n_337),
.B1(n_371),
.B2(n_323),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_403),
.B(n_323),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_449),
.C(n_460),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_391),
.B(n_356),
.C(n_340),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_393),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_469),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_388),
.B(n_356),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_455),
.B(n_457),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_389),
.A2(n_361),
.B1(n_367),
.B2(n_359),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_426),
.B(n_373),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_415),
.A2(n_350),
.B1(n_368),
.B2(n_361),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_458),
.A2(n_423),
.B1(n_383),
.B2(n_420),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_408),
.B(n_331),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_461),
.A2(n_396),
.B(n_379),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_389),
.A2(n_367),
.B1(n_359),
.B2(n_357),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_405),
.B(n_373),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g494 ( 
.A(n_467),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_404),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_473),
.A2(n_482),
.B1(n_492),
.B2(n_495),
.Y(n_520)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_474),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_434),
.B(n_400),
.Y(n_475)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_475),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_466),
.A2(n_420),
.B1(n_397),
.B2(n_384),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_476),
.A2(n_479),
.B(n_480),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_434),
.B(n_422),
.Y(n_478)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_406),
.B(n_401),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_461),
.A2(n_406),
.B(n_401),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_466),
.A2(n_382),
.B1(n_416),
.B2(n_399),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_481),
.A2(n_497),
.B(n_503),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_437),
.A2(n_423),
.B1(n_408),
.B2(n_378),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_483),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_450),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_493),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_429),
.B(n_408),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_488),
.C(n_496),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_SL g487 ( 
.A1(n_432),
.A2(n_395),
.B(n_390),
.C(n_381),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_490),
.B(n_506),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_390),
.C(n_418),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_444),
.B(n_385),
.Y(n_489)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_489),
.Y(n_547)
);

A2O1A1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_432),
.A2(n_424),
.B(n_394),
.C(n_402),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_437),
.A2(n_423),
.B1(n_387),
.B2(n_425),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_435),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_452),
.A2(n_380),
.B1(n_413),
.B2(n_377),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_448),
.B(n_392),
.C(n_398),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_442),
.A2(n_407),
.B(n_409),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_451),
.B(n_380),
.Y(n_498)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_498),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_421),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_499),
.A2(n_509),
.B(n_443),
.Y(n_529)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_501),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_465),
.A2(n_417),
.B1(n_427),
.B2(n_410),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_502),
.A2(n_430),
.B1(n_433),
.B2(n_459),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_457),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_451),
.B(n_410),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_505),
.B(n_462),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_446),
.A2(n_319),
.B(n_414),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_447),
.A2(n_438),
.B1(n_456),
.B2(n_453),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_507),
.A2(n_442),
.B1(n_453),
.B2(n_458),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_443),
.B(n_386),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_514),
.A2(n_524),
.B1(n_526),
.B2(n_532),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_448),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_516),
.B(n_519),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_484),
.Y(n_519)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_522),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_482),
.A2(n_470),
.B1(n_454),
.B2(n_439),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_491),
.A2(n_454),
.B1(n_439),
.B2(n_460),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_500),
.B(n_440),
.C(n_449),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_527),
.B(n_538),
.C(n_542),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_484),
.B(n_440),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_528),
.B(n_540),
.Y(n_579)
);

INVxp33_ASAP7_75t_L g555 ( 
.A(n_529),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_498),
.B(n_441),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_530),
.B(n_537),
.Y(n_572)
);

NAND4xp25_ASAP7_75t_SL g531 ( 
.A(n_505),
.B(n_446),
.C(n_345),
.D(n_455),
.Y(n_531)
);

BUFx12f_ASAP7_75t_L g568 ( 
.A(n_531),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_491),
.A2(n_507),
.B1(n_492),
.B2(n_473),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_533),
.A2(n_544),
.B1(n_494),
.B2(n_501),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_491),
.A2(n_460),
.B1(n_449),
.B2(n_433),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_534),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_479),
.A2(n_445),
.B(n_431),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_535),
.A2(n_536),
.B(n_480),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_479),
.A2(n_431),
.B(n_459),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_494),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_500),
.B(n_462),
.C(n_445),
.Y(n_538)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_539),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_484),
.B(n_331),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_471),
.B(n_463),
.Y(n_541)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_541),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_500),
.B(n_464),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_496),
.B(n_464),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_546),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_507),
.A2(n_436),
.B1(n_468),
.B2(n_463),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_490),
.Y(n_545)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_545),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_496),
.B(n_327),
.Y(n_546)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_549),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_548),
.B(n_472),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_L g609 ( 
.A(n_550),
.B(n_508),
.C(n_509),
.Y(n_609)
);

XOR2x2_ASAP7_75t_L g552 ( 
.A(n_542),
.B(n_486),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_552),
.B(n_556),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_SL g553 ( 
.A(n_528),
.B(n_486),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_SL g595 ( 
.A(n_553),
.B(n_583),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_525),
.A2(n_503),
.B(n_506),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_554),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_518),
.A2(n_525),
.B(n_515),
.Y(n_556)
);

CKINVDCx14_ASAP7_75t_R g557 ( 
.A(n_523),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_557),
.A2(n_558),
.B1(n_481),
.B2(n_474),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_511),
.B(n_471),
.Y(n_559)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_559),
.Y(n_592)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_523),
.Y(n_564)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_564),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_535),
.A2(n_476),
.B(n_481),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_565),
.B(n_570),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_518),
.A2(n_490),
.B(n_487),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_566),
.B(n_581),
.Y(n_608)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_541),
.Y(n_569)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_569),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_511),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_539),
.Y(n_571)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_571),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_536),
.Y(n_574)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_574),
.Y(n_588)
);

AOI322xp5_ASAP7_75t_L g577 ( 
.A1(n_548),
.A2(n_493),
.A3(n_475),
.B1(n_478),
.B2(n_485),
.C1(n_499),
.C2(n_489),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_577),
.B(n_582),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_519),
.B(n_495),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_578),
.B(n_540),
.Y(n_585)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_513),
.Y(n_580)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_580),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_515),
.A2(n_487),
.B(n_497),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_536),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_516),
.B(n_497),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_584),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_585),
.B(n_552),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_578),
.B(n_512),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_586),
.B(n_579),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_576),
.A2(n_520),
.B1(n_532),
.B2(n_524),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_589),
.A2(n_591),
.B1(n_599),
.B2(n_603),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_564),
.A2(n_520),
.B1(n_526),
.B2(n_510),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_572),
.B(n_472),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_593),
.B(n_598),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_551),
.B(n_512),
.C(n_543),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_559),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_584),
.A2(n_547),
.B1(n_510),
.B2(n_544),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_600),
.A2(n_554),
.B1(n_568),
.B2(n_560),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_551),
.B(n_546),
.C(n_538),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_601),
.B(n_553),
.C(n_579),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_561),
.A2(n_517),
.B1(n_547),
.B2(n_534),
.Y(n_603)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_606),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_561),
.A2(n_517),
.B1(n_521),
.B2(n_502),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_607),
.A2(n_609),
.B1(n_611),
.B2(n_562),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_555),
.A2(n_574),
.B1(n_571),
.B2(n_567),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_555),
.A2(n_558),
.B1(n_573),
.B2(n_566),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_613),
.Y(n_621)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_611),
.Y(n_614)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_614),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_SL g644 ( 
.A(n_615),
.B(n_616),
.Y(n_644)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_596),
.Y(n_617)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_617),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_598),
.B(n_586),
.C(n_601),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_618),
.B(n_619),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_603),
.B(n_563),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_585),
.B(n_563),
.C(n_575),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_622),
.B(n_626),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_594),
.A2(n_549),
.B(n_556),
.Y(n_624)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_624),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_625),
.Y(n_650)
);

XOR2x2_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_581),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_592),
.B(n_560),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_627),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_608),
.B(n_575),
.C(n_573),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_628),
.B(n_638),
.C(n_595),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_597),
.A2(n_580),
.B1(n_476),
.B2(n_569),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_629),
.B(n_631),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_630),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.Y(n_640)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_596),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_591),
.B(n_583),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_632),
.B(n_637),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g634 ( 
.A1(n_589),
.A2(n_565),
.B1(n_568),
.B2(n_487),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_604),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_590),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_600),
.A2(n_568),
.B1(n_487),
.B2(n_477),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_641),
.B(n_653),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_633),
.A2(n_612),
.B(n_587),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_646),
.A2(n_654),
.B(n_645),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_628),
.B(n_618),
.C(n_615),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_647),
.B(n_648),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_622),
.B(n_587),
.C(n_610),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_619),
.B(n_610),
.C(n_608),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_651),
.B(n_652),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_626),
.B(n_602),
.C(n_607),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_616),
.B(n_621),
.C(n_620),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_621),
.B(n_588),
.C(n_595),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_654),
.B(n_657),
.C(n_638),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_614),
.B(n_588),
.C(n_527),
.Y(n_657)
);

FAx1_ASAP7_75t_L g659 ( 
.A(n_624),
.B(n_590),
.CI(n_605),
.CON(n_659),
.SN(n_659)
);

CKINVDCx16_ASAP7_75t_R g671 ( 
.A(n_659),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_658),
.B(n_632),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_660),
.B(n_663),
.Y(n_687)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_643),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_661),
.B(n_664),
.Y(n_679)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_651),
.B(n_634),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_650),
.A2(n_623),
.B1(n_627),
.B2(n_617),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_639),
.B(n_637),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_665),
.B(n_668),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_649),
.B(n_653),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_666),
.B(n_667),
.Y(n_683)
);

XNOR2xp5_ASAP7_75t_L g667 ( 
.A(n_648),
.B(n_630),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_647),
.B(n_508),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_669),
.A2(n_641),
.B(n_652),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_657),
.B(n_568),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_670),
.B(n_674),
.Y(n_691)
);

AOI21xp33_ASAP7_75t_L g689 ( 
.A1(n_673),
.A2(n_677),
.B(n_412),
.Y(n_689)
);

XNOR2xp5_ASAP7_75t_L g674 ( 
.A(n_656),
.B(n_531),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_659),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_SL g685 ( 
.A1(n_675),
.A2(n_412),
.B1(n_428),
.B2(n_414),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_655),
.A2(n_487),
.B1(n_428),
.B2(n_412),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_662),
.A2(n_644),
.B(n_659),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_678),
.A2(n_681),
.B(n_682),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_680),
.B(n_685),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_668),
.A2(n_640),
.B(n_642),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_676),
.A2(n_640),
.B(n_639),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_663),
.B(n_667),
.C(n_672),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_686),
.B(n_688),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_R g688 ( 
.A(n_671),
.B(n_327),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_689),
.B(n_690),
.Y(n_697)
);

OAI21xp33_ASAP7_75t_L g690 ( 
.A1(n_675),
.A2(n_428),
.B(n_414),
.Y(n_690)
);

MAJIxp5_ASAP7_75t_L g692 ( 
.A(n_686),
.B(n_660),
.C(n_670),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_692),
.B(n_694),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g694 ( 
.A(n_683),
.B(n_674),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_684),
.B(n_665),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_695),
.A2(n_679),
.B(n_357),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_SL g696 ( 
.A1(n_687),
.A2(n_345),
.B(n_319),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_696),
.A2(n_701),
.B(n_354),
.Y(n_706)
);

MAJIxp5_ASAP7_75t_L g700 ( 
.A(n_687),
.B(n_359),
.C(n_367),
.Y(n_700)
);

XNOR2xp5_ASAP7_75t_L g703 ( 
.A(n_700),
.B(n_690),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_691),
.B(n_386),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_693),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_702),
.B(n_703),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_704),
.B(n_705),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_698),
.B(n_351),
.Y(n_705)
);

MAJIxp5_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_701),
.C(n_699),
.Y(n_710)
);

MAJIxp5_ASAP7_75t_L g712 ( 
.A(n_710),
.B(n_707),
.C(n_709),
.Y(n_712)
);

BUFx24_ASAP7_75t_SL g711 ( 
.A(n_708),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_711),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_713),
.B(n_712),
.Y(n_714)
);

AOI21xp33_ASAP7_75t_L g715 ( 
.A1(n_714),
.A2(n_697),
.B(n_351),
.Y(n_715)
);

MAJIxp5_ASAP7_75t_L g716 ( 
.A(n_715),
.B(n_354),
.C(n_697),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_716),
.A2(n_351),
.B(n_707),
.Y(n_717)
);


endmodule