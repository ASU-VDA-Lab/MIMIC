module fake_jpeg_2221_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_60),
.Y(n_119)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_55),
.Y(n_112)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_62),
.B(n_70),
.Y(n_148)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g125 ( 
.A(n_65),
.Y(n_125)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_27),
.B(n_16),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_27),
.B(n_0),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_36),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_46),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_20),
.Y(n_120)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_102),
.Y(n_122)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_99),
.B(n_101),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_104),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_43),
.B1(n_45),
.B2(n_36),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_106),
.A2(n_116),
.B1(n_117),
.B2(n_128),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_111),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_43),
.B1(n_45),
.B2(n_36),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_30),
.B1(n_51),
.B2(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_158),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_51),
.B1(n_30),
.B2(n_26),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_127),
.A2(n_131),
.B1(n_138),
.B2(n_101),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_66),
.A2(n_20),
.B1(n_23),
.B2(n_47),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_58),
.A2(n_19),
.B1(n_28),
.B2(n_31),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_129),
.A2(n_146),
.B1(n_48),
.B2(n_4),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_51),
.B1(n_30),
.B2(n_26),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_61),
.A2(n_34),
.B1(n_35),
.B2(n_44),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_89),
.B(n_34),
.C(n_35),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_145),
.B(n_149),
.C(n_73),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_77),
.A2(n_28),
.B1(n_19),
.B2(n_47),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_64),
.B(n_44),
.C(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_55),
.B(n_31),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_55),
.B(n_23),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_74),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_54),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_42),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_167),
.B(n_172),
.Y(n_240)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_168),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_115),
.A2(n_68),
.B1(n_63),
.B2(n_87),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_169),
.A2(n_189),
.B(n_218),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_170),
.B(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_147),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_193),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_74),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_104),
.B1(n_103),
.B2(n_100),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_173),
.A2(n_194),
.B1(n_209),
.B2(n_118),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_159),
.B(n_87),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_174),
.B(n_177),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

AO21x2_ASAP7_75t_L g264 ( 
.A1(n_176),
.A2(n_3),
.B(n_4),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_102),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_178),
.Y(n_233)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_121),
.B(n_94),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_180),
.B(n_185),
.Y(n_248)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_181),
.Y(n_239)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_143),
.A2(n_131),
.B1(n_127),
.B2(n_88),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_184),
.A2(n_215),
.B1(n_220),
.B2(n_14),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_134),
.B(n_80),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_15),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_190),
.Y(n_222)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_136),
.Y(n_187)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_122),
.A2(n_130),
.B1(n_112),
.B2(n_137),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_75),
.Y(n_190)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_117),
.A2(n_73),
.B(n_69),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_192),
.A2(n_141),
.B(n_4),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_93),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_91),
.B1(n_37),
.B2(n_33),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_205),
.Y(n_243)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_125),
.Y(n_199)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_0),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_204),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_109),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_211),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_140),
.B(n_113),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_140),
.B(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_219),
.Y(n_250)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_155),
.A2(n_37),
.B1(n_33),
.B2(n_69),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_2),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_212),
.B(n_188),
.C(n_171),
.Y(n_262)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_213),
.B(n_216),
.Y(n_267)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_217),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_106),
.A2(n_37),
.B1(n_33),
.B2(n_52),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_154),
.B(n_135),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_112),
.A2(n_37),
.B1(n_52),
.B2(n_48),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_109),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_113),
.B(n_3),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_3),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_220),
.A2(n_150),
.B1(n_144),
.B2(n_133),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_226),
.A2(n_231),
.B1(n_241),
.B2(n_261),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_184),
.A2(n_150),
.B1(n_144),
.B2(n_133),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_170),
.B(n_124),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_235),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_164),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_237),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_164),
.B(n_124),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_188),
.A2(n_132),
.B1(n_160),
.B2(n_136),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_177),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_269),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_262),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_176),
.A2(n_160),
.B1(n_132),
.B2(n_48),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_253),
.A2(n_265),
.B1(n_212),
.B2(n_168),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_255),
.B(n_272),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_251),
.B(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_197),
.B(n_3),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_266),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_264),
.A2(n_271),
.B1(n_226),
.B2(n_231),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_6),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_204),
.B(n_6),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_185),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_205),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_174),
.CI(n_196),
.CON(n_273),
.SN(n_273)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_273),
.B(n_301),
.Y(n_325)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_274),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_196),
.B(n_216),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_277),
.A2(n_278),
.B(n_279),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_192),
.B(n_196),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_280),
.B(n_298),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_206),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_292),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_180),
.C(n_183),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_304),
.C(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_283),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_256),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_287),
.Y(n_327)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_286),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_178),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_288),
.A2(n_306),
.B1(n_309),
.B2(n_292),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_234),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_196),
.B(n_202),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_290),
.A2(n_295),
.B(n_311),
.Y(n_345)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_242),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

AO22x1_ASAP7_75t_L g292 ( 
.A1(n_247),
.A2(n_191),
.B1(n_182),
.B2(n_178),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_243),
.B(n_212),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_297),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_233),
.B(n_193),
.Y(n_295)
);

BUFx8_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_296),
.A2(n_239),
.B1(n_270),
.B2(n_224),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_250),
.B(n_179),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_234),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_250),
.A2(n_193),
.B(n_166),
.C(n_200),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_299),
.B(n_300),
.Y(n_349)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_234),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_195),
.C(n_219),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_240),
.B(n_213),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_305),
.B(n_308),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_261),
.A2(n_264),
.B1(n_248),
.B2(n_267),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_207),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_313),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_251),
.B(n_198),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_264),
.A2(n_214),
.B1(n_175),
.B2(n_210),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_267),
.A2(n_217),
.B(n_211),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_241),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_312),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_268),
.A2(n_181),
.B(n_187),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_254),
.B(n_264),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_210),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_316),
.Y(n_347)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_211),
.B(n_208),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_248),
.B(n_208),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_249),
.B(n_239),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_240),
.B(n_175),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_SL g337 ( 
.A(n_318),
.B(n_232),
.C(n_246),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_222),
.B(n_8),
.C(n_9),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_313),
.A2(n_264),
.B1(n_265),
.B2(n_254),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_321),
.A2(n_326),
.B1(n_332),
.B2(n_340),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_310),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_322),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_323),
.A2(n_343),
.B(n_338),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_285),
.A2(n_278),
.B1(n_302),
.B2(n_312),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_263),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_328),
.B(n_276),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_296),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_330),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_296),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_354),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_239),
.B(n_246),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_338),
.A2(n_316),
.B(n_295),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_294),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_346),
.C(n_351),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_306),
.A2(n_271),
.B1(n_249),
.B2(n_260),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_285),
.A2(n_228),
.B1(n_238),
.B2(n_260),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_342),
.A2(n_352),
.B1(n_360),
.B2(n_309),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_238),
.C(n_227),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_227),
.C(n_257),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_302),
.A2(n_258),
.B1(n_225),
.B2(n_224),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_258),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_355),
.C(n_289),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_296),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_257),
.C(n_252),
.Y(n_355)
);

AO22x1_ASAP7_75t_L g357 ( 
.A1(n_288),
.A2(n_317),
.B1(n_287),
.B2(n_277),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_361),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_292),
.A2(n_279),
.B1(n_299),
.B2(n_275),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_276),
.B(n_252),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_331),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_356),
.Y(n_367)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_273),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_377),
.C(n_379),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_348),
.A2(n_314),
.B1(n_316),
.B2(n_311),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_372),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_375),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_303),
.Y(n_374)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_320),
.Y(n_376)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_301),
.C(n_287),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_378),
.A2(n_380),
.B(n_323),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_273),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_293),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_308),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_351),
.Y(n_398)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_383),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_331),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_342),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_344),
.A2(n_317),
.B1(n_315),
.B2(n_295),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_319),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_307),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_390),
.C(n_355),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_300),
.C(n_284),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_291),
.Y(n_392)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_392),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_334),
.B(n_286),
.Y(n_393)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_393),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_320),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_394),
.A2(n_396),
.B1(n_397),
.B2(n_329),
.Y(n_427)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_346),
.B(n_283),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_344),
.A2(n_274),
.B1(n_225),
.B2(n_270),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_398),
.B(n_382),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_364),
.A2(n_332),
.B1(n_385),
.B2(n_389),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_414),
.B1(n_417),
.B2(n_357),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_341),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_406),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_341),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_371),
.A2(n_345),
.B(n_326),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_407),
.A2(n_426),
.B(n_378),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_370),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_364),
.A2(n_333),
.B1(n_340),
.B2(n_360),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_392),
.Y(n_416)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_416),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_389),
.A2(n_333),
.B1(n_347),
.B2(n_349),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_393),
.Y(n_418)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_418),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_353),
.C(n_327),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_422),
.C(n_429),
.Y(n_439)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_324),
.Y(n_421)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_327),
.C(n_345),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_347),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_427),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_373),
.B(n_327),
.C(n_320),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_425),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_441),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_399),
.A2(n_414),
.B1(n_408),
.B2(n_357),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_432),
.A2(n_407),
.B1(n_410),
.B2(n_416),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_365),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_433),
.B(n_434),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_424),
.B(n_375),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_436),
.B(n_448),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_437),
.A2(n_402),
.B(n_423),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_369),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_388),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_379),
.C(n_371),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_419),
.C(n_429),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_445),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_362),
.Y(n_444)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_406),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_418),
.B1(n_410),
.B2(n_397),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_409),
.B(n_386),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_362),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_453),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_380),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_451),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_395),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_350),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_421),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_455),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_420),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_457),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_458),
.B(n_460),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_422),
.C(n_403),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_403),
.C(n_415),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_462),
.B(n_467),
.Y(n_489)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_464),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_446),
.A2(n_452),
.B1(n_438),
.B2(n_447),
.Y(n_466)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_466),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_415),
.C(n_426),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_401),
.C(n_354),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_469),
.B(n_470),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_438),
.A2(n_321),
.B1(n_352),
.B2(n_402),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_401),
.C(n_330),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_478),
.C(n_443),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_428),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_474),
.B(n_452),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_476),
.A2(n_449),
.B(n_444),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_391),
.C(n_368),
.Y(n_478)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_479),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_456),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_483),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_450),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_494),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_435),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_487),
.Y(n_502)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_486),
.A2(n_469),
.B1(n_472),
.B2(n_460),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_435),
.Y(n_487)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_488),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_448),
.C(n_436),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_492),
.B(n_493),
.C(n_458),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_442),
.C(n_437),
.Y(n_493)
);

AO21x1_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_446),
.B(n_432),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_491),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_481),
.A2(n_463),
.B1(n_477),
.B2(n_467),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_504),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_490),
.A2(n_400),
.B1(n_367),
.B2(n_383),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_501),
.A2(n_13),
.B1(n_14),
.B2(n_510),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_505),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_473),
.Y(n_504)
);

XOR2x1_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_465),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_468),
.C(n_465),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_507),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_486),
.A2(n_468),
.B1(n_225),
.B2(n_11),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_9),
.C(n_10),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_509),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_11),
.C(n_12),
.Y(n_509)
);

NOR2x1_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_493),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_511),
.A2(n_521),
.B(n_506),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_484),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_512),
.B(n_514),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_505),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_495),
.C(n_481),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_518),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_494),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_504),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_502),
.A2(n_488),
.B(n_479),
.Y(n_521)
);

AO21x1_ASAP7_75t_L g524 ( 
.A1(n_522),
.A2(n_499),
.B(n_501),
.Y(n_524)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_524),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_509),
.Y(n_525)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_525),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_527),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_516),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_528),
.A2(n_529),
.B(n_530),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_508),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_534),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_535),
.A2(n_536),
.B(n_537),
.Y(n_539)
);

OAI21x1_ASAP7_75t_SL g536 ( 
.A1(n_533),
.A2(n_523),
.B(n_513),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_512),
.Y(n_537)
);

OAI321xp33_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_531),
.A3(n_520),
.B1(n_517),
.B2(n_526),
.C(n_514),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_526),
.C(n_519),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_539),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_14),
.Y(n_542)
);


endmodule