module fake_jpeg_12622_n_444 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_444);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_444;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_14),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_57),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_58),
.B(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_64),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_15),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_68),
.B(n_69),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_73),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_79),
.Y(n_136)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_81),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_20),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2x1_ASAP7_75t_SL g176 ( 
.A(n_82),
.B(n_101),
.Y(n_176)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_89),
.B(n_90),
.Y(n_144)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_94),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_43),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_105),
.Y(n_118)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_34),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_20),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_104),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_20),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_112),
.Y(n_163)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_111),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_34),
.B(n_0),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_39),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_113),
.B(n_114),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_115),
.B(n_54),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_43),
.B1(n_44),
.B2(n_29),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_122),
.A2(n_149),
.B1(n_177),
.B2(n_185),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_43),
.B1(n_39),
.B2(n_27),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_123),
.A2(n_125),
.B1(n_131),
.B2(n_147),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_25),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_124),
.B(n_152),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_61),
.A2(n_39),
.B1(n_27),
.B2(n_18),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_36),
.B(n_50),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_129),
.A2(n_173),
.B(n_180),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_92),
.B1(n_114),
.B2(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_166),
.B1(n_172),
.B2(n_109),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_72),
.A2(n_27),
.B1(n_18),
.B2(n_23),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_56),
.B(n_24),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_159),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_100),
.A2(n_18),
.B1(n_23),
.B2(n_31),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_71),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_148),
.B(n_171),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_59),
.A2(n_19),
.B1(n_30),
.B2(n_50),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_86),
.B(n_35),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_60),
.B(n_45),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_71),
.A2(n_37),
.B(n_24),
.C(n_45),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_63),
.B(n_42),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_184),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_23),
.B1(n_35),
.B2(n_38),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_37),
.C(n_42),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_7),
.C(n_97),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_67),
.A2(n_38),
.B1(n_32),
.B2(n_30),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_106),
.B(n_32),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_175),
.B(n_178),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_55),
.A2(n_19),
.B1(n_54),
.B2(n_48),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_66),
.B(n_54),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_74),
.A2(n_54),
.B1(n_48),
.B2(n_2),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_78),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_66),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_182),
.A2(n_183),
.B1(n_113),
.B2(n_7),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_84),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_84),
.B(n_3),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_98),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_93),
.B(n_5),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_181),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_78),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_168),
.B1(n_118),
.B2(n_186),
.Y(n_248)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_189),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_93),
.B1(n_97),
.B2(n_113),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_190),
.A2(n_220),
.B1(n_227),
.B2(n_235),
.Y(n_288)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_192),
.Y(n_279)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_57),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_198),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_130),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_197),
.A2(n_204),
.B1(n_209),
.B2(n_236),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_199),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_144),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_201),
.B(n_207),
.Y(n_271)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_156),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_210),
.B(n_216),
.Y(n_272)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_164),
.B1(n_159),
.B2(n_184),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_151),
.B1(n_142),
.B2(n_126),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_135),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_176),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_217),
.B(n_226),
.Y(n_283)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_155),
.A2(n_139),
.B1(n_179),
.B2(n_121),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_152),
.B(n_124),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_222),
.B(n_229),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_224),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_140),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_151),
.Y(n_225)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_187),
.A2(n_170),
.B1(n_178),
.B2(n_160),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_117),
.B(n_138),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_162),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_230),
.B(n_239),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_128),
.Y(n_231)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_231),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_119),
.B(n_121),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_165),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_179),
.A2(n_175),
.B1(n_139),
.B2(n_127),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_167),
.A2(n_176),
.B1(n_146),
.B2(n_128),
.Y(n_236)
);

OR2x2_ASAP7_75t_SL g237 ( 
.A(n_153),
.B(n_165),
.Y(n_237)
);

OR2x2_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_241),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

BUFx24_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_146),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_148),
.B(n_118),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_250),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_126),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_167),
.A2(n_137),
.B1(n_168),
.B2(n_154),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_157),
.A2(n_158),
.B1(n_141),
.B2(n_161),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_225),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_137),
.Y(n_247)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_132),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_249),
.A2(n_225),
.B(n_231),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_118),
.Y(n_250)
);

AOI221xp5_ASAP7_75t_L g319 ( 
.A1(n_251),
.A2(n_261),
.B1(n_286),
.B2(n_256),
.C(n_284),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_171),
.Y(n_255)
);

A2O1A1O1Ixp25_ASAP7_75t_L g310 ( 
.A1(n_255),
.A2(n_265),
.B(n_268),
.C(n_280),
.D(n_284),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_217),
.A2(n_174),
.B1(n_126),
.B2(n_142),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_258),
.A2(n_290),
.B1(n_287),
.B2(n_292),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_212),
.A2(n_174),
.B1(n_186),
.B2(n_200),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_263),
.B1(n_274),
.B2(n_278),
.Y(n_302)
);

AOI32xp33_ASAP7_75t_L g261 ( 
.A1(n_213),
.A2(n_174),
.A3(n_200),
.B1(n_203),
.B2(n_232),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_228),
.A2(n_204),
.B1(n_203),
.B2(n_202),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_221),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_194),
.B(n_195),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_233),
.A2(n_246),
.B1(n_198),
.B2(n_242),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_196),
.A2(n_220),
.B1(n_235),
.B2(n_190),
.Y(n_278)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_196),
.B(n_223),
.Y(n_280)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_240),
.Y(n_284)
);

AND2x6_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_239),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_189),
.A2(n_193),
.B1(n_219),
.B2(n_218),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_278),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_234),
.A2(n_238),
.B1(n_215),
.B2(n_191),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_294),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_214),
.A2(n_226),
.B1(n_205),
.B2(n_206),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_249),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_298),
.B(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_265),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_303),
.B(n_313),
.Y(n_353)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_270),
.B1(n_263),
.B2(n_291),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_308),
.B1(n_324),
.B2(n_329),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_316),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_275),
.B(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_247),
.B1(n_245),
.B2(n_241),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_208),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_293),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_281),
.Y(n_315)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_315),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_260),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_317),
.A2(n_327),
.B1(n_328),
.B2(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_318),
.B(n_319),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_252),
.B(n_255),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_320),
.A2(n_310),
.B(n_306),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_252),
.B(n_283),
.C(n_280),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_279),
.C(n_296),
.Y(n_341)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_322),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_252),
.B(n_283),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_323),
.B(n_325),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_251),
.B(n_294),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_272),
.B(n_271),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_326),
.Y(n_359)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_254),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_253),
.A2(n_256),
.B1(n_286),
.B2(n_268),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_262),
.B(n_264),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_331),
.A2(n_325),
.B(n_300),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_259),
.A2(n_267),
.B1(n_297),
.B2(n_266),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_332),
.A2(n_279),
.B1(n_266),
.B2(n_296),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_302),
.A2(n_259),
.B1(n_267),
.B2(n_297),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_337),
.A2(n_352),
.B1(n_356),
.B2(n_357),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_334),
.C(n_344),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_321),
.C(n_320),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_341),
.C(n_354),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_305),
.A2(n_317),
.B1(n_314),
.B2(n_308),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_350),
.A2(n_318),
.B1(n_328),
.B2(n_330),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_302),
.A2(n_316),
.B1(n_299),
.B2(n_301),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_354),
.A2(n_344),
.B(n_343),
.Y(n_369)
);

NOR2x1_ASAP7_75t_R g355 ( 
.A(n_310),
.B(n_313),
.Y(n_355)
);

FAx1_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_334),
.CI(n_338),
.CON(n_378),
.SN(n_378)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_317),
.A2(n_312),
.B1(n_300),
.B2(n_325),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_312),
.A2(n_311),
.B1(n_315),
.B2(n_322),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g360 ( 
.A(n_339),
.B(n_331),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_360),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_374),
.B1(n_333),
.B2(n_336),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_345),
.Y(n_364)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_371),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_332),
.B1(n_327),
.B2(n_304),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_368),
.A2(n_379),
.B1(n_359),
.B2(n_358),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_369),
.A2(n_378),
.B(n_366),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_373),
.C(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_342),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_375),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_338),
.A2(n_350),
.B1(n_335),
.B2(n_353),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_376),
.B(n_380),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_357),
.B(n_353),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_377),
.A2(n_333),
.B(n_334),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_346),
.A2(n_337),
.B1(n_355),
.B2(n_349),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_346),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_365),
.A2(n_336),
.B1(n_355),
.B2(n_351),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_381),
.A2(n_386),
.B1(n_396),
.B2(n_361),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_390),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_384),
.A2(n_376),
.B(n_378),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_340),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_388),
.C(n_391),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_368),
.C(n_375),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_358),
.C(n_373),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_377),
.B1(n_362),
.B2(n_361),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_369),
.B(n_378),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_360),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_379),
.B1(n_363),
.B2(n_372),
.Y(n_396)
);

AOI21xp33_ASAP7_75t_L g398 ( 
.A1(n_389),
.A2(n_378),
.B(n_380),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_398),
.A2(n_409),
.B(n_410),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_400),
.A2(n_407),
.B(n_397),
.Y(n_417)
);

FAx1_ASAP7_75t_SL g401 ( 
.A(n_389),
.B(n_360),
.CI(n_364),
.CON(n_401),
.SN(n_401)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_404),
.Y(n_413)
);

BUFx12f_ASAP7_75t_SL g403 ( 
.A(n_391),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_403),
.A2(n_382),
.B(n_392),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_391),
.B(n_360),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_393),
.Y(n_405)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_405),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_406),
.A2(n_382),
.B1(n_393),
.B2(n_397),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_384),
.A2(n_395),
.B(n_390),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_408),
.A2(n_381),
.B(n_383),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_367),
.C(n_371),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_412),
.B(n_417),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_399),
.A2(n_396),
.B1(n_386),
.B2(n_392),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_414),
.A2(n_416),
.B1(n_402),
.B2(n_407),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_415),
.A2(n_394),
.B1(n_401),
.B2(n_404),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_410),
.A2(n_387),
.B1(n_394),
.B2(n_385),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_409),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_400),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_418),
.B(n_402),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_423),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_406),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_422),
.B(n_411),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g424 ( 
.A(n_417),
.B(n_414),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_424),
.A2(n_426),
.B(n_412),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_408),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_427),
.C(n_423),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_413),
.Y(n_432)
);

AO21x1_ASAP7_75t_L g437 ( 
.A1(n_429),
.A2(n_432),
.B(n_428),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_430),
.B(n_425),
.Y(n_435)
);

AOI21xp33_ASAP7_75t_L g433 ( 
.A1(n_421),
.A2(n_401),
.B(n_403),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_433),
.B(n_427),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_434),
.B(n_431),
.C(n_409),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_435),
.B(n_437),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_436),
.B(n_438),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_439),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_441),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_440),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_443),
.B(n_431),
.Y(n_444)
);


endmodule